//
// Conformal-LEC Version 20.10-d213 (02-Sep-2020)
//
module top(RI9871f50_143,RI9871e60_141,RI9871ed8_142,RI986f520_53,RI986f610_55,RI9872220_149,RI9872130_147,RI9871d70_139,RI986ddb0_3,
        RI986dcc0_1,RI9871de8_140,RI986df90_7,RI986dea0_5,RI986f8e0_61,RI9871fc8_144,RI9872040_145,RI986f430_51,RI986f340_49,RI9871c80_137,
        RI9871cf8_138,RI9871b18_134,RI986e260_13,RI986e350_15,RI9871c08_136,RI9871b90_135,RI98721a8_148,RI986e170_11,RI986e080_9,RI986f9d0_63,
        RI986e0f8_10,RI986e2d8_14,RI986e3c8_16,RI986dd38_2,RI986e1e8_12,RI986f4a8_52,RI986f3b8_50,RI986f598_54,RI986df18_6,RI986de28_4,
        RI986f688_56,RI986e008_8,RI986f958_62,RI986f700_57,RI98718c0_129,RI98720b8_146,RI986e710_23,RI986e620_21,RI986e530_19,RI986e440_17,
        RI986f7f0_59,RI98719b0_131,RI9871a28_132,RI9871aa0_133,RI9871938_130,RI9872310_151,RI9872298_150,RI986f160_45,RI98726d0_159,RI9872748_160,
        RI986f070_43,RI986ef80_41,RI986f250_47,RI98725e0_157,RI9872658_158,RI986ebc0_33,RI986ecb0_35,RI9872388_152,RI98727c0_161,RI986eda0_37,
        RI986ee90_39,RI9872478_154,RI9872400_153,RI986e800_25,RI986e8f0_27,RI98724f0_155,RI9872568_156,RI986e9e0_29,RI986ead0_31,RI98728b0_163,
        RI9872838_162,RI98715f0_123,RI9871500_121,RI98729a0_165,RI9872928_164,RI98717d0_127,RI9872a18_166,RI9872a90_167,RI98716e0_125,RI9871410_119,
        RI9871320_117,RI9872b08_168,RI9872b80_169,RI9871140_113,RI9871230_115,RI9872bf8_170,RI9872c70_171,RI9871050_111,RI9870c90_103,RI9872d60_173,
        RI9872ce8_172,RI9870ba0_101,RI9870e70_107,RI9872e50_175,RI9872dd8_174,RI98709c0_97,RI9870d80_105,RI9872f40_177,RI9872ec8_176,RI9870ab0_99,
        RI9870f60_109,RI9872fb8_178,RI9873030_179,RI9870150_79,RI9870060_77,RI986fe80_73,RI98730a8_180,RI9873120_181,RI986ff70_75,RI9873210_183,
        RI9873198_182,RI986fca0_69,RI986fd90_71,RI9873288_184,RI9873300_185,RI986fbb0_67,RI986fac0_65,RI98707e0_93,RI98733f0_187,RI9873378_186,
        RI98708d0_95,RI98734e0_189,RI9873468_188,RI98706f0_91,RI9870600_89,RI9873558_190,RI98735d0_191,RI9870240_81,RI9870330_83,RI9870510_87,
        RI9873648_192,RI9870420_85,RI986fa48_64,RI986f778_58,RI986f868_60,RI986e698_22,RI986e788_24,RI986e4b8_18,RI986e5a8_20,RI986f1d8_46,
        RI986f2c8_48,RI986f0e8_44,RI986eff8_42,RI986ec38_34,RI986ed28_36,RI986ee18_38,RI986ef08_40,RI986e878_26,RI986e968_28,RI986ea58_30,
        RI986eb48_32,RI9871668_124,RI9871578_122,RI9871758_126,RI9871848_128,RI9871488_120,RI9871398_118,RI98711b8_114,RI98712a8_116,RI98710c8_112,
        RI9870d08_104,RI9870c18_102,RI9870ee8_108,RI9870a38_98,RI9870df8_106,RI9870b28_100,RI9870fd8_110,RI98701c8_80,RI98700d8_78,RI986fef8_74,
        RI986ffe8_76,RI986fd18_70,RI986fe08_72,RI986fc28_68,RI986fb38_66,RI9870858_94,RI9870948_96,RI9870768_92,RI9870678_90,RI98702b8_82,
        RI98703a8_84,RI9870588_88,RI9870498_86,RI9874ae8_236,RI9874f20_245,RI98745c0_225,RI9874a70_235,RI9874548_224,RI98736c0_193,RI9873e40_209,
        RI9874c50_239,RI9874188_216,RI9874278_218,RI9873f30_211,RI9874ea8_244,RI98743e0_221,RI98744d0_223,RI9875358_254,RI9873b70_203,RI98749f8_234,
        RI9875178_250,RI9874458_222,RI9874098_214,RI9873eb8_210,RI9874818_230,RI9874db8_242,RI9875088_248,RI9874638_226,RI9874b60_237,RI9873738_194,
        RI9874cc8_240,RI9873918_198,RI9873cd8_206,RI9873be8_204,RI9875010_247,RI9875100_249,RI9874980_233,RI98747a0_229,RI9874020_213,RI9874110_215,
        RI98737b0_195,RI9874f98_246,RI9874bd8_238,RI9874890_231,RI9873fa8_212,RI9873a08_200,RI9873af8_202,RI98742f0_219,RI98751f0_251,RI9874200_217,
        RI98738a0_197,RI9873828_196,RI9875268_252,RI9874368_220,RI9873a80_201,RI9874728_228,RI9873d50_207,RI9873990_199,RI9874908_232,RI9874d40_241,
        RI98746b0_227,RI9874e30_243,RI9873c60_205,RI98752e0_253,RI9875448_256,RI98753d0_255,RI9873dc8_208,R_101_8a8e950,R_102_8a8f868,R_103_8a8f910,
        R_104_8a8f9b8,R_105_8a8fa60,R_106_8a8fb08,R_107_8a8fbb0,R_108_8a8fc58,R_109_8a8fd00,R_10a_8a8fda8,R_10b_8a8fe50,R_10c_8a8fef8,R_10d_8a8ffa0,
        R_10e_8a90048,R_10f_8a900f0,R_110_8a90198,R_111_8a90240,R_112_8a902e8,R_113_8a90390,R_114_8a90438,R_115_8a904e0,R_116_8a90588,R_117_8a90630,
        R_118_8a906d8,R_119_8a90780,R_11a_8a90828,R_11b_8a908d0,R_11c_8a90978,R_11d_8a90a20,R_11e_8a90ac8,R_11f_8a90b70,R_120_8a90c18,R_121_8a90cc0,
        R_122_8a90d68,R_123_8a90e10,R_124_8a90eb8,R_125_8a90f60,R_126_8a91008,R_127_8a910b0,R_128_8a91158,R_129_8a91200,R_12a_8a912a8,R_12b_8a91350,
        R_12c_8a913f8,R_12d_8a914a0,R_12e_8a91548,R_12f_8a915f0,R_130_8a91698,R_131_8a91740,R_132_8a917e8,R_133_8a91890,R_134_8a91938,R_135_8a919e0,
        R_136_8a91a88,R_137_8a91b30,R_138_8a91bd8,R_139_8a91c80,R_13a_8a91d28,R_13b_8a91dd0,R_13c_8a91e78,R_13d_8a91f20,R_13e_8a91fc8,R_13f_8a92070,
        R_140_8a92118,R_141_8a921c0,R_142_8a92268,R_143_8a92310,R_144_8a923b8,R_145_8a92460,R_146_8a92508,R_147_8a925b0,R_148_8a92658,R_149_8a92700,
        R_14a_8a927a8,R_14b_8a92850,R_14c_8a928f8,R_14d_8a929a0,R_14e_8a92a48,R_14f_8a92af0,R_150_8a92b98,R_151_8a92c40,R_152_8a92ce8,R_153_8a92d90,
        R_154_8a92e38,R_155_8a92ee0);
input RI9871f50_143,RI9871e60_141,RI9871ed8_142,RI986f520_53,RI986f610_55,RI9872220_149,RI9872130_147,RI9871d70_139,RI986ddb0_3,
        RI986dcc0_1,RI9871de8_140,RI986df90_7,RI986dea0_5,RI986f8e0_61,RI9871fc8_144,RI9872040_145,RI986f430_51,RI986f340_49,RI9871c80_137,
        RI9871cf8_138,RI9871b18_134,RI986e260_13,RI986e350_15,RI9871c08_136,RI9871b90_135,RI98721a8_148,RI986e170_11,RI986e080_9,RI986f9d0_63,
        RI986e0f8_10,RI986e2d8_14,RI986e3c8_16,RI986dd38_2,RI986e1e8_12,RI986f4a8_52,RI986f3b8_50,RI986f598_54,RI986df18_6,RI986de28_4,
        RI986f688_56,RI986e008_8,RI986f958_62,RI986f700_57,RI98718c0_129,RI98720b8_146,RI986e710_23,RI986e620_21,RI986e530_19,RI986e440_17,
        RI986f7f0_59,RI98719b0_131,RI9871a28_132,RI9871aa0_133,RI9871938_130,RI9872310_151,RI9872298_150,RI986f160_45,RI98726d0_159,RI9872748_160,
        RI986f070_43,RI986ef80_41,RI986f250_47,RI98725e0_157,RI9872658_158,RI986ebc0_33,RI986ecb0_35,RI9872388_152,RI98727c0_161,RI986eda0_37,
        RI986ee90_39,RI9872478_154,RI9872400_153,RI986e800_25,RI986e8f0_27,RI98724f0_155,RI9872568_156,RI986e9e0_29,RI986ead0_31,RI98728b0_163,
        RI9872838_162,RI98715f0_123,RI9871500_121,RI98729a0_165,RI9872928_164,RI98717d0_127,RI9872a18_166,RI9872a90_167,RI98716e0_125,RI9871410_119,
        RI9871320_117,RI9872b08_168,RI9872b80_169,RI9871140_113,RI9871230_115,RI9872bf8_170,RI9872c70_171,RI9871050_111,RI9870c90_103,RI9872d60_173,
        RI9872ce8_172,RI9870ba0_101,RI9870e70_107,RI9872e50_175,RI9872dd8_174,RI98709c0_97,RI9870d80_105,RI9872f40_177,RI9872ec8_176,RI9870ab0_99,
        RI9870f60_109,RI9872fb8_178,RI9873030_179,RI9870150_79,RI9870060_77,RI986fe80_73,RI98730a8_180,RI9873120_181,RI986ff70_75,RI9873210_183,
        RI9873198_182,RI986fca0_69,RI986fd90_71,RI9873288_184,RI9873300_185,RI986fbb0_67,RI986fac0_65,RI98707e0_93,RI98733f0_187,RI9873378_186,
        RI98708d0_95,RI98734e0_189,RI9873468_188,RI98706f0_91,RI9870600_89,RI9873558_190,RI98735d0_191,RI9870240_81,RI9870330_83,RI9870510_87,
        RI9873648_192,RI9870420_85,RI986fa48_64,RI986f778_58,RI986f868_60,RI986e698_22,RI986e788_24,RI986e4b8_18,RI986e5a8_20,RI986f1d8_46,
        RI986f2c8_48,RI986f0e8_44,RI986eff8_42,RI986ec38_34,RI986ed28_36,RI986ee18_38,RI986ef08_40,RI986e878_26,RI986e968_28,RI986ea58_30,
        RI986eb48_32,RI9871668_124,RI9871578_122,RI9871758_126,RI9871848_128,RI9871488_120,RI9871398_118,RI98711b8_114,RI98712a8_116,RI98710c8_112,
        RI9870d08_104,RI9870c18_102,RI9870ee8_108,RI9870a38_98,RI9870df8_106,RI9870b28_100,RI9870fd8_110,RI98701c8_80,RI98700d8_78,RI986fef8_74,
        RI986ffe8_76,RI986fd18_70,RI986fe08_72,RI986fc28_68,RI986fb38_66,RI9870858_94,RI9870948_96,RI9870768_92,RI9870678_90,RI98702b8_82,
        RI98703a8_84,RI9870588_88,RI9870498_86,RI9874ae8_236,RI9874f20_245,RI98745c0_225,RI9874a70_235,RI9874548_224,RI98736c0_193,RI9873e40_209,
        RI9874c50_239,RI9874188_216,RI9874278_218,RI9873f30_211,RI9874ea8_244,RI98743e0_221,RI98744d0_223,RI9875358_254,RI9873b70_203,RI98749f8_234,
        RI9875178_250,RI9874458_222,RI9874098_214,RI9873eb8_210,RI9874818_230,RI9874db8_242,RI9875088_248,RI9874638_226,RI9874b60_237,RI9873738_194,
        RI9874cc8_240,RI9873918_198,RI9873cd8_206,RI9873be8_204,RI9875010_247,RI9875100_249,RI9874980_233,RI98747a0_229,RI9874020_213,RI9874110_215,
        RI98737b0_195,RI9874f98_246,RI9874bd8_238,RI9874890_231,RI9873fa8_212,RI9873a08_200,RI9873af8_202,RI98742f0_219,RI98751f0_251,RI9874200_217,
        RI98738a0_197,RI9873828_196,RI9875268_252,RI9874368_220,RI9873a80_201,RI9874728_228,RI9873d50_207,RI9873990_199,RI9874908_232,RI9874d40_241,
        RI98746b0_227,RI9874e30_243,RI9873c60_205,RI98752e0_253,RI9875448_256,RI98753d0_255,RI9873dc8_208;
output R_101_8a8e950,R_102_8a8f868,R_103_8a8f910,R_104_8a8f9b8,R_105_8a8fa60,R_106_8a8fb08,R_107_8a8fbb0,R_108_8a8fc58,R_109_8a8fd00,
        R_10a_8a8fda8,R_10b_8a8fe50,R_10c_8a8fef8,R_10d_8a8ffa0,R_10e_8a90048,R_10f_8a900f0,R_110_8a90198,R_111_8a90240,R_112_8a902e8,R_113_8a90390,
        R_114_8a90438,R_115_8a904e0,R_116_8a90588,R_117_8a90630,R_118_8a906d8,R_119_8a90780,R_11a_8a90828,R_11b_8a908d0,R_11c_8a90978,R_11d_8a90a20,
        R_11e_8a90ac8,R_11f_8a90b70,R_120_8a90c18,R_121_8a90cc0,R_122_8a90d68,R_123_8a90e10,R_124_8a90eb8,R_125_8a90f60,R_126_8a91008,R_127_8a910b0,
        R_128_8a91158,R_129_8a91200,R_12a_8a912a8,R_12b_8a91350,R_12c_8a913f8,R_12d_8a914a0,R_12e_8a91548,R_12f_8a915f0,R_130_8a91698,R_131_8a91740,
        R_132_8a917e8,R_133_8a91890,R_134_8a91938,R_135_8a919e0,R_136_8a91a88,R_137_8a91b30,R_138_8a91bd8,R_139_8a91c80,R_13a_8a91d28,R_13b_8a91dd0,
        R_13c_8a91e78,R_13d_8a91f20,R_13e_8a91fc8,R_13f_8a92070,R_140_8a92118,R_141_8a921c0,R_142_8a92268,R_143_8a92310,R_144_8a923b8,R_145_8a92460,
        R_146_8a92508,R_147_8a925b0,R_148_8a92658,R_149_8a92700,R_14a_8a927a8,R_14b_8a92850,R_14c_8a928f8,R_14d_8a929a0,R_14e_8a92a48,R_14f_8a92af0,
        R_150_8a92b98,R_151_8a92c40,R_152_8a92ce8,R_153_8a92d90,R_154_8a92e38,R_155_8a92ee0;

wire \342_ZERO , \343_ONE , \344 , \345 , \346 , \347 , \348 , \349 , \350 ,
         \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 ,
         \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 ,
         \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 ,
         \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 ,
         \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 ,
         \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 ,
         \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 ,
         \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 ,
         \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 ,
         \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 ,
         \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 ,
         \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 ,
         \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 ,
         \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 ,
         \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 ,
         \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 ,
         \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 ,
         \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 ,
         \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 ,
         \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 ,
         \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 ,
         \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 ,
         \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 ,
         \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 ,
         \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 ,
         \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 ,
         \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 ,
         \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 ,
         \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 ,
         \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 ,
         \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 ,
         \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 ,
         \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 ,
         \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 ,
         \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 ,
         \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 ,
         \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 ,
         \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 ,
         \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 ,
         \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 ,
         \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 ,
         \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 ,
         \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 ,
         \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 ,
         \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 ,
         \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 ,
         \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 ,
         \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 ,
         \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 ,
         \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 ,
         \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 ,
         \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 ,
         \871 , \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 ,
         \881 , \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 ,
         \891 , \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 ,
         \901 , \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 ,
         \911 , \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 ,
         \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 ,
         \931 , \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 ,
         \941 , \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 ,
         \951 , \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 ,
         \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 ,
         \971 , \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 ,
         \981 , \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 ,
         \991 , \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 ,
         \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 ,
         \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 ,
         \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 ,
         \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 ,
         \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 ,
         \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 ,
         \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 ,
         \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 ,
         \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 ,
         \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 ,
         \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 ,
         \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 ,
         \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 ,
         \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 ,
         \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 ,
         \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 ,
         \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 ,
         \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 ,
         \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 ,
         \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 ,
         \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 ,
         \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 ,
         \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 ,
         \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 ,
         \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 ,
         \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 ,
         \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 ,
         \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 ,
         \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 ,
         \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 ,
         \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 ,
         \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 ,
         \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 ,
         \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 ,
         \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 ,
         \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 ,
         \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 ,
         \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 ,
         \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 ,
         \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 ,
         \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 ,
         \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 ,
         \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 ,
         \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 ,
         \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 ,
         \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 ,
         \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 ,
         \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 ,
         \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 ,
         \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 ,
         \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 ,
         \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 ,
         \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 ,
         \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 ,
         \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 ,
         \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 ,
         \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 ,
         \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 ,
         \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 ,
         \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 ,
         \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 ,
         \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 ,
         \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 ,
         \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 ,
         \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 ,
         \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 ,
         \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 ,
         \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 ,
         \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 ,
         \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 ,
         \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 ,
         \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 ,
         \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 ,
         \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 ,
         \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 ,
         \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 ,
         \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 ,
         \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 ,
         \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 ,
         \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 ,
         \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 ,
         \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 ,
         \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 ,
         \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 ,
         \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 ,
         \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 ,
         \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 ,
         \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 ,
         \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 ,
         \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 ,
         \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 ,
         \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 ,
         \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 ,
         \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 ,
         \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 ,
         \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 ,
         \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 ,
         \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 ,
         \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 ,
         \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 ,
         \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 ,
         \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 ,
         \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 ,
         \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 ,
         \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 ,
         \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 ,
         \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 ,
         \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 ,
         \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 ,
         \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 ,
         \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 ,
         \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 ,
         \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 ,
         \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 ,
         \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 ,
         \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 ,
         \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 ,
         \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 ,
         \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 ,
         \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 ,
         \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 ,
         \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 ,
         \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 ,
         \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 ,
         \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 ,
         \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 ,
         \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 ,
         \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 ,
         \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 ,
         \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 ,
         \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 ,
         \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 ,
         \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 ,
         \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 ,
         \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 ,
         \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 ,
         \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 ,
         \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 ,
         \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 ,
         \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 ,
         \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 ,
         \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 ,
         \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 ,
         \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 ,
         \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 ,
         \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 ,
         \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 ,
         \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 ,
         \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 ,
         \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 ,
         \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 ,
         \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 ,
         \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 ,
         \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 ,
         \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 ,
         \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 ,
         \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 ,
         \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 ,
         \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 ,
         \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 ,
         \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 ,
         \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 ,
         \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 ,
         \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 ,
         \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 ,
         \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 ,
         \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 ,
         \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 ,
         \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 ,
         \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 ,
         \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 ,
         \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 ,
         \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 ,
         \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 ,
         \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 ,
         \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 ,
         \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 ,
         \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 ,
         \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 ,
         \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 ,
         \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 ,
         \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 ,
         \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 ,
         \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 ,
         \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 ,
         \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 ,
         \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 ,
         \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 ,
         \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 ,
         \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 ,
         \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 ,
         \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 ,
         \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 ,
         \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 ,
         \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 ,
         \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 ,
         \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 ,
         \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 ,
         \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 ,
         \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 ,
         \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 ,
         \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 ,
         \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 ,
         \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 ,
         \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 ,
         \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 ,
         \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 ,
         \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 ,
         \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 ,
         \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 ,
         \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 ,
         \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 ,
         \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 ,
         \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 ,
         \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 ,
         \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 ,
         \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 ,
         \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 ,
         \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 ,
         \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 ,
         \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 ,
         \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 ,
         \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 ,
         \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 ,
         \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 ,
         \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 ,
         \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 ,
         \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 ,
         \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 ,
         \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 ,
         \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 ,
         \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 ,
         \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 ,
         \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 ,
         \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 ,
         \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 ,
         \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 ,
         \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 ,
         \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 ,
         \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 ,
         \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 ,
         \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 ,
         \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 ,
         \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 ,
         \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 ,
         \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 ,
         \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 ,
         \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 ,
         \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 ,
         \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 ,
         \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 ,
         \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 ,
         \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 ,
         \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 ,
         \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 ,
         \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 ,
         \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 ,
         \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 ,
         \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 ,
         \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 ,
         \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 ,
         \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 ,
         \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 ,
         \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 ,
         \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 ,
         \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 ,
         \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 ,
         \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 ,
         \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 ,
         \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 ,
         \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 ,
         \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 ,
         \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 ,
         \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 ,
         \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 ,
         \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 ,
         \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 ,
         \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 ,
         \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 ,
         \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 ,
         \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 ,
         \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 ,
         \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 ,
         \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 ,
         \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 ,
         \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 ,
         \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 ,
         \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 ,
         \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 ,
         \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 ,
         \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 ,
         \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 ,
         \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 ,
         \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 ,
         \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 ,
         \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 ,
         \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 ,
         \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 ,
         \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 ,
         \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 ,
         \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 ,
         \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 ,
         \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 ,
         \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 ,
         \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 ,
         \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 ,
         \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 ,
         \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 ,
         \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 ,
         \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 ,
         \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 ,
         \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 ,
         \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 ,
         \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 ,
         \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 ,
         \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 ,
         \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 ,
         \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 ,
         \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 ,
         \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 ,
         \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 ,
         \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 ,
         \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 ,
         \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 ,
         \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 ,
         \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 ,
         \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 ,
         \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 ,
         \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 ,
         \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 ,
         \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 ,
         \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 ,
         \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 ,
         \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 ,
         \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 ,
         \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 ,
         \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 ,
         \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 ,
         \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 ,
         \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 ,
         \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 ,
         \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 ,
         \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 ,
         \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 ,
         \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 ,
         \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 ,
         \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 ,
         \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 ,
         \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 ,
         \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 ,
         \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 ,
         \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 ,
         \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 ,
         \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 ,
         \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 ,
         \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 ,
         \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 ,
         \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 ,
         \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 ,
         \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 ,
         \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 ,
         \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 ,
         \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 ,
         \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 ,
         \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 ,
         \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 ,
         \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 ,
         \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 ,
         \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 ,
         \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 ,
         \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 ,
         \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 ,
         \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 ,
         \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 ,
         \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 ,
         \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 ,
         \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 ,
         \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 ,
         \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 ,
         \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 ,
         \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 ,
         \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 ,
         \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 ,
         \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 ,
         \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 ,
         \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 ,
         \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 ,
         \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 ,
         \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 ,
         \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 ,
         \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 ,
         \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 ,
         \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 ,
         \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 ,
         \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 ,
         \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 ,
         \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 ,
         \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 ,
         \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 ,
         \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 ,
         \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 ,
         \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 ,
         \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 ,
         \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 ,
         \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 ,
         \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 ,
         \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 ,
         \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 ,
         \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 ,
         \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 ,
         \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 ,
         \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 ,
         \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 ,
         \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 ,
         \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 ,
         \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 ,
         \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 ,
         \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 ,
         \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 ,
         \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 ,
         \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 ,
         \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 ,
         \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 ,
         \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 ,
         \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 ,
         \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 ,
         \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 ,
         \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 ,
         \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 ,
         \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 ,
         \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 ,
         \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 ,
         \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 ,
         \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 ,
         \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 ,
         \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 ,
         \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 ,
         \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 ,
         \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 ,
         \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 ,
         \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 ,
         \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 ,
         \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 ,
         \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 ,
         \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 ,
         \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 ,
         \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 ,
         \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 ,
         \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 ,
         \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 ,
         \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 ,
         \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 ,
         \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 ,
         \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 ,
         \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 ,
         \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 ,
         \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 ,
         \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 ,
         \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 ,
         \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 ,
         \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 ,
         \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 ,
         \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 ,
         \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 ,
         \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 ,
         \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 ,
         \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 ,
         \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 ,
         \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 ,
         \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 ,
         \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 ,
         \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 ,
         \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 ,
         \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 ,
         \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 ,
         \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 ,
         \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 ,
         \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 ,
         \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 ,
         \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 ,
         \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 ,
         \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 ,
         \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 ,
         \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 ,
         \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 ,
         \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 ,
         \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 ,
         \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 ,
         \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 ,
         \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 ,
         \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 ,
         \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 ,
         \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 ,
         \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 ,
         \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 ,
         \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 ,
         \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 ,
         \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 ,
         \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 ,
         \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 ,
         \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 ,
         \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 ,
         \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 ,
         \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 ,
         \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 ,
         \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 ,
         \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 ,
         \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 ,
         \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 ,
         \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 ,
         \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 ,
         \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 ,
         \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 ,
         \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 ,
         \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 ,
         \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 ,
         \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 ,
         \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 ,
         \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 ,
         \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 ,
         \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 ,
         \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 ,
         \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 ,
         \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 ,
         \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 ,
         \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 ,
         \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 ,
         \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 ,
         \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 ,
         \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 ,
         \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 ,
         \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 ,
         \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 ,
         \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 ,
         \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 ,
         \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 ,
         \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 ,
         \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 ,
         \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 ,
         \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 ,
         \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 ,
         \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 ,
         \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 ,
         \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 ,
         \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 ,
         \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 ,
         \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 ,
         \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 ,
         \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 ,
         \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 ,
         \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 ,
         \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 ,
         \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 ,
         \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 ,
         \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 ,
         \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 ,
         \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 ,
         \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 ,
         \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 ,
         \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 ,
         \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 ,
         \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 ,
         \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 ,
         \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 ,
         \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 ,
         \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 ,
         \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 ,
         \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 ,
         \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 ,
         \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 ,
         \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 ,
         \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 ,
         \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 ,
         \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 ,
         \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 ,
         \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 ,
         \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 ,
         \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 ,
         \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 ,
         \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 ,
         \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 ,
         \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 ,
         \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 ,
         \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 ,
         \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 ,
         \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 ,
         \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 ,
         \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 ,
         \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 ,
         \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 ,
         \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 ,
         \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 ,
         \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 ,
         \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 ,
         \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 ,
         \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 ,
         \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 ,
         \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 ,
         \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 ,
         \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 ,
         \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 ,
         \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 ,
         \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 ,
         \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 ,
         \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 ,
         \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 ,
         \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 ,
         \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 ,
         \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 ,
         \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 ,
         \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 ,
         \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 ,
         \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 ,
         \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 ,
         \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 ,
         \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 ,
         \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 ,
         \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 ,
         \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 ,
         \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 ,
         \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 ,
         \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 ,
         \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 ,
         \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 ,
         \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 ,
         \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 ,
         \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 ,
         \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 ,
         \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 ,
         \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 ,
         \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 ,
         \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 ,
         \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 ,
         \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 ,
         \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 ,
         \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 ,
         \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 ,
         \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 ,
         \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 ,
         \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 ,
         \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 ,
         \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 ,
         \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 ,
         \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 ,
         \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 ,
         \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 ,
         \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 ,
         \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 ,
         \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 ,
         \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 ,
         \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 ,
         \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 ,
         \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 ,
         \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 ,
         \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 ,
         \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 ,
         \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 ,
         \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 ,
         \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 ,
         \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 ,
         \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 ,
         \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 ,
         \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 ,
         \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 ,
         \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 ,
         \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 ,
         \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 ,
         \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 ,
         \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 ,
         \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 ,
         \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 ,
         \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 ,
         \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 ,
         \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 ,
         \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 ,
         \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 ,
         \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 ,
         \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 ,
         \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 ,
         \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 ,
         \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 ,
         \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 ,
         \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 ,
         \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 ,
         \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 ,
         \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 ,
         \7861 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 ,
         \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 ,
         \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 ,
         \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 ,
         \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 ,
         \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 ,
         \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 ,
         \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 ,
         \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 ,
         \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 ,
         \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 ,
         \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 ,
         \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 ,
         \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 ,
         \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 ,
         \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 ,
         \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 ,
         \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 ,
         \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 ,
         \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 ,
         \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 ,
         \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 ,
         \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 ,
         \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 ,
         \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 ,
         \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 ,
         \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 ,
         \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 ,
         \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 ,
         \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 ,
         \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 ,
         \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 ,
         \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 ,
         \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 ,
         \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 ,
         \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 ,
         \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 ,
         \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 ,
         \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 ,
         \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 ,
         \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 ,
         \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 ,
         \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 ,
         \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 ,
         \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 ,
         \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 ,
         \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 ,
         \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 ,
         \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 ,
         \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 ,
         \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 ,
         \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 ,
         \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 ,
         \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 ,
         \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 ,
         \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 ,
         \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 ,
         \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 ,
         \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 ,
         \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 ,
         \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 ,
         \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 ,
         \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 ,
         \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 ,
         \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 ,
         \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 ,
         \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 ,
         \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 ,
         \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 ,
         \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 ,
         \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 ,
         \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 ,
         \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 ,
         \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 ,
         \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 ,
         \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 ,
         \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 ,
         \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 ,
         \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 ,
         \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 ,
         \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 ,
         \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 ,
         \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 ,
         \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 ,
         \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 ,
         \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 ,
         \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 ,
         \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 ,
         \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 ,
         \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 ,
         \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 ,
         \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 ,
         \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 ,
         \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 ,
         \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 ,
         \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 ,
         \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 ,
         \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 ,
         \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 ,
         \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 ,
         \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 ,
         \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 ,
         \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 ,
         \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 ,
         \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 ,
         \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 ,
         \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 ,
         \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 ,
         \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 ,
         \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 ,
         \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 ,
         \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 ,
         \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 ,
         \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 ,
         \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 ,
         \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 ,
         \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 ,
         \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 ,
         \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 ,
         \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 ,
         \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 ,
         \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 ,
         \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 ,
         \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 ,
         \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 ,
         \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 ,
         \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 ,
         \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 ,
         \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 ,
         \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 ,
         \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 ,
         \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 ,
         \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 ,
         \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 ,
         \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 ,
         \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 ,
         \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 ,
         \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 ,
         \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 ,
         \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 ,
         \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 ,
         \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 ,
         \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 ,
         \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 ,
         \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 ,
         \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 ,
         \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 ,
         \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 ,
         \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 ,
         \9351 , \9352 , \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 ,
         \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 ,
         \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 ,
         \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 ,
         \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 ,
         \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 ,
         \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 ,
         \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 ,
         \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 ,
         \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 ,
         \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 ,
         \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 ,
         \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 ,
         \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 ,
         \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 ,
         \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 ,
         \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 ,
         \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 ,
         \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 ,
         \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 ,
         \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 ,
         \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 ,
         \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 ,
         \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 ,
         \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 ,
         \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 ,
         \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 ,
         \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 ,
         \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 ,
         \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 ,
         \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 ,
         \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 ,
         \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 ,
         \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 ,
         \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 ,
         \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 ,
         \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 ,
         \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 ,
         \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 ,
         \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 ,
         \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 ,
         \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 ,
         \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 ,
         \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 ,
         \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 ,
         \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 ,
         \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 ,
         \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 ,
         \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 ,
         \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 ,
         \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 ,
         \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 ,
         \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 ,
         \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 ,
         \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 ,
         \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 ,
         \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 ,
         \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 ,
         \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 ,
         \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 ,
         \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 ,
         \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 ,
         \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 ,
         \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 ,
         \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 ,
         \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 ,
         \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 ,
         \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 ,
         \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 ,
         \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 ,
         \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 ,
         \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 ,
         \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 ,
         \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 ,
         \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 ,
         \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 ,
         \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 ,
         \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 ,
         \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 ,
         \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 ,
         \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 ,
         \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 ,
         \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 ,
         \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 ,
         \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 ,
         \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 ,
         \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 ,
         \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 ,
         \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 ,
         \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 ,
         \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 ,
         \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 ,
         \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 ,
         \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 ,
         \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 ,
         \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 ,
         \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 ,
         \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 ,
         \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 ,
         \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 ,
         \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 ,
         \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 ,
         \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 ,
         \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 ,
         \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 ,
         \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 ,
         \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 ,
         \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 ,
         \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 ,
         \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 ,
         \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 ,
         \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 ,
         \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 ,
         \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 ,
         \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 ,
         \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 ,
         \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 ,
         \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 ,
         \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 ,
         \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 ,
         \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 ,
         \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 ,
         \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 ,
         \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 ,
         \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 ,
         \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 ,
         \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 ,
         \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 ,
         \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 ,
         \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 ,
         \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 ,
         \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 ,
         \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 ,
         \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 ,
         \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 ,
         \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 ,
         \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 ,
         \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 ,
         \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 ,
         \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 ,
         \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 ,
         \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 ,
         \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 ,
         \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 ,
         \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 ,
         \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 ,
         \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 ,
         \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 ,
         \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 ,
         \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 ,
         \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 ,
         \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 ,
         \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 ,
         \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 ,
         \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 ,
         \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 ,
         \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 ,
         \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 ,
         \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 ,
         \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 ,
         \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 ,
         \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 ,
         \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 ,
         \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 ,
         \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 ,
         \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 ,
         \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 ,
         \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 ,
         \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 ,
         \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 ,
         \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 ,
         \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 ,
         \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 ,
         \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 ,
         \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 ,
         \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 ,
         \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 ,
         \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 ,
         \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 ,
         \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 ,
         \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 ,
         \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 ,
         \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 ,
         \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 ,
         \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 ,
         \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 ,
         \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 ,
         \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 ,
         \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 ,
         \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 ,
         \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 ,
         \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 ,
         \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 ,
         \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 ,
         \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 ,
         \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 ,
         \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 ,
         \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 ,
         \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 ,
         \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 ,
         \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 ,
         \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 ,
         \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 ,
         \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 ,
         \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 ,
         \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 ,
         \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 ,
         \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 ,
         \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 ,
         \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 ,
         \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 ,
         \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 ,
         \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 ,
         \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 ,
         \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 ,
         \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 ,
         \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 ,
         \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 ,
         \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 ,
         \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 ,
         \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 ,
         \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 ,
         \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 ,
         \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 ,
         \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 ,
         \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 ,
         \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 ,
         \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 ,
         \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 ,
         \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 ,
         \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 ,
         \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 ,
         \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 ,
         \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 ,
         \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 ,
         \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 ,
         \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 ,
         \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 ,
         \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 ,
         \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 ,
         \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 ,
         \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 ,
         \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 ,
         \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 ,
         \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 ,
         \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 ,
         \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 ,
         \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 ,
         \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 ,
         \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 ,
         \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 ,
         \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 ,
         \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 ,
         \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 ,
         \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 ,
         \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 ,
         \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 ,
         \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 ,
         \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 ,
         \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 ,
         \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 ,
         \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 ,
         \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 ,
         \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 ,
         \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 ,
         \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 ,
         \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 ,
         \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 ,
         \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 ,
         \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 ,
         \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 ,
         \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 ,
         \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 ,
         \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 ,
         \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 ,
         \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 ,
         \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 ,
         \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 ,
         \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 ,
         \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 ,
         \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 ,
         \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 ,
         \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 ,
         \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 ,
         \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 ,
         \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 ,
         \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 ,
         \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 ,
         \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 ,
         \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 ,
         \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 ,
         \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 ,
         \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 ,
         \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 ,
         \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 ,
         \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 ,
         \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 ,
         \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 ,
         \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 ,
         \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 ,
         \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 ,
         \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 ,
         \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 ,
         \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 ,
         \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 ,
         \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 ,
         \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 ,
         \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 ,
         \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 ,
         \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 ,
         \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 ,
         \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 ,
         \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 ,
         \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 ,
         \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 ,
         \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 ,
         \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 ,
         \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 ,
         \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 ,
         \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 ,
         \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 ,
         \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 ,
         \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 ,
         \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 ,
         \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 ,
         \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 ,
         \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 ,
         \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 ,
         \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 ,
         \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 ,
         \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 ,
         \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 ,
         \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 ,
         \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 ,
         \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 ,
         \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 ,
         \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 ,
         \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 ,
         \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 ,
         \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 ,
         \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 ,
         \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 ,
         \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 ,
         \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 ,
         \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 ,
         \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 ,
         \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 ,
         \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 ,
         \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 ,
         \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 ,
         \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 ,
         \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 ,
         \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 ,
         \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 ,
         \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 ,
         \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 ,
         \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 ,
         \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 ,
         \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 ,
         \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 ,
         \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 ,
         \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 ,
         \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 ,
         \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 ,
         \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 ,
         \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 ,
         \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 ,
         \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 ,
         \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 ,
         \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 ,
         \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 ,
         \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 ,
         \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 ,
         \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 ,
         \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 ,
         \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 ,
         \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 ,
         \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 ,
         \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 ,
         \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 ,
         \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 ,
         \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 ,
         \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 ,
         \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 ,
         \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 ,
         \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 ,
         \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 ,
         \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 ,
         \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 ,
         \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 ,
         \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 ,
         \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 ,
         \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 ,
         \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 ,
         \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 ,
         \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 ,
         \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 ,
         \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 ,
         \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 ,
         \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 ,
         \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 ,
         \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 ,
         \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 ,
         \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 ,
         \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 ,
         \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 ,
         \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 ,
         \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 ,
         \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 ,
         \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 ,
         \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 ,
         \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 ,
         \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 ,
         \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 ,
         \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 ,
         \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 ,
         \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 ,
         \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 ,
         \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 ,
         \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 ,
         \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 ,
         \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 ,
         \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 ,
         \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 ,
         \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 ,
         \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 ,
         \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 ,
         \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 ,
         \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 ,
         \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 ,
         \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 ,
         \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 ,
         \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 ,
         \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 ,
         \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 ,
         \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 ,
         \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 ,
         \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 ,
         \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 ,
         \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 ,
         \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 ,
         \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 ,
         \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 ,
         \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 ,
         \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 ,
         \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 ,
         \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 ,
         \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 ,
         \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 ,
         \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 ,
         \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 ,
         \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 ,
         \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 ,
         \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 ,
         \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 ,
         \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 ,
         \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 ,
         \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 ,
         \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 ,
         \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 ,
         \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 ,
         \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 ,
         \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 ,
         \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 ,
         \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 ,
         \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 ,
         \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 ,
         \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 ,
         \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 ,
         \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 ,
         \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 ,
         \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 ,
         \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 ,
         \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 ,
         \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 ,
         \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 ,
         \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 ,
         \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 ,
         \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 ,
         \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 ,
         \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 ,
         \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 ,
         \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 ,
         \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 ,
         \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 ,
         \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 ,
         \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 ,
         \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 ,
         \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 ,
         \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 ,
         \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 ,
         \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 ,
         \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 ,
         \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 ,
         \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 ,
         \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 ,
         \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 ,
         \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 ,
         \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 ,
         \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 ,
         \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 ,
         \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 ,
         \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 ,
         \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 ,
         \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 ,
         \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 ,
         \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 ,
         \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 ,
         \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 ,
         \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 ,
         \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 ,
         \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 ,
         \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 ,
         \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 ,
         \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 ,
         \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 ,
         \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 ,
         \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 ,
         \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 ,
         \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 ,
         \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 ,
         \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 ,
         \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 ,
         \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 ,
         \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 ,
         \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 ,
         \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 ,
         \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 ,
         \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 ,
         \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 ,
         \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 ,
         \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 ,
         \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 ,
         \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 ,
         \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 ,
         \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 ,
         \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 ,
         \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 ,
         \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 ,
         \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 ,
         \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 ,
         \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 ,
         \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 ,
         \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 ,
         \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 ,
         \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 ,
         \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 ,
         \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 ,
         \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 ,
         \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 ,
         \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 ,
         \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 ,
         \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 ,
         \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 ,
         \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 ,
         \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 ,
         \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 ,
         \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 ,
         \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 ,
         \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 ,
         \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 ,
         \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 ,
         \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 ,
         \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 ,
         \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 ,
         \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 ,
         \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 ,
         \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 ,
         \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 ,
         \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 ,
         \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 ,
         \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 ,
         \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 ,
         \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 ,
         \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 ,
         \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 ,
         \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 ,
         \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 ,
         \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 ,
         \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 ,
         \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 ,
         \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 ,
         \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 ,
         \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 ,
         \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 ,
         \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 ,
         \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 ,
         \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 ,
         \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 ,
         \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 ,
         \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 ,
         \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 ,
         \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 ,
         \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 ,
         \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 ,
         \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 ,
         \15311 , \15312 , \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 ,
         \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 ,
         \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 ,
         \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 ,
         \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 ,
         \15361 , \15362 , \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 ,
         \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 ,
         \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 ,
         \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 ,
         \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 ,
         \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 ,
         \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 ,
         \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 ,
         \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 ,
         \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 ,
         \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 ,
         \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 ,
         \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 ,
         \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 ,
         \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 ,
         \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 ,
         \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 ,
         \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 ,
         \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 ,
         \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 ,
         \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 ,
         \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 ,
         \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 ,
         \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 ,
         \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 ,
         \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 ,
         \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 ,
         \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 ,
         \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 ,
         \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 ,
         \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 ,
         \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 ,
         \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 ,
         \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 ,
         \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 ,
         \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 ,
         \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 ,
         \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 ,
         \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 ,
         \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 ,
         \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 ,
         \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 ,
         \15781 , \15782 , \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 ,
         \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 ,
         \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 ,
         \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 ,
         \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 ,
         \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 ,
         \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 ,
         \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 ,
         \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 ,
         \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 ,
         \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 ,
         \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 ,
         \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 ,
         \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 ,
         \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 ,
         \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 ,
         \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 ,
         \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 ,
         \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 ,
         \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 ,
         \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 ,
         \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 ,
         \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 ,
         \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 ,
         \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 ,
         \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 ,
         \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 ,
         \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 ,
         \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 ,
         \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 ,
         \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 ,
         \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 ,
         \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 ,
         \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 ,
         \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 ,
         \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 ,
         \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 ,
         \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 ,
         \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 ,
         \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 ,
         \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 ,
         \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 ,
         \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 ,
         \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 ,
         \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 ,
         \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 ,
         \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 ,
         \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 ,
         \16261 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 ,
         \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 ,
         \16281 , \16282 , \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 ,
         \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 ,
         \16301 , \16302 , \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 ,
         \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 ,
         \16321 , \16322 , \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 ,
         \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 ,
         \16341 , \16342 , \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 ,
         \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 ,
         \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 ,
         \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 ,
         \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 ,
         \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 ,
         \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 ,
         \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 ,
         \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 ,
         \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 ,
         \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 ,
         \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 ,
         \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 ,
         \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 ,
         \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 ,
         \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 ,
         \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 ,
         \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 ,
         \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 ,
         \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 ,
         \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 ,
         \16551 , \16552 , \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 ,
         \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 ,
         \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 ,
         \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 ,
         \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 ,
         \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 ,
         \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 ,
         \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 ,
         \16631 , \16632 , \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 ,
         \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 ,
         \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 ,
         \16661 , \16662 , \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 ,
         \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 ,
         \16681 , \16682 , \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 ,
         \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 ,
         \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 ,
         \16711 , \16712 , \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 ,
         \16721 , \16722 , \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 ,
         \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 ,
         \16741 , \16742 , \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 ,
         \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 ,
         \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 ,
         \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 ,
         \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 ,
         \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 ,
         \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 ,
         \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 ,
         \16821 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 ,
         \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 ,
         \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 ,
         \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 ,
         \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 ,
         \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 ,
         \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 ,
         \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 ,
         \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 ,
         \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 ,
         \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 ,
         \16931 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 ,
         \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 ,
         \16951 , \16952 , \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 ,
         \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 ,
         \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 ,
         \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 ,
         \16991 , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 ,
         \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 ,
         \17011 , \17012 , \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 ,
         \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 ,
         \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 ,
         \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 ,
         \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 ,
         \17061 , \17062 , \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 ,
         \17071 , \17072 , \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 ,
         \17081 , \17082 , \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 ,
         \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 ,
         \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 ,
         \17111 , \17112 , \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 ,
         \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 ,
         \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 ,
         \17141 , \17142 , \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 ,
         \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 ,
         \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 ,
         \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 ,
         \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 ,
         \17191 , \17192 , \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 ,
         \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 ,
         \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 ,
         \17221 , \17222 , \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 ,
         \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 ,
         \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 ,
         \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 ,
         \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 ,
         \17271 , \17272 , \17273 , \17274 , \17275 , \17276 , \17277 , \17278 , \17279 , \17280 ,
         \17281 , \17282 , \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 ,
         \17291 , \17292 , \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 ,
         \17301 , \17302 , \17303 , \17304 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 ,
         \17311 , \17312 , \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 ,
         \17321 , \17322 , \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 , \17330 ,
         \17331 , \17332 , \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 ,
         \17341 , \17342 , \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 ,
         \17351 , \17352 , \17353 , \17354 , \17355 , \17356 , \17357 , \17358 , \17359 , \17360 ,
         \17361 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 ,
         \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 ,
         \17381 , \17382 , \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 ,
         \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 ,
         \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 ,
         \17411 , \17412 , \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 ,
         \17421 , \17422 , \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 ,
         \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 ,
         \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 ,
         \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 ,
         \17461 , \17462 , \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 ,
         \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 ,
         \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 ,
         \17491 , \17492 , \17493 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 ,
         \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 ,
         \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 ,
         \17521 , \17522 , \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 ,
         \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 ,
         \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 ,
         \17551 , \17552 , \17553 , \17554 , \17555 , \17556 , \17557 , \17558 , \17559 , \17560 ,
         \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 ,
         \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 ,
         \17581 , \17582 , \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 ,
         \17591 , \17592 , \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 ,
         \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 ,
         \17611 , \17612 , \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 ,
         \17621 , \17622 , \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 ,
         \17631 , \17632 , \17633 , \17634 , \17635 , \17636 , \17637 , \17638 , \17639 , \17640 ,
         \17641 , \17642 , \17643 , \17644 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 ,
         \17651 , \17652 , \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 ,
         \17661 , \17662 , \17663 , \17664 , \17665 , \17666 , \17667 , \17668 , \17669 , \17670 ,
         \17671 , \17672 , \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 ,
         \17681 , \17682 , \17683 , \17684 , \17685 , \17686 , \17687 , \17688 , \17689 , \17690 ,
         \17691 , \17692 , \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 ,
         \17701 , \17702 , \17703 , \17704 , \17705 , \17706 , \17707 , \17708 , \17709 , \17710 ,
         \17711 , \17712 , \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 ,
         \17721 , \17722 , \17723 , \17724 , \17725 , \17726 , \17727 , \17728 , \17729 , \17730 ,
         \17731 , \17732 , \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 ,
         \17741 , \17742 , \17743 , \17744 , \17745 , \17746 , \17747 , \17748 , \17749 , \17750 ,
         \17751 , \17752 , \17753 , \17754 , \17755 , \17756 , \17757 , \17758 , \17759 , \17760 ,
         \17761 , \17762 , \17763 , \17764 , \17765 , \17766 , \17767 , \17768 , \17769 , \17770 ,
         \17771 , \17772 , \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 ,
         \17781 , \17782 , \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 ,
         \17791 , \17792 , \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 ,
         \17801 , \17802 , \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 ,
         \17811 , \17812 , \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 ,
         \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 ,
         \17831 , \17832 , \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 ,
         \17841 , \17842 , \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 ,
         \17851 , \17852 , \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 ,
         \17861 , \17862 , \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 ,
         \17871 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 ,
         \17881 , \17882 , \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 ,
         \17891 , \17892 , \17893 , \17894 , \17895 , \17896 , \17897 , \17898 , \17899 , \17900 ,
         \17901 , \17902 , \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 ,
         \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 ,
         \17921 , \17922 , \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 ,
         \17931 , \17932 , \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 ,
         \17941 , \17942 , \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 ,
         \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 ,
         \17961 , \17962 , \17963 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 ,
         \17971 , \17972 , \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 ,
         \17981 , \17982 , \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 ,
         \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 ,
         \18001 , \18002 , \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 ,
         \18011 , \18012 , \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 ,
         \18021 , \18022 , \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 ,
         \18031 , \18032 , \18033 , \18034 , \18035 , \18036 , \18037 , \18038 , \18039 , \18040 ,
         \18041 , \18042 , \18043 , \18044 , \18045 , \18046 , \18047 , \18048 , \18049 , \18050 ,
         \18051 , \18052 , \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 ,
         \18061 , \18062 , \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 ,
         \18071 , \18072 , \18073 , \18074 , \18075 , \18076 , \18077 , \18078 , \18079 , \18080 ,
         \18081 , \18082 , \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 ,
         \18091 , \18092 , \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 ,
         \18101 , \18102 , \18103 , \18104 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 ,
         \18111 , \18112 , \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 ,
         \18121 , \18122 , \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 , \18130 ,
         \18131 , \18132 , \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 ,
         \18141 , \18142 , \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 ,
         \18151 , \18152 , \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 ,
         \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 ,
         \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 ,
         \18181 , \18182 , \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 ,
         \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 ,
         \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 ,
         \18211 , \18212 , \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 ,
         \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 ,
         \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 ,
         \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 ,
         \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 ,
         \18261 , \18262 , \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 ,
         \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 ,
         \18281 , \18282 , \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 ,
         \18291 , \18292 , \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 ,
         \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 ,
         \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 ,
         \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 ,
         \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 ,
         \18341 , \18342 , \18343 , \18344 , \18345 , \18346 , \18347 , \18348 , \18349 , \18350 ,
         \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 ,
         \18361 , \18362 , \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 ,
         \18371 , \18372 , \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 ,
         \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 ,
         \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 ,
         \18401 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 ,
         \18411 , \18412 , \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 ,
         \18421 , \18422 , \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 ,
         \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 ,
         \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 ,
         \18451 , \18452 , \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 ,
         \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 ,
         \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 ,
         \18481 , \18482 , \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 ,
         \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 ,
         \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 ,
         \18511 , \18512 , \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 ,
         \18521 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 ,
         \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 ,
         \18541 , \18542 , \18543 , \18544 , \18545 , \18546 , \18547 , \18548 , \18549 , \18550 ,
         \18551 , \18552 , \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 ,
         \18561 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 ,
         \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 ,
         \18581 , \18582 , \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 ,
         \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 ,
         \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 ,
         \18611 , \18612 , \18613 , \18614 , \18615 , \18616 , \18617 , \18618 , \18619 , \18620 ,
         \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 ,
         \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 ,
         \18641 , \18642 , \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 ,
         \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 ,
         \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 ,
         \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 ,
         \18681 , \18682 , \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 ,
         \18691 , \18692 , \18693 , \18694 , \18695 , \18696 , \18697 , \18698 , \18699 , \18700 ,
         \18701 , \18702 , \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 ,
         \18711 , \18712 , \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 ,
         \18721 , \18722 , \18723 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 ,
         \18731 , \18732 , \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 ,
         \18741 , \18742 , \18743 , \18744 , \18745 , \18746 , \18747 , \18748 , \18749 , \18750 ,
         \18751 , \18752 , \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 ,
         \18761 , \18762 , \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 ,
         \18771 , \18772 , \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 ,
         \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 ,
         \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 ,
         \18801 , \18802 , \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 ,
         \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 ,
         \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 ,
         \18831 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 ,
         \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 ,
         \18851 , \18852 , \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 ,
         \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 ,
         \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 ,
         \18881 , \18882 , \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 ,
         \18891 , \18892 , \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 ,
         \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 ,
         \18911 , \18912 , \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 ,
         \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 ,
         \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 ,
         \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 ,
         \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 ,
         \18961 , \18962 , \18963 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 ,
         \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 ,
         \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 ,
         \18991 , \18992 , \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 ,
         \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 ,
         \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 ,
         \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 , \19028 , \19029 , \19030 ,
         \19031 , \19032 , \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 ,
         \19041 , \19042 , \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 ,
         \19051 , \19052 , \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19059 , \19060 ,
         \19061 , \19062 , \19063 , \19064 , \19065 , \19066 , \19067 , \19068 , \19069 , \19070 ,
         \19071 , \19072 , \19073 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 ,
         \19081 , \19082 , \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 , \19090 ,
         \19091 , \19092 , \19093 , \19094 , \19095 , \19096 , \19097 , \19098 , \19099 , \19100 ,
         \19101 , \19102 , \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 ,
         \19111 , \19112 , \19113 , \19114 , \19115 , \19116 , \19117 , \19118 , \19119 , \19120 ,
         \19121 , \19122 , \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 ,
         \19131 , \19132 , \19133 , \19134 , \19135 , \19136 , \19137 , \19138 , \19139 , \19140 ,
         \19141 , \19142 , \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 ,
         \19151 , \19152 , \19153 , \19154 , \19155 , \19156 , \19157 , \19158 , \19159 , \19160 ,
         \19161 , \19162 , \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 ,
         \19171 , \19172 , \19173 , \19174 , \19175 , \19176 , \19177 , \19178 , \19179 , \19180 ,
         \19181 , \19182 , \19183 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 ,
         \19191 , \19192 , \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 , \19200 ,
         \19201 , \19202 , \19203 , \19204 , \19205 , \19206 , \19207 , \19208 , \19209 , \19210 ,
         \19211 , \19212 , \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 ,
         \19221 , \19222 , \19223 , \19224 , \19225 , \19226 , \19227 , \19228 , \19229 , \19230 ,
         \19231 , \19232 , \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 ,
         \19241 , \19242 , \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 ,
         \19251 , \19252 , \19253 , \19254 , \19255 , \19256 , \19257 , \19258 , \19259 , \19260 ,
         \19261 , \19262 , \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 ,
         \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 ,
         \19281 , \19282 , \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 ,
         \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 ,
         \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 ,
         \19311 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 ,
         \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 ,
         \19331 , \19332 , \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 ,
         \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 ,
         \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 ,
         \19361 , \19362 , \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 ,
         \19371 , \19372 , \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 ,
         \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 ,
         \19391 , \19392 , \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 ,
         \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 ,
         \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 ,
         \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 ,
         \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 ,
         \19441 , \19442 , \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 ,
         \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 ,
         \19461 , \19462 , \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 ,
         \19471 , \19472 , \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 ,
         \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 ,
         \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 ,
         \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 ,
         \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 ,
         \19521 , \19522 , \19523 , \19524 , \19525 , \19526 , \19527 , \19528 , \19529 , \19530 ,
         \19531 , \19532 , \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 ,
         \19541 , \19542 , \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 ,
         \19551 , \19552 , \19553 , \19554 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 ,
         \19561 , \19562 , \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 ,
         \19571 , \19572 , \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 , \19580 ,
         \19581 , \19582 , \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 ,
         \19591 , \19592 , \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 ,
         \19601 , \19602 , \19603 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 ,
         \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 ,
         \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 ,
         \19631 , \19632 , \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 ,
         \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 ,
         \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 ,
         \19661 , \19662 , \19663 , \19664 , \19665 , \19666 , \19667 , \19668 , \19669 , \19670 ,
         \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 ,
         \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 ,
         \19691 , \19692 , \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 ,
         \19701 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 ,
         \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 ,
         \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 ,
         \19731 , \19732 , \19733 , \19734 , \19735 , \19736 , \19737 , \19738 , \19739 , \19740 ,
         \19741 , \19742 , \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 ,
         \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 ,
         \19761 , \19762 , \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 ,
         \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 ,
         \19781 , \19782 , \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 ,
         \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 ,
         \19801 , \19802 , \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 ,
         \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 ,
         \19821 , \19822 , \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 ,
         \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 ,
         \19841 , \19842 , \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 ,
         \19851 , \19852 , \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 ,
         \19861 , \19862 , \19863 , \19864 , \19865 , \19866 , \19867 , \19868 , \19869 , \19870 ,
         \19871 , \19872 , \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 ,
         \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 ,
         \19891 , \19892 , \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 ,
         \19901 , \19902 , \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 ,
         \19911 , \19912 , \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 ,
         \19921 , \19922 , \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 ,
         \19931 , \19932 , \19933 , \19934 , \19935 , \19936 , \19937 , \19938 , \19939 , \19940 ,
         \19941 , \19942 , \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 ,
         \19951 , \19952 , \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 ,
         \19961 , \19962 , \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 ,
         \19971 , \19972 , \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 ,
         \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 ,
         \19991 , \19992 , \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 ,
         \20001 , \20002 , \20003 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 ,
         \20011 , \20012 , \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 ,
         \20021 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 ,
         \20031 , \20032 , \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 ,
         \20041 , \20042 , \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 ,
         \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 ,
         \20061 , \20062 , \20063 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 ,
         \20071 , \20072 , \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 ,
         \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 ,
         \20091 , \20092 , \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 ,
         \20101 , \20102 , \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 ,
         \20111 , \20112 , \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 ,
         \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 ,
         \20131 , \20132 , \20133 , \20134 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 ,
         \20141 , \20142 , \20143 , \20144 , \20145 , \20146 , \20147 , \20148 , \20149 , \20150 ,
         \20151 , \20152 , \20153 , \20154 , \20155 , \20156 , \20157 , \20158 , \20159 , \20160 ,
         \20161 , \20162 , \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 ,
         \20171 , \20172 , \20173 , \20174 , \20175 , \20176 , \20177 , \20178 , \20179 , \20180 ,
         \20181 , \20182 , \20183 , \20184 , \20185 , \20186 , \20187 , \20188 , \20189 , \20190 ,
         \20191 , \20192 , \20193 , \20194 , \20195 , \20196 , \20197 , \20198 , \20199 , \20200 ,
         \20201 , \20202 , \20203 , \20204 , \20205 , \20206 , \20207 , \20208 , \20209 , \20210 ,
         \20211 , \20212 , \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 ,
         \20221 , \20222 , \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 ,
         \20231 , \20232 , \20233 , \20234 , \20235 , \20236 , \20237 , \20238 , \20239 , \20240 ,
         \20241 , \20242 , \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 ,
         \20251 , \20252 , \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 ,
         \20261 , \20262 , \20263 , \20264 , \20265 , \20266 , \20267 , \20268 , \20269 , \20270 ,
         \20271 , \20272 , \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 ,
         \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 ,
         \20291 , \20292 , \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 ,
         \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 ,
         \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 ,
         \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 ,
         \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 ,
         \20341 , \20342 , \20343 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 ,
         \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 ,
         \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 ,
         \20371 , \20372 , \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 ,
         \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 ,
         \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 ,
         \20401 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 ,
         \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 ,
         \20421 , \20422 , \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 ,
         \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 ,
         \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 ,
         \20451 , \20452 , \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 ,
         \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 ,
         \20471 , \20472 , \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 ,
         \20481 , \20482 , \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 ,
         \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 ,
         \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 ,
         \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 ,
         \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 ,
         \20531 , \20532 , \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 , \20540 ,
         \20541 , \20542 , \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 ,
         \20551 , \20552 , \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 ,
         \20561 , \20562 , \20563 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 ,
         \20571 , \20572 , \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 ,
         \20581 , \20582 , \20583 , \20584 , \20585 , \20586 , \20587 , \20588 , \20589 , \20590 ,
         \20591 , \20592 , \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 ,
         \20601 , \20602 , \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 ,
         \20611 , \20612 , \20613 , \20614 , \20615 , \20616 , \20617 , \20618 , \20619 , \20620 ,
         \20621 , \20622 , \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 ,
         \20631 , \20632 , \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 ,
         \20641 , \20642 , \20643 , \20644 , \20645 , \20646 , \20647 , \20648 , \20649 , \20650 ,
         \20651 , \20652 , \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 ,
         \20661 , \20662 , \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 ,
         \20671 , \20672 , \20673 , \20674 , \20675 , \20676 , \20677 , \20678 , \20679 , \20680 ,
         \20681 , \20682 , \20683 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 ,
         \20691 , \20692 , \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 ,
         \20701 , \20702 , \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20710 ,
         \20711 , \20712 , \20713 , \20714 , \20715 , \20716 , \20717 , \20718 , \20719 , \20720 ,
         \20721 , \20722 , \20723 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 ,
         \20731 , \20732 , \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 ,
         \20741 , \20742 , \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 ,
         \20751 , \20752 , \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 ,
         \20761 , \20762 , \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 ,
         \20771 , \20772 , \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 ,
         \20781 , \20782 , \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 ,
         \20791 , \20792 , \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 ,
         \20801 , \20802 , \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 ,
         \20811 , \20812 , \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 ,
         \20821 , \20822 , \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 ,
         \20831 , \20832 , \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 ,
         \20841 , \20842 , \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 ,
         \20851 , \20852 , \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 ,
         \20861 , \20862 , \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 ,
         \20871 , \20872 , \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 ,
         \20881 , \20882 , \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 ,
         \20891 , \20892 , \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 ,
         \20901 , \20902 , \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 ,
         \20911 , \20912 , \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 ,
         \20921 , \20922 , \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 ,
         \20931 , \20932 , \20933 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 ,
         \20941 , \20942 , \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 ,
         \20951 , \20952 , \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 ,
         \20961 , \20962 , \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 ,
         \20971 , \20972 , \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 ,
         \20981 , \20982 , \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 ,
         \20991 , \20992 , \20993 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 ,
         \21001 , \21002 , \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 ,
         \21011 , \21012 , \21013 , \21014 , \21015 , \21016 , \21017 , \21018 , \21019 , \21020 ,
         \21021 , \21022 , \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 ,
         \21031 , \21032 , \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 ,
         \21041 , \21042 , \21043 , \21044 , \21045 , \21046 , \21047 , \21048 , \21049 , \21050 ,
         \21051 , \21052 , \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 ,
         \21061 , \21062 , \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 ,
         \21071 , \21072 , \21073 , \21074 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 ,
         \21081 , \21082 , \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 ,
         \21091 , \21092 , \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 , \21100 ,
         \21101 , \21102 , \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 ,
         \21111 , \21112 , \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 ,
         \21121 , \21122 , \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 ,
         \21131 , \21132 , \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 ,
         \21141 , \21142 , \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 ,
         \21151 , \21152 , \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 ,
         \21161 , \21162 , \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 ,
         \21171 , \21172 , \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 ,
         \21181 , \21182 , \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 ,
         \21191 , \21192 , \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 ,
         \21201 , \21202 , \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 ,
         \21211 , \21212 , \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 ,
         \21221 , \21222 , \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 ,
         \21231 , \21232 , \21233 , \21234 , \21235 , \21236 , \21237 , \21238 , \21239 , \21240 ,
         \21241 , \21242 , \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 ,
         \21251 , \21252 , \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 ,
         \21261 , \21262 , \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 ,
         \21271 , \21272 , \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 ,
         \21281 , \21282 , \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 ,
         \21291 , \21292 , \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 ,
         \21301 , \21302 , \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 ,
         \21311 , \21312 , \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 ,
         \21321 , \21322 , \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 ,
         \21331 , \21332 , \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 ,
         \21341 , \21342 , \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 ,
         \21351 , \21352 , \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 ,
         \21361 , \21362 , \21363 , \21364 , \21365 , \21366 , \21367 , \21368 , \21369 , \21370 ,
         \21371 , \21372 , \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 ,
         \21381 , \21382 , \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 ,
         \21391 , \21392 , \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 ,
         \21401 , \21402 , \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 ,
         \21411 , \21412 , \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 ,
         \21421 , \21422 , \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 ,
         \21431 , \21432 , \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 ,
         \21441 , \21442 , \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 ,
         \21451 , \21452 , \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 ,
         \21461 , \21462 , \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 ,
         \21471 , \21472 , \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 ,
         \21481 , \21482 , \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 ,
         \21491 , \21492 , \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 ,
         \21501 , \21502 , \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 ,
         \21511 , \21512 , \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 ,
         \21521 , \21522 , \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 ,
         \21531 , \21532 , \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 ,
         \21541 , \21542 , \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 ,
         \21551 , \21552 , \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 ,
         \21561 , \21562 , \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 ,
         \21571 , \21572 , \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 ,
         \21581 , \21582 , \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 ,
         \21591 , \21592 , \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 ,
         \21601 , \21602 , \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 ,
         \21611 , \21612 , \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 ,
         \21621 , \21622 , \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 ,
         \21631 , \21632 , \21633 , \21634 , \21635 , \21636 , \21637 , \21638 , \21639 , \21640 ,
         \21641 , \21642 , \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 ,
         \21651 , \21652 , \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 ,
         \21661 , \21662 , \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 ,
         \21671 , \21672 , \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 ,
         \21681 , \21682 , \21683 , \21684 , \21685 , \21686 , \21687 , \21688 , \21689 , \21690 ,
         \21691 , \21692 , \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 ,
         \21701 , \21702 , \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 ,
         \21711 , \21712 , \21713 , \21714 , \21715 , \21716 , \21717 , \21718 , \21719 , \21720 ,
         \21721 , \21722 , \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 ,
         \21731 , \21732 , \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 ,
         \21741 , \21742 , \21743 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 ,
         \21751 , \21752 , \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 ,
         \21761 , \21762 , \21763 , \21764 , \21765 , \21766 , \21767 , \21768 , \21769 , \21770 ,
         \21771 , \21772 , \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 ,
         \21781 , \21782 , \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 ,
         \21791 , \21792 , \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 ,
         \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 ,
         \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 ,
         \21821 , \21822 , \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 ,
         \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 ,
         \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 ,
         \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 ,
         \21861 , \21862 , \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 ,
         \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 ,
         \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 ,
         \21891 , \21892 , \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 ,
         \21901 , \21902 , \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 ,
         \21911 , \21912 , \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 ,
         \21921 , \21922 , \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 ,
         \21931 , \21932 , \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 ,
         \21941 , \21942 , \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 ,
         \21951 , \21952 , \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 ,
         \21961 , \21962 , \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 ,
         \21971 , \21972 , \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 ,
         \21981 , \21982 , \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 ,
         \21991 , \21992 , \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 ,
         \22001 , \22002 , \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 ,
         \22011 , \22012 , \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 ,
         \22021 , \22022 , \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 ,
         \22031 , \22032 , \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 ,
         \22041 , \22042 , \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 ,
         \22051 , \22052 , \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 ,
         \22061 , \22062 , \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 ,
         \22071 , \22072 , \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 ,
         \22081 , \22082 , \22083 , \22084 , \22085 , \22086 , \22087 , \22088 , \22089 , \22090 ,
         \22091 , \22092 , \22093 , \22094 , \22095 , \22096 , \22097 , \22098 , \22099 , \22100 ,
         \22101 , \22102 , \22103 , \22104 , \22105 , \22106 , \22107 , \22108 , \22109 , \22110 ,
         \22111 , \22112 , \22113 , \22114 , \22115 , \22116 , \22117 , \22118 , \22119 , \22120 ,
         \22121 , \22122 , \22123 , \22124 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 ,
         \22131 , \22132 , \22133 , \22134 , \22135 , \22136 , \22137 , \22138 , \22139 , \22140 ,
         \22141 , \22142 , \22143 , \22144 , \22145 , \22146 , \22147 , \22148 , \22149 , \22150 ,
         \22151 , \22152 , \22153 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 ,
         \22161 , \22162 , \22163 , \22164 , \22165 , \22166 , \22167 , \22168 , \22169 , \22170 ,
         \22171 , \22172 , \22173 , \22174 , \22175 , \22176 , \22177 , \22178 , \22179 , \22180 ,
         \22181 , \22182 , \22183 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 ,
         \22191 , \22192 , \22193 , \22194 , \22195 , \22196 , \22197 , \22198 , \22199 , \22200 ,
         \22201 , \22202 , \22203 , \22204 , \22205 , \22206 , \22207 , \22208 , \22209 , \22210 ,
         \22211 , \22212 , \22213 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 ,
         \22221 , \22222 , \22223 , \22224 , \22225 , \22226 , \22227 , \22228 , \22229 , \22230 ,
         \22231 , \22232 , \22233 , \22234 , \22235 , \22236 , \22237 , \22238 , \22239 , \22240 ,
         \22241 , \22242 , \22243 , \22244 , \22245 , \22246 , \22247 , \22248 , \22249 , \22250 ,
         \22251 , \22252 , \22253 , \22254 , \22255 , \22256 , \22257 , \22258 , \22259 , \22260 ,
         \22261 , \22262 , \22263 , \22264 , \22265 , \22266 , \22267 , \22268 , \22269 , \22270 ,
         \22271 , \22272 , \22273 , \22274 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 ,
         \22281 , \22282 , \22283 , \22284 , \22285 , \22286 , \22287 , \22288 , \22289 , \22290 ,
         \22291 , \22292 , \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , \22299 , \22300 ,
         \22301 , \22302 , \22303 , \22304 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 ,
         \22311 , \22312 , \22313 , \22314 , \22315 , \22316 , \22317 , \22318 , \22319 , \22320 ,
         \22321 , \22322 , \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , \22329 , \22330 ,
         \22331 , \22332 , \22333 , \22334 , \22335 , \22336 , \22337 , \22338 , \22339 , \22340 ,
         \22341 , \22342 , \22343 , \22344 , \22345 , \22346 , \22347 , \22348 , \22349 , \22350 ,
         \22351 , \22352 , \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , \22359 , \22360 ,
         \22361 , \22362 , \22363 , \22364 , \22365 , \22366 , \22367 , \22368 , \22369 , \22370 ,
         \22371 , \22372 , \22373 , \22374 , \22375 , \22376 , \22377 , \22378 , \22379 , \22380 ,
         \22381 , \22382 , \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 ,
         \22391 , \22392 , \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 ,
         \22401 , \22402 , \22403 , \22404 , \22405 , \22406 , \22407 , \22408 , \22409 , \22410 ,
         \22411 , \22412 , \22413 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 ,
         \22421 , \22422 , \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 ,
         \22431 , \22432 , \22433 , \22434 , \22435 , \22436 , \22437 , \22438 , \22439 , \22440 ,
         \22441 , \22442 , \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 ,
         \22451 , \22452 , \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 ,
         \22461 , \22462 , \22463 , \22464 , \22465 , \22466 , \22467 , \22468 , \22469 , \22470 ,
         \22471 , \22472 , \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 ,
         \22481 , \22482 , \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 ,
         \22491 , \22492 , \22493 , \22494 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 ,
         \22501 , \22502 , \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 ,
         \22511 , \22512 , \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 , \22520 ,
         \22521 , \22522 , \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 ,
         \22531 , \22532 , \22533 , \22534 , \22535 , \22536 , \22537 , \22538 , \22539 , \22540 ,
         \22541 , \22542 , \22543 , \22544 , \22545 , \22546 , \22547 , \22548 , \22549 , \22550 ,
         \22551 , \22552 , \22553 , \22554 , \22555 , \22556 , \22557 , \22558 , \22559 , \22560 ,
         \22561 , \22562 , \22563 , \22564 , \22565 , \22566 , \22567 , \22568 , \22569 , \22570 ,
         \22571 , \22572 , \22573 , \22574 , \22575 , \22576 , \22577 , \22578 , \22579 , \22580 ,
         \22581 , \22582 , \22583 , \22584 , \22585 , \22586 , \22587 , \22588 , \22589 , \22590 ,
         \22591 , \22592 , \22593 , \22594 , \22595 , \22596 , \22597 , \22598 , \22599 , \22600 ,
         \22601 , \22602 , \22603 , \22604 , \22605 , \22606 , \22607 , \22608 , \22609 , \22610 ,
         \22611 , \22612 , \22613 , \22614 , \22615 , \22616 , \22617 , \22618 , \22619 , \22620 ,
         \22621 , \22622 , \22623 , \22624 , \22625 , \22626 , \22627 , \22628 , \22629 , \22630 ,
         \22631 , \22632 , \22633 , \22634 , \22635 , \22636 , \22637 , \22638 , \22639 , \22640 ,
         \22641 , \22642 , \22643 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 ,
         \22651 , \22652 , \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 ,
         \22661 , \22662 , \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 ,
         \22671 , \22672 , \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 ,
         \22681 , \22682 , \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 ,
         \22691 , \22692 , \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 ,
         \22701 , \22702 , \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 ,
         \22711 , \22712 , \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 ,
         \22721 , \22722 , \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 ,
         \22731 , \22732 , \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 ,
         \22741 , \22742 , \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 ,
         \22751 , \22752 , \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 ,
         \22761 , \22762 , \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 ,
         \22771 , \22772 , \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 ,
         \22781 , \22782 , \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 ,
         \22791 , \22792 , \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 ,
         \22801 , \22802 , \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 ,
         \22811 , \22812 , \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 ,
         \22821 , \22822 , \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 ,
         \22831 , \22832 , \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 ,
         \22841 , \22842 , \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 ,
         \22851 , \22852 , \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 ,
         \22861 , \22862 , \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 ,
         \22871 , \22872 , \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 ,
         \22881 , \22882 , \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 ,
         \22891 , \22892 , \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899 , \22900 ,
         \22901 , \22902 , \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 ,
         \22911 , \22912 , \22913 , \22914 , \22915 , \22916 , \22917 , \22918 , \22919 , \22920 ,
         \22921 , \22922 , \22923 , \22924 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 ,
         \22931 , \22932 , \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 ,
         \22941 , \22942 , \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 , \22950 ,
         \22951 , \22952 , \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 ,
         \22961 , \22962 , \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 ,
         \22971 , \22972 , \22973 , \22974 , \22975 , \22976 , \22977 , \22978 , \22979 , \22980 ,
         \22981 , \22982 , \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 ,
         \22991 , \22992 , \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 ,
         \23001 , \23002 , \23003 , \23004 , \23005 , \23006 , \23007 , \23008 , \23009 , \23010 ,
         \23011 , \23012 , \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 ,
         \23021 , \23022 , \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 ,
         \23031 , \23032 , \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 ,
         \23041 , \23042 , \23043 , \23044 , \23045 , \23046 , \23047 , \23048 , \23049 , \23050 ,
         \23051 , \23052 , \23053 , \23054 , \23055 , \23056 , \23057 , \23058 , \23059 , \23060 ,
         \23061 , \23062 , \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 ,
         \23071 , \23072 , \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 ,
         \23081 , \23082 , \23083 , \23084 , \23085 , \23086 , \23087 , \23088 , \23089 , \23090 ,
         \23091 , \23092 , \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 ,
         \23101 , \23102 , \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 ,
         \23111 , \23112 , \23113 , \23114 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 ,
         \23121 , \23122 , \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 ,
         \23131 , \23132 , \23133 , \23134 , \23135 , \23136 , \23137 , \23138 , \23139 , \23140 ,
         \23141 , \23142 , \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 ,
         \23151 , \23152 , \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 ,
         \23161 , \23162 , \23163 , \23164 , \23165 , \23166 , \23167 , \23168 , \23169 , \23170 ,
         \23171 , \23172 , \23173 , \23174 , \23175 , \23176 , \23177 , \23178 , \23179 , \23180 ,
         \23181 , \23182 , \23183 , \23184 , \23185 , \23186 , \23187 , \23188 , \23189 , \23190 ,
         \23191 , \23192 , \23193 , \23194 , \23195 , \23196 , \23197 , \23198 , \23199 , \23200 ,
         \23201 , \23202 , \23203 , \23204 , \23205 , \23206 , \23207 , \23208 , \23209 , \23210 ,
         \23211 , \23212 , \23213 , \23214 , \23215 , \23216 , \23217 , \23218 , \23219 , \23220 ,
         \23221 , \23222 , \23223 , \23224 , \23225 , \23226 , \23227 , \23228 , \23229 , \23230 ,
         \23231 , \23232 , \23233 , \23234 , \23235 , \23236 , \23237 , \23238 , \23239 , \23240 ,
         \23241 , \23242 , \23243 , \23244 , \23245 , \23246 , \23247 , \23248 , \23249 , \23250 ,
         \23251 , \23252 , \23253 , \23254 , \23255 , \23256 , \23257 , \23258 , \23259 , \23260 ,
         \23261 , \23262 , \23263 , \23264 , \23265 , \23266 , \23267 , \23268 , \23269 , \23270 ,
         \23271 , \23272 , \23273 , \23274 , \23275 , \23276 , \23277 , \23278 , \23279 , \23280 ,
         \23281 , \23282 , \23283 , \23284 , \23285 , \23286 , \23287 , \23288 , \23289 , \23290 ,
         \23291 , \23292 , \23293 , \23294 , \23295 , \23296 , \23297 , \23298 , \23299 , \23300 ,
         \23301 , \23302 , \23303 , \23304 , \23305 , \23306 , \23307 , \23308 , \23309 , \23310 ,
         \23311 , \23312 , \23313 , \23314 , \23315 , \23316 , \23317 , \23318 , \23319 , \23320 ,
         \23321 , \23322 , \23323 , \23324 , \23325 , \23326 , \23327 , \23328 , \23329 , \23330 ,
         \23331 , \23332 , \23333 , \23334 , \23335 , \23336 , \23337 , \23338 , \23339 , \23340 ,
         \23341 , \23342 , \23343 , \23344 , \23345 , \23346 , \23347 , \23348 , \23349 , \23350 ,
         \23351 , \23352 , \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 ,
         \23361 , \23362 , \23363 , \23364 , \23365 , \23366 , \23367 , \23368 , \23369 , \23370 ,
         \23371 , \23372 , \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 ,
         \23381 , \23382 , \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 ,
         \23391 , \23392 , \23393 , \23394 , \23395 , \23396 , \23397 , \23398 , \23399 , \23400 ,
         \23401 , \23402 , \23403 , \23404 , \23405 , \23406 , \23407 , \23408 , \23409 , \23410 ,
         \23411 , \23412 , \23413 , \23414 , \23415 , \23416 , \23417 , \23418 , \23419 , \23420 ,
         \23421 , \23422 , \23423 , \23424 , \23425 , \23426 , \23427 , \23428 , \23429 , \23430 ,
         \23431 , \23432 , \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 ,
         \23441 , \23442 , \23443 , \23444 , \23445 , \23446 , \23447 , \23448 , \23449 , \23450 ,
         \23451 , \23452 , \23453 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 ,
         \23461 , \23462 , \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 , \23470 ,
         \23471 , \23472 , \23473 , \23474 , \23475 , \23476 , \23477 , \23478 , \23479 , \23480 ,
         \23481 , \23482 , \23483 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 ,
         \23491 , \23492 , \23493 , \23494 , \23495 , \23496 , \23497 , \23498 , \23499 , \23500 ,
         \23501 , \23502 , \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 ,
         \23511 , \23512 , \23513 , \23514 , \23515 , \23516 , \23517 , \23518 , \23519 , \23520 ,
         \23521 , \23522 , \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 ,
         \23531 , \23532 , \23533 , \23534 , \23535 , \23536 , \23537 , \23538 , \23539 , \23540 ,
         \23541 , \23542 , \23543 , \23544 , \23545 , \23546 , \23547 , \23548 , \23549 , \23550 ,
         \23551 , \23552 , \23553 , \23554 , \23555 , \23556 , \23557 , \23558 , \23559 , \23560 ,
         \23561 , \23562 , \23563 , \23564 , \23565 , \23566 , \23567 , \23568 , \23569 , \23570 ,
         \23571 , \23572 , \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 ,
         \23581 , \23582 , \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 ,
         \23591 , \23592 , \23593 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 ,
         \23601 , \23602 , \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 ,
         \23611 , \23612 , \23613 , \23614 , \23615 , \23616 , \23617 , \23618 , \23619 , \23620 ,
         \23621 , \23622 , \23623 , \23624 , \23625 , \23626 , \23627 , \23628 , \23629 , \23630 ,
         \23631 , \23632 , \23633 , \23634 , \23635 , \23636 , \23637 , \23638 , \23639 , \23640 ,
         \23641 , \23642 , \23643 , \23644 , \23645 , \23646 , \23647 , \23648 , \23649 , \23650 ,
         \23651 , \23652 , \23653 , \23654 , \23655 , \23656 , \23657 , \23658 , \23659 , \23660 ,
         \23661 , \23662 , \23663 , \23664 , \23665 , \23666 , \23667 , \23668 , \23669 , \23670 ,
         \23671 , \23672 , \23673 , \23674 , \23675 , \23676 , \23677 , \23678 , \23679 , \23680 ,
         \23681 , \23682 , \23683 , \23684 , \23685 , \23686 , \23687 , \23688 , \23689 , \23690 ,
         \23691 , \23692 , \23693 , \23694 , \23695 , \23696 , \23697 , \23698 , \23699 , \23700 ,
         \23701 , \23702 , \23703 , \23704 , \23705 , \23706 , \23707 , \23708 , \23709 , \23710 ,
         \23711 , \23712 , \23713 , \23714 , \23715 , \23716 , \23717 , \23718 , \23719 , \23720 ,
         \23721 , \23722 , \23723 , \23724 , \23725 , \23726 , \23727 , \23728 , \23729 , \23730 ,
         \23731 , \23732 , \23733 , \23734 , \23735 , \23736 , \23737 , \23738 , \23739 , \23740 ,
         \23741 , \23742 , \23743 , \23744 , \23745 , \23746 , \23747 , \23748 , \23749 , \23750 ,
         \23751 , \23752 , \23753 , \23754 , \23755 , \23756 , \23757 , \23758 , \23759 , \23760 ,
         \23761 , \23762 , \23763 , \23764 , \23765 , \23766 , \23767 , \23768 , \23769 , \23770 ,
         \23771 , \23772 , \23773 , \23774 , \23775 , \23776 , \23777 , \23778 , \23779 , \23780 ,
         \23781 , \23782 , \23783 , \23784 , \23785 , \23786 , \23787 , \23788 , \23789 , \23790 ,
         \23791 , \23792 , \23793 , \23794 , \23795 , \23796 , \23797 , \23798 , \23799 , \23800 ,
         \23801 , \23802 , \23803 , \23804 , \23805 , \23806 , \23807 , \23808 , \23809 , \23810 ,
         \23811 , \23812 , \23813 , \23814 , \23815 , \23816 , \23817 , \23818 , \23819 , \23820 ,
         \23821 , \23822 , \23823 , \23824 , \23825 , \23826 , \23827 , \23828 , \23829 , \23830 ,
         \23831 , \23832 , \23833 , \23834 , \23835 , \23836 , \23837 , \23838 , \23839 , \23840 ,
         \23841 , \23842 , \23843 , \23844 , \23845 , \23846 , \23847 , \23848 , \23849 , \23850 ,
         \23851 , \23852 , \23853 , \23854 , \23855 , \23856 , \23857 , \23858 , \23859 , \23860 ,
         \23861 , \23862 , \23863 , \23864 , \23865 , \23866 , \23867 , \23868 , \23869 , \23870 ,
         \23871 , \23872 , \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 ,
         \23881 , \23882 , \23883 , \23884 , \23885 , \23886 , \23887 , \23888 , \23889 , \23890 ,
         \23891 , \23892 , \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 ,
         \23901 , \23902 , \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 ,
         \23911 , \23912 , \23913 , \23914 , \23915 , \23916 , \23917 , \23918 , \23919 , \23920 ,
         \23921 , \23922 , \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 ,
         \23931 , \23932 , \23933 , \23934 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 ,
         \23941 , \23942 , \23943 , \23944 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 ,
         \23951 , \23952 , \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 ,
         \23961 , \23962 , \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 , \23970 ,
         \23971 , \23972 , \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 ,
         \23981 , \23982 , \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 ,
         \23991 , \23992 , \23993 , \23994 , \23995 , \23996 , \23997 , \23998 , \23999 , \24000 ,
         \24001 , \24002 , \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 ,
         \24011 , \24012 , \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 ,
         \24021 , \24022 , \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 ,
         \24031 , \24032 , \24033 , \24034 , \24035 , \24036 , \24037 , \24038 , \24039 , \24040 ,
         \24041 , \24042 , \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 ,
         \24051 , \24052 , \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 ,
         \24061 , \24062 , \24063 , \24064 , \24065 , \24066 , \24067 , \24068 , \24069 , \24070 ,
         \24071 , \24072 , \24073 , \24074 , \24075 , \24076 , \24077 , \24078 , \24079 , \24080 ,
         \24081 , \24082 , \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 ,
         \24091 , \24092 , \24093 , \24094 , \24095 , \24096 , \24097 , \24098 , \24099 , \24100 ,
         \24101 , \24102 , \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 ,
         \24111 , \24112 , \24113 , \24114 , \24115 , \24116 , \24117 , \24118 , \24119 , \24120 ,
         \24121 , \24122 , \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 ,
         \24131 , \24132 , \24133 , \24134 , \24135 , \24136 , \24137 , \24138 , \24139 , \24140 ,
         \24141 , \24142 , \24143 , \24144 , \24145 , \24146 , \24147 , \24148 , \24149 , \24150 ,
         \24151 , \24152 , \24153 , \24154 , \24155 , \24156 , \24157 , \24158 , \24159 , \24160 ,
         \24161 , \24162 , \24163 , \24164 , \24165 , \24166 , \24167 , \24168 , \24169 , \24170 ,
         \24171 , \24172 , \24173 , \24174 , \24175 , \24176 , \24177 , \24178 , \24179 , \24180 ,
         \24181 , \24182 , \24183 , \24184 , \24185 , \24186 , \24187 , \24188 , \24189 , \24190 ,
         \24191 , \24192 , \24193 , \24194 , \24195 , \24196 , \24197 , \24198 , \24199 , \24200 ,
         \24201 , \24202 , \24203 , \24204 , \24205 , \24206 , \24207 , \24208 , \24209 , \24210 ,
         \24211 , \24212 , \24213 , \24214 , \24215 , \24216 , \24217 , \24218 , \24219 , \24220 ,
         \24221 , \24222 , \24223 , \24224 , \24225 , \24226 , \24227 , \24228 , \24229 , \24230 ,
         \24231 , \24232 , \24233 , \24234 , \24235 , \24236 , \24237 , \24238 , \24239 , \24240 ,
         \24241 , \24242 , \24243 , \24244 , \24245 , \24246 , \24247 , \24248 , \24249 , \24250 ,
         \24251 , \24252 , \24253 , \24254 , \24255 , \24256 , \24257 , \24258 , \24259 , \24260 ,
         \24261 , \24262 , \24263 , \24264 , \24265 , \24266 , \24267 , \24268 , \24269 , \24270 ,
         \24271 , \24272 , \24273 , \24274 , \24275 , \24276 , \24277 , \24278 , \24279 , \24280 ,
         \24281 , \24282 , \24283 , \24284 , \24285 , \24286 , \24287 , \24288 , \24289 , \24290 ,
         \24291 , \24292 , \24293 , \24294 , \24295 , \24296 , \24297 , \24298 , \24299 , \24300 ,
         \24301 , \24302 , \24303 , \24304 , \24305 , \24306 , \24307 , \24308 , \24309 , \24310 ,
         \24311 , \24312 , \24313 , \24314 , \24315 , \24316 , \24317 , \24318 , \24319 , \24320 ,
         \24321 , \24322 , \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 ,
         \24331 , \24332 , \24333 , \24334 , \24335 , \24336 , \24337 , \24338 , \24339 , \24340 ,
         \24341 , \24342 , \24343 , \24344 , \24345 , \24346 , \24347 , \24348 , \24349 , \24350 ,
         \24351 , \24352 , \24353 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 ,
         \24361 , \24362 , \24363 , \24364 , \24365 , \24366 , \24367 , \24368 , \24369 , \24370 ,
         \24371 , \24372 , \24373 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , \24380 ,
         \24381 , \24382 , \24383 , \24384 , \24385 , \24386 , \24387 , \24388 , \24389 , \24390 ,
         \24391 , \24392 , \24393 , \24394 , \24395 , \24396 , \24397 , \24398 , \24399 , \24400 ,
         \24401 , \24402 , \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 ,
         \24411 , \24412 , \24413 , \24414 , \24415 , \24416 , \24417 , \24418 , \24419 , \24420 ,
         \24421 , \24422 , \24423 , \24424 , \24425 , \24426 , \24427 , \24428 , \24429 , \24430 ,
         \24431 , \24432 , \24433 , \24434 , \24435 , \24436 , \24437 , \24438 , \24439 , \24440 ,
         \24441 , \24442 , \24443 , \24444 , \24445 , \24446 , \24447 , \24448 , \24449 , \24450 ,
         \24451 , \24452 , \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 ,
         \24461 , \24462 , \24463 , \24464 , \24465 , \24466 , \24467 , \24468 , \24469 , \24470 ,
         \24471 , \24472 , \24473 , \24474 , \24475 , \24476 , \24477 , \24478 , \24479 , \24480 ,
         \24481 , \24482 , \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 ,
         \24491 , \24492 , \24493 , \24494 , \24495 , \24496 , \24497 , \24498 , \24499 , \24500 ,
         \24501 , \24502 , \24503 , \24504 , \24505 , \24506 , \24507 , \24508 , \24509 , \24510 ,
         \24511 , \24512 , \24513 , \24514 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 ,
         \24521 , \24522 , \24523 , \24524 , \24525 , \24526 , \24527 , \24528 , \24529 , \24530 ,
         \24531 , \24532 , \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 ,
         \24541 , \24542 , \24543 , \24544 , \24545 , \24546 , \24547 , \24548 , \24549 , \24550 ,
         \24551 , \24552 , \24553 , \24554 , \24555 , \24556 , \24557 , \24558 , \24559 , \24560 ,
         \24561 , \24562 , \24563 , \24564 , \24565 , \24566 , \24567 , \24568 , \24569 , \24570 ,
         \24571 , \24572 , \24573 , \24574 , \24575 , \24576 , \24577 , \24578 , \24579 , \24580 ,
         \24581 , \24582 , \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 ,
         \24591 , \24592 , \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 ,
         \24601 , \24602 , \24603 , \24604 , \24605 , \24606 , \24607 , \24608 , \24609 , \24610 ,
         \24611 , \24612 , \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 ,
         \24621 , \24622 , \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 ,
         \24631 , \24632 , \24633 , \24634 , \24635 , \24636 , \24637 , \24638 , \24639 , \24640 ,
         \24641 , \24642 , \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 ,
         \24651 , \24652 , \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 ,
         \24661 , \24662 , \24663 , \24664 , \24665 , \24666 , \24667 , \24668 , \24669 , \24670 ,
         \24671 , \24672 , \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 ,
         \24681 , \24682 , \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 ,
         \24691 , \24692 , \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 ,
         \24701 , \24702 , \24703 , \24704 , \24705 , \24706 , \24707 , \24708 , \24709 , \24710 ,
         \24711 , \24712 , \24713 , \24714 , \24715 , \24716 , \24717 , \24718 , \24719 , \24720 ,
         \24721 , \24722 , \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 ,
         \24731 , \24732 , \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 ,
         \24741 , \24742 , \24743 , \24744 , \24745 , \24746 , \24747 , \24748 , \24749 , \24750 ,
         \24751 , \24752 , \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 ,
         \24761 , \24762 , \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 , \24770 ,
         \24771 , \24772 , \24773 , \24774 , \24775 , \24776 , \24777 , \24778 , \24779 , \24780 ,
         \24781 , \24782 , \24783 , \24784 , \24785 , \24786 , \24787 , \24788 , \24789 , \24790 ,
         \24791 , \24792 , \24793 , \24794 , \24795 , \24796 , \24797 , \24798 , \24799 , \24800 ,
         \24801 , \24802 , \24803 , \24804 , \24805 , \24806 , \24807 , \24808 , \24809 , \24810 ,
         \24811 , \24812 , \24813 , \24814 , \24815 , \24816 , \24817 , \24818 , \24819 , \24820 ,
         \24821 , \24822 , \24823 , \24824 , \24825 , \24826 , \24827 , \24828 , \24829 , \24830 ,
         \24831 , \24832 , \24833 , \24834 , \24835 , \24836 , \24837 , \24838 , \24839 , \24840 ,
         \24841 , \24842 , \24843 , \24844 , \24845 , \24846 , \24847 , \24848 , \24849 , \24850 ,
         \24851 , \24852 , \24853 , \24854 , \24855 , \24856 , \24857 , \24858 , \24859 , \24860 ,
         \24861 , \24862 , \24863 , \24864 , \24865 , \24866 , \24867 , \24868 , \24869 , \24870 ,
         \24871 , \24872 , \24873 , \24874 , \24875 , \24876 , \24877 , \24878 , \24879 , \24880 ,
         \24881 , \24882 , \24883 , \24884 , \24885 , \24886 , \24887 , \24888 , \24889 , \24890 ,
         \24891 , \24892 , \24893 , \24894 , \24895 , \24896 , \24897 , \24898 , \24899 , \24900 ,
         \24901 , \24902 , \24903 , \24904 , \24905 , \24906 , \24907 , \24908 , \24909 , \24910 ,
         \24911 , \24912 , \24913 , \24914 , \24915 , \24916 , \24917 , \24918 , \24919 , \24920 ,
         \24921 , \24922 , \24923 , \24924 , \24925 , \24926 , \24927 , \24928 , \24929 , \24930 ,
         \24931 , \24932 , \24933 , \24934 , \24935 , \24936 , \24937 , \24938 , \24939 , \24940 ,
         \24941 , \24942 , \24943 , \24944 , \24945 , \24946 , \24947 , \24948 , \24949 , \24950 ,
         \24951 , \24952 , \24953 , \24954 , \24955 , \24956 , \24957 , \24958 , \24959 , \24960 ,
         \24961 , \24962 , \24963 , \24964 , \24965 , \24966 , \24967 , \24968 , \24969 , \24970 ,
         \24971 , \24972 , \24973 , \24974 , \24975 , \24976 , \24977 , \24978 , \24979 , \24980 ,
         \24981 , \24982 , \24983 , \24984 , \24985 , \24986 , \24987 , \24988 , \24989 , \24990 ,
         \24991 , \24992 , \24993 , \24994 , \24995 , \24996 , \24997 , \24998 , \24999 , \25000 ,
         \25001 , \25002 , \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 ,
         \25011 , \25012 , \25013 , \25014 , \25015 , \25016 , \25017 , \25018 , \25019 , \25020 ,
         \25021 , \25022 , \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 ,
         \25031 , \25032 , \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 ,
         \25041 , \25042 , \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 ,
         \25051 , \25052 , \25053 , \25054 , \25055 , \25056 , \25057 , \25058 , \25059 , \25060 ,
         \25061 , \25062 , \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 ,
         \25071 , \25072 , \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 ,
         \25081 , \25082 , \25083 , \25084 , \25085 , \25086 , \25087 , \25088 , \25089 , \25090 ,
         \25091 , \25092 , \25093 , \25094 , \25095 , \25096 , \25097 , \25098 , \25099 , \25100 ,
         \25101 , \25102 , \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 ,
         \25111 , \25112 , \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 ,
         \25121 , \25122 , \25123 , \25124 , \25125 , \25126 , \25127 , \25128 , \25129 , \25130 ,
         \25131 , \25132 , \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 ,
         \25141 , \25142 , \25143 , \25144 , \25145 , \25146 , \25147 , \25148 , \25149 , \25150 ,
         \25151 , \25152 , \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 ,
         \25161 , \25162 , \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 ,
         \25171 , \25172 , \25173 , \25174 , \25175 , \25176 , \25177 , \25178 , \25179 , \25180 ,
         \25181 , \25182 , \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 ,
         \25191 , \25192 , \25193 , \25194 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 ,
         \25201 , \25202 , \25203 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 ,
         \25211 , \25212 , \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 ,
         \25221 , \25222 , \25223 , \25224 , \25225 , \25226 , \25227 , \25228 , \25229 , \25230 ,
         \25231 , \25232 , \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 ,
         \25241 , \25242 , \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 ,
         \25251 , \25252 , \25253 , \25254 , \25255 , \25256 , \25257 , \25258 , \25259 , \25260 ,
         \25261 , \25262 , \25263 , \25264 , \25265 , \25266 , \25267 , \25268 , \25269 , \25270 ,
         \25271 , \25272 , \25273 , \25274 , \25275 , \25276 , \25277 , \25278 , \25279 , \25280 ,
         \25281 , \25282 , \25283 , \25284 , \25285 , \25286 , \25287 , \25288 , \25289 , \25290 ,
         \25291 , \25292 , \25293 , \25294 , \25295 , \25296 , \25297 , \25298 , \25299 , \25300 ,
         \25301 , \25302 , \25303 , \25304 , \25305 , \25306 , \25307 , \25308 , \25309 , \25310 ,
         \25311 , \25312 , \25313 , \25314 , \25315 , \25316 , \25317 , \25318 , \25319 , \25320 ,
         \25321 , \25322 , \25323 , \25324 , \25325 , \25326 , \25327 , \25328 , \25329 , \25330 ,
         \25331 , \25332 , \25333 , \25334 , \25335 , \25336 , \25337 , \25338 , \25339 , \25340 ,
         \25341 , \25342 , \25343 , \25344 , \25345 , \25346 , \25347 , \25348 , \25349 , \25350 ,
         \25351 , \25352 , \25353 , \25354 , \25355 , \25356 , \25357 , \25358 , \25359 , \25360 ,
         \25361 , \25362 , \25363 , \25364 , \25365 , \25366 , \25367 , \25368 , \25369 , \25370 ,
         \25371 , \25372 , \25373 , \25374 , \25375 , \25376 , \25377 , \25378 , \25379 , \25380 ,
         \25381 , \25382 , \25383 , \25384 , \25385 , \25386 , \25387 , \25388 , \25389 , \25390 ,
         \25391 , \25392 , \25393 , \25394 , \25395 , \25396 , \25397 , \25398 , \25399 , \25400 ,
         \25401 , \25402 , \25403 , \25404 , \25405 , \25406 , \25407 , \25408 , \25409 , \25410 ,
         \25411 , \25412 , \25413 , \25414 , \25415 , \25416 , \25417 , \25418 , \25419 , \25420 ,
         \25421 , \25422 , \25423 , \25424 , \25425 , \25426 , \25427 , \25428 , \25429 , \25430 ,
         \25431 , \25432 , \25433 , \25434 , \25435 , \25436 , \25437 , \25438 , \25439 , \25440 ,
         \25441 , \25442 , \25443 , \25444 , \25445 , \25446 , \25447 , \25448 , \25449 , \25450 ,
         \25451 , \25452 , \25453 , \25454 , \25455 , \25456 , \25457 , \25458 , \25459 , \25460 ,
         \25461 , \25462 , \25463 , \25464 , \25465 , \25466 , \25467 , \25468 , \25469 , \25470 ,
         \25471 , \25472 , \25473 , \25474 , \25475 , \25476 , \25477 , \25478 , \25479 , \25480 ,
         \25481 , \25482 , \25483 , \25484 , \25485 , \25486 , \25487 , \25488 , \25489 , \25490 ,
         \25491 , \25492 , \25493 , \25494 , \25495 , \25496 , \25497 , \25498 , \25499 , \25500 ,
         \25501 , \25502 , \25503 , \25504 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 ,
         \25511 , \25512 , \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 ,
         \25521 , \25522 , \25523 , \25524 , \25525 , \25526 , \25527 , \25528 , \25529 , \25530 ,
         \25531 , \25532 , \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 ,
         \25541 , \25542 , \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 ,
         \25551 , \25552 , \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 ,
         \25561 , \25562 , \25563 , \25564 , \25565 , \25566 , \25567 , \25568 , \25569 , \25570 ,
         \25571 , \25572 , \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 ,
         \25581 , \25582 , \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 ,
         \25591 , \25592 , \25593 , \25594 , \25595 , \25596 , \25597 , \25598 , \25599 , \25600 ,
         \25601 , \25602 , \25603 , \25604 , \25605 , \25606 , \25607 , \25608 , \25609 , \25610 ,
         \25611 , \25612 , \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 ,
         \25621 , \25622 , \25623 , \25624 , \25625 , \25626 , \25627 , \25628 , \25629 , \25630 ,
         \25631 , \25632 , \25633 , \25634 , \25635 , \25636 , \25637 , \25638 , \25639 , \25640 ,
         \25641 , \25642 , \25643 , \25644 , \25645 , \25646 , \25647 , \25648 , \25649 , \25650 ,
         \25651 , \25652 , \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 ,
         \25661 , \25662 , \25663 , \25664 , \25665 , \25666 , \25667 , \25668 , \25669 , \25670 ,
         \25671 , \25672 , \25673 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 ,
         \25681 , \25682 , \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 , \25690 ,
         \25691 , \25692 , \25693 , \25694 , \25695 , \25696 , \25697 , \25698 , \25699 , \25700 ,
         \25701 , \25702 , \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 ,
         \25711 , \25712 , \25713 , \25714 , \25715 , \25716 , \25717 , \25718 , \25719 , \25720 ,
         \25721 , \25722 , \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 ,
         \25731 , \25732 , \25733 , \25734 , \25735 , \25736 , \25737 , \25738 , \25739 , \25740 ,
         \25741 , \25742 , \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 ,
         \25751 , \25752 , \25753 , \25754 , \25755 , \25756 , \25757 , \25758 , \25759 , \25760 ,
         \25761 , \25762 , \25763 , \25764 , \25765 , \25766 , \25767 , \25768 , \25769 , \25770 ,
         \25771 , \25772 , \25773 , \25774 , \25775 , \25776 , \25777 , \25778 , \25779 , \25780 ,
         \25781 , \25782 , \25783 , \25784 , \25785 , \25786 , \25787 , \25788 , \25789 , \25790 ,
         \25791 , \25792 , \25793 , \25794 , \25795 , \25796 , \25797 , \25798 , \25799 , \25800 ,
         \25801 , \25802 , \25803 , \25804 , \25805 , \25806 , \25807 , \25808 , \25809 , \25810 ,
         \25811 , \25812 , \25813 , \25814 , \25815 , \25816 , \25817 , \25818 , \25819 , \25820 ,
         \25821 , \25822 , \25823 , \25824 , \25825 , \25826 , \25827 , \25828 , \25829 , \25830 ,
         \25831 , \25832 , \25833 , \25834 , \25835 , \25836 , \25837 , \25838 , \25839 , \25840 ,
         \25841 , \25842 , \25843 , \25844 , \25845 , \25846 , \25847 , \25848 , \25849 , \25850 ,
         \25851 , \25852 , \25853 , \25854 , \25855 , \25856 , \25857 , \25858 , \25859 , \25860 ,
         \25861 , \25862 , \25863 , \25864 , \25865 , \25866 , \25867 , \25868 , \25869 , \25870 ,
         \25871 , \25872 , \25873 , \25874 , \25875 , \25876 , \25877 , \25878 , \25879 , \25880 ,
         \25881 , \25882 , \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 ,
         \25891 , \25892 , \25893 , \25894 , \25895 , \25896 , \25897 , \25898 , \25899 , \25900 ,
         \25901 , \25902 , \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 ,
         \25911 , \25912 , \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 ,
         \25921 , \25922 , \25923 , \25924 , \25925 , \25926 , \25927 , \25928 , \25929 , \25930 ,
         \25931 , \25932 , \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 ,
         \25941 , \25942 , \25943 , \25944 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 ,
         \25951 , \25952 , \25953 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 ,
         \25961 , \25962 , \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 ,
         \25971 , \25972 , \25973 , \25974 , \25975 , \25976 , \25977 , \25978 , \25979 , \25980 ,
         \25981 , \25982 , \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 ,
         \25991 , \25992 , \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 ,
         \26001 , \26002 , \26003 , \26004 , \26005 , \26006 , \26007 , \26008 , \26009 , \26010 ,
         \26011 , \26012 , \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 ,
         \26021 , \26022 , \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 ,
         \26031 , \26032 , \26033 , \26034 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 ,
         \26041 , \26042 , \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 ,
         \26051 , \26052 , \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 , \26060 ,
         \26061 , \26062 , \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 ,
         \26071 , \26072 , \26073 , \26074 , \26075 , \26076 , \26077 , \26078 , \26079 , \26080 ,
         \26081 , \26082 , \26083 , \26084 , \26085 , \26086 , \26087 , \26088 , \26089 , \26090 ,
         \26091 , \26092 , \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 ,
         \26101 , \26102 , \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 ,
         \26111 , \26112 , \26113 , \26114 , \26115 , \26116 , \26117 , \26118 , \26119 , \26120 ,
         \26121 , \26122 , \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 ,
         \26131 , \26132 , \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 ,
         \26141 , \26142 , \26143 , \26144 , \26145 , \26146 , \26147 , \26148 , \26149 , \26150 ,
         \26151 , \26152 , \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 ,
         \26161 , \26162 , \26163 , \26164 , \26165 , \26166 , \26167 , \26168 , \26169 , \26170 ,
         \26171 , \26172 , \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 ,
         \26181 , \26182 , \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 ,
         \26191 , \26192 , \26193 , \26194 , \26195 , \26196 , \26197 , \26198 , \26199 , \26200 ,
         \26201 , \26202 , \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 ,
         \26211 , \26212 , \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 ,
         \26221 , \26222 , \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 ,
         \26231 , \26232 , \26233 , \26234 , \26235 , \26236 , \26237 , \26238 , \26239 , \26240 ,
         \26241 , \26242 , \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 ,
         \26251 , \26252 , \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 ,
         \26261 , \26262 , \26263 , \26264 , \26265 , \26266 , \26267 , \26268 , \26269 , \26270 ,
         \26271 , \26272 , \26273 , \26274 , \26275 , \26276 , \26277 , \26278 , \26279 , \26280 ,
         \26281 , \26282 , \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 ,
         \26291 , \26292 , \26293 , \26294 , \26295 , \26296 , \26297 , \26298 , \26299 , \26300 ,
         \26301 , \26302 , \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 ,
         \26311 , \26312 , \26313 , \26314 , \26315 , \26316 , \26317 , \26318 , \26319 , \26320 ,
         \26321 , \26322 , \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 ,
         \26331 , \26332 , \26333 , \26334 , \26335 , \26336 , \26337 , \26338 , \26339 , \26340 ,
         \26341 , \26342 , \26343 , \26344 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 ,
         \26351 , \26352 , \26353 , \26354 , \26355 , \26356 , \26357 , \26358 , \26359 , \26360 ,
         \26361 , \26362 , \26363 , \26364 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 ,
         \26371 , \26372 , \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 ,
         \26381 , \26382 , \26383 , \26384 , \26385 , \26386 , \26387 , \26388 , \26389 , \26390 ,
         \26391 , \26392 , \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 ,
         \26401 , \26402 , \26403 , \26404 , \26405 , \26406 , \26407 , \26408 , \26409 , \26410 ,
         \26411 , \26412 , \26413 , \26414 , \26415 , \26416 , \26417 , \26418 , \26419 , \26420 ,
         \26421 , \26422 , \26423 , \26424 , \26425 , \26426 , \26427 , \26428 , \26429 , \26430 ,
         \26431 , \26432 , \26433 , \26434 , \26435 , \26436 , \26437 , \26438 , \26439 , \26440 ,
         \26441 , \26442 , \26443 , \26444 , \26445 , \26446 , \26447 , \26448 , \26449 , \26450 ,
         \26451 , \26452 , \26453 , \26454 , \26455 , \26456 , \26457 , \26458 , \26459 , \26460 ,
         \26461 , \26462 , \26463 , \26464 , \26465 , \26466 , \26467 , \26468 , \26469 , \26470 ,
         \26471 , \26472 , \26473 , \26474 , \26475 , \26476 , \26477 , \26478 , \26479 , \26480 ,
         \26481 , \26482 , \26483 , \26484 , \26485 , \26486 , \26487 , \26488 , \26489 , \26490 ,
         \26491 , \26492 , \26493 , \26494 , \26495 , \26496 , \26497 , \26498 , \26499 , \26500 ,
         \26501 , \26502 , \26503 , \26504 , \26505 , \26506 , \26507 , \26508 , \26509 , \26510 ,
         \26511 , \26512 , \26513 , \26514 , \26515 , \26516 , \26517 , \26518 , \26519 , \26520 ,
         \26521 , \26522 , \26523 , \26524 , \26525 , \26526 , \26527 , \26528 , \26529 , \26530 ,
         \26531 , \26532 , \26533 , \26534 , \26535 , \26536 , \26537 , \26538 , \26539 , \26540 ,
         \26541 , \26542 , \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , \26549 , \26550 ,
         \26551 , \26552 , \26553 , \26554 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 ,
         \26561 , \26562 , \26563 , \26564 , \26565 , \26566 , \26567 , \26568 , \26569 , \26570 ,
         \26571 , \26572 , \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 ,
         \26581 , \26582 , \26583 , \26584 , \26585 , \26586 , \26587 , \26588 , \26589 , \26590 ,
         \26591 , \26592 , \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , \26600 ,
         \26601 , \26602 , \26603 , \26604 , \26605 , \26606 , \26607 , \26608 , \26609 , \26610 ,
         \26611 , \26612 , \26613 , \26614 , \26615 , \26616 , \26617 , \26618 , \26619 , \26620 ,
         \26621 , \26622 , \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 ,
         \26631 , \26632 , \26633 , \26634 , \26635 , \26636 , \26637 , \26638 , \26639 , \26640 ,
         \26641 , \26642 , \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 ,
         \26651 , \26652 , \26653 , \26654 , \26655 , \26656 , \26657 , \26658 , \26659 , \26660 ,
         \26661 , \26662 , \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , \26669 , \26670 ,
         \26671 , \26672 , \26673 , \26674 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 ,
         \26681 , \26682 , \26683 , \26684 , \26685 , \26686 , \26687 , \26688 , \26689 , \26690 ,
         \26691 , \26692 , \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 ,
         \26701 , \26702 , \26703 , \26704 , \26705 , \26706 , \26707 , \26708 , \26709 , \26710 ,
         \26711 , \26712 , \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , \26720 ,
         \26721 , \26722 , \26723 , \26724 , \26725 , \26726 , \26727 , \26728 , \26729 , \26730 ,
         \26731 , \26732 , \26733 , \26734 , \26735 , \26736 , \26737 , \26738 , \26739 , \26740 ,
         \26741 , \26742 , \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 ,
         \26751 , \26752 , \26753 , \26754 , \26755 , \26756 , \26757 , \26758 , \26759 , \26760 ,
         \26761 , \26762 , \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 ,
         \26771 , \26772 , \26773 , \26774 , \26775 , \26776 , \26777 , \26778 , \26779 , \26780 ,
         \26781 , \26782 , \26783 , \26784 , \26785 , \26786 , \26787 , \26788 , \26789 , \26790 ,
         \26791 , \26792 , \26793 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 ,
         \26801 , \26802 , \26803 , \26804 , \26805 , \26806 , \26807 , \26808 , \26809 , \26810 ,
         \26811 , \26812 , \26813 , \26814 , \26815 , \26816 , \26817 , \26818 , \26819 , \26820 ,
         \26821 , \26822 , \26823 , \26824 , \26825 , \26826 , \26827 , \26828 , \26829 , \26830 ,
         \26831 , \26832 , \26833 , \26834 , \26835 , \26836 , \26837 , \26838 , \26839 , \26840 ,
         \26841 , \26842 , \26843 , \26844 , \26845 , \26846 , \26847 , \26848 , \26849 , \26850 ,
         \26851 , \26852 , \26853 , \26854 , \26855 , \26856 , \26857 , \26858 , \26859 , \26860 ,
         \26861 , \26862 , \26863 , \26864 , \26865 , \26866 , \26867 , \26868 , \26869 , \26870 ,
         \26871 , \26872 , \26873 , \26874 , \26875 , \26876 , \26877 , \26878 , \26879 , \26880 ,
         \26881 , \26882 , \26883 , \26884 , \26885 , \26886 , \26887 , \26888 , \26889 , \26890 ,
         \26891 , \26892 , \26893 , \26894 , \26895 , \26896 , \26897 , \26898 , \26899 , \26900 ,
         \26901 , \26902 , \26903 , \26904 , \26905 , \26906 , \26907 , \26908 , \26909 , \26910 ,
         \26911 , \26912 , \26913 , \26914 , \26915 , \26916 , \26917 , \26918 , \26919 , \26920 ,
         \26921 , \26922 , \26923 , \26924 , \26925 , \26926 , \26927 , \26928 , \26929 , \26930 ,
         \26931 , \26932 , \26933 , \26934 , \26935 , \26936 , \26937 , \26938 , \26939 , \26940 ,
         \26941 , \26942 , \26943 , \26944 , \26945 , \26946 , \26947 , \26948 , \26949 , \26950 ,
         \26951 , \26952 , \26953 , \26954 , \26955 , \26956 , \26957 , \26958 , \26959 , \26960 ,
         \26961 , \26962 , \26963 , \26964 , \26965 , \26966 , \26967 , \26968 , \26969 , \26970 ,
         \26971 , \26972 , \26973 , \26974 , \26975 , \26976 , \26977 , \26978 , \26979 , \26980 ,
         \26981 , \26982 , \26983 , \26984 , \26985 , \26986 , \26987 , \26988 , \26989 , \26990 ,
         \26991 , \26992 , \26993 , \26994 , \26995 , \26996 , \26997 , \26998 , \26999 , \27000 ,
         \27001 , \27002 , \27003 , \27004 , \27005 , \27006 , \27007 , \27008 , \27009 , \27010 ,
         \27011 , \27012 , \27013 , \27014 , \27015 , \27016 , \27017 , \27018 , \27019 , \27020 ,
         \27021 , \27022 , \27023 , \27024 , \27025 , \27026 , \27027 , \27028 , \27029 , \27030 ,
         \27031 , \27032 , \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 , \27040 ,
         \27041 , \27042 , \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 ,
         \27051 , \27052 , \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 ,
         \27061 , \27062 , \27063 , \27064 , \27065 , \27066 , \27067 , \27068 , \27069 , \27070 ,
         \27071 , \27072 , \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 ,
         \27081 , \27082 , \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 ,
         \27091 , \27092 , \27093 , \27094 , \27095 , \27096 , \27097 , \27098 , \27099 , \27100 ,
         \27101 , \27102 , \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 ,
         \27111 , \27112 , \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 ,
         \27121 , \27122 , \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 ,
         \27131 , \27132 , \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 ,
         \27141 , \27142 , \27143 , \27144 , \27145 , \27146 , \27147 , \27148 , \27149 , \27150 ,
         \27151 , \27152 , \27153 , \27154 , \27155 , \27156 , \27157 , \27158 , \27159 , \27160 ,
         \27161 , \27162 , \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 ,
         \27171 , \27172 , \27173 , \27174 , \27175 , \27176 , \27177 , \27178 , \27179 , \27180 ,
         \27181 , \27182 , \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 ,
         \27191 , \27192 , \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 ,
         \27201 , \27202 , \27203 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 ,
         \27211 , \27212 , \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 ,
         \27221 , \27222 , \27223 , \27224 , \27225 , \27226 , \27227 , \27228 , \27229 , \27230 ,
         \27231 , \27232 , \27233 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 ,
         \27241 , \27242 , \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 ,
         \27251 , \27252 , \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 ,
         \27261 , \27262 , \27263 , \27264 , \27265 , \27266 , \27267 , \27268 , \27269 , \27270 ,
         \27271 , \27272 , \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 ,
         \27281 , \27282 , \27283 , \27284 , \27285 , \27286 , \27287 , \27288 , \27289 , \27290 ,
         \27291 , \27292 , \27293 , \27294 , \27295 , \27296 , \27297 , \27298 , \27299 , \27300 ,
         \27301 , \27302 , \27303 , \27304 , \27305 , \27306 , \27307 , \27308 , \27309 , \27310 ,
         \27311 , \27312 , \27313 , \27314 , \27315 , \27316 , \27317 , \27318 , \27319 , \27320 ,
         \27321 , \27322 , \27323 , \27324 , \27325 , \27326 , \27327 , \27328 , \27329 , \27330 ,
         \27331 , \27332 , \27333 , \27334 , \27335 , \27336 , \27337 , \27338 , \27339 , \27340 ,
         \27341 , \27342 , \27343 , \27344 , \27345 , \27346 , \27347 , \27348 , \27349 , \27350 ,
         \27351 , \27352 , \27353 , \27354 , \27355 , \27356 , \27357 , \27358 , \27359 , \27360 ,
         \27361 , \27362 , \27363 , \27364 , \27365 , \27366 , \27367 , \27368 , \27369 , \27370 ,
         \27371 , \27372 , \27373 , \27374 , \27375 , \27376 , \27377 , \27378 , \27379 , \27380 ,
         \27381 , \27382 , \27383 , \27384 , \27385 , \27386 , \27387 , \27388 , \27389 , \27390 ,
         \27391 , \27392 , \27393 , \27394 , \27395 , \27396 , \27397 , \27398 , \27399 , \27400 ,
         \27401 , \27402 , \27403 , \27404 , \27405 , \27406 , \27407 , \27408 , \27409 , \27410 ,
         \27411 , \27412 , \27413 , \27414 , \27415 , \27416 , \27417 , \27418 , \27419 , \27420 ,
         \27421 , \27422 , \27423 , \27424 , \27425 , \27426 , \27427 , \27428 , \27429 , \27430 ,
         \27431 , \27432 , \27433 , \27434 , \27435 , \27436 , \27437 , \27438 , \27439 , \27440 ,
         \27441 , \27442 , \27443 , \27444 , \27445 , \27446 , \27447 , \27448 , \27449 , \27450 ,
         \27451 , \27452 , \27453 , \27454 , \27455 , \27456 , \27457 , \27458 , \27459 , \27460 ,
         \27461 , \27462 , \27463 , \27464 , \27465 , \27466 , \27467 , \27468 , \27469 , \27470 ,
         \27471 , \27472 , \27473 , \27474 , \27475 , \27476 , \27477 , \27478 , \27479 , \27480 ,
         \27481 , \27482 , \27483 , \27484 , \27485 , \27486 , \27487 , \27488 , \27489 , \27490 ,
         \27491 , \27492 , \27493 , \27494 , \27495 , \27496 , \27497 , \27498 , \27499 , \27500 ,
         \27501 , \27502 , \27503 , \27504 , \27505 , \27506 , \27507 , \27508 , \27509 , \27510 ,
         \27511 , \27512 , \27513 , \27514 , \27515 , \27516 , \27517 , \27518 , \27519 , \27520 ,
         \27521 , \27522 , \27523 , \27524 , \27525 , \27526 , \27527 , \27528 , \27529 , \27530 ,
         \27531 , \27532 , \27533 , \27534 , \27535 , \27536 , \27537 , \27538 , \27539 , \27540 ,
         \27541 , \27542 , \27543 , \27544 , \27545 , \27546 , \27547 , \27548 , \27549 , \27550 ,
         \27551 , \27552 , \27553 , \27554 , \27555 , \27556 , \27557 , \27558 , \27559 , \27560 ,
         \27561 , \27562 , \27563 , \27564 , \27565 , \27566 , \27567 , \27568 , \27569 , \27570 ,
         \27571 , \27572 , \27573 , \27574 , \27575 , \27576 , \27577 , \27578 , \27579 , \27580 ,
         \27581 , \27582 , \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 ,
         \27591 , \27592 , \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 ,
         \27601 , \27602 , \27603 , \27604 , \27605 , \27606 , \27607 , \27608 , \27609 , \27610 ,
         \27611 , \27612 , \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 ,
         \27621 , \27622 , \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 ,
         \27631 , \27632 , \27633 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 ,
         \27641 , \27642 , \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 ,
         \27651 , \27652 , \27653 , \27654 , \27655 , \27656 , \27657 , \27658 , \27659 , \27660 ,
         \27661 , \27662 , \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 ,
         \27671 , \27672 , \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 ,
         \27681 , \27682 , \27683 , \27684 , \27685 , \27686 , \27687 , \27688 , \27689 , \27690 ,
         \27691 , \27692 , \27693 , \27694 , \27695 , \27696 , \27697 , \27698 , \27699 , \27700 ,
         \27701 , \27702 , \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 ,
         \27711 , \27712 , \27713 , \27714 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 ,
         \27721 , \27722 , \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 ,
         \27731 , \27732 , \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 , \27740 ,
         \27741 , \27742 , \27743 , \27744 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 ,
         \27751 , \27752 , \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 ,
         \27761 , \27762 , \27763 , \27764 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 ,
         \27771 , \27772 , \27773 , \27774 , \27775 , \27776 , \27777 , \27778 , \27779 , \27780 ,
         \27781 , \27782 , \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 ,
         \27791 , \27792 , \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 ,
         \27801 , \27802 , \27803 , \27804 , \27805 , \27806 , \27807 , \27808 , \27809 , \27810 ,
         \27811 , \27812 , \27813 , \27814 , \27815 , \27816 , \27817 , \27818 , \27819 , \27820 ,
         \27821 , \27822 , \27823 , \27824 , \27825 , \27826 , \27827 , \27828 , \27829 , \27830 ,
         \27831 , \27832 , \27833 , \27834 , \27835 , \27836 , \27837 , \27838 , \27839 , \27840 ,
         \27841 , \27842 , \27843 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 ,
         \27851 , \27852 , \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 , \27860 ,
         \27861 , \27862 , \27863 , \27864 , \27865 , \27866 , \27867 , \27868 , \27869 , \27870 ,
         \27871 , \27872 , \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 ,
         \27881 , \27882 , \27883 , \27884 , \27885 , \27886 , \27887 , \27888 , \27889 , \27890 ,
         \27891 , \27892 , \27893 , \27894 , \27895 , \27896 , \27897 , \27898 , \27899 , \27900 ,
         \27901 , \27902 , \27903 , \27904 , \27905 , \27906 , \27907 , \27908 , \27909 , \27910 ,
         \27911 , \27912 , \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 ,
         \27921 , \27922 , \27923 , \27924 , \27925 , \27926 , \27927 , \27928 , \27929 , \27930 ,
         \27931 , \27932 , \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 ,
         \27941 , \27942 , \27943 , \27944 , \27945 , \27946 , \27947 , \27948 , \27949 , \27950 ,
         \27951 , \27952 , \27953 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 ,
         \27961 , \27962 , \27963 , \27964 , \27965 , \27966 , \27967 , \27968 , \27969 , \27970 ,
         \27971 , \27972 , \27973 , \27974 , \27975 , \27976 , \27977 , \27978 , \27979 , \27980 ,
         \27981 , \27982 , \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 ,
         \27991 , \27992 , \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 ,
         \28001 , \28002 , \28003 , \28004 , \28005 , \28006 , \28007 , \28008 , \28009 , \28010 ,
         \28011 , \28012 , \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 ,
         \28021 , \28022 , \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 ,
         \28031 , \28032 , \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 ,
         \28041 , \28042 , \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 ,
         \28051 , \28052 , \28053 , \28054 , \28055 , \28056 , \28057 , \28058 , \28059 , \28060 ,
         \28061 , \28062 , \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 ,
         \28071 , \28072 , \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 ,
         \28081 , \28082 , \28083 , \28084 , \28085 , \28086 , \28087 , \28088 , \28089 , \28090 ,
         \28091 , \28092 , \28093 , \28094 , \28095 , \28096 , \28097 , \28098 , \28099 , \28100 ,
         \28101 , \28102 , \28103 , \28104 , \28105 , \28106 , \28107 , \28108 , \28109 , \28110 ,
         \28111 , \28112 , \28113 , \28114 , \28115 , \28116 , \28117 , \28118 , \28119 , \28120 ,
         \28121 , \28122 , \28123 , \28124 , \28125 , \28126 , \28127 , \28128 , \28129 , \28130 ,
         \28131 , \28132 , \28133 , \28134 , \28135 , \28136 , \28137 , \28138 , \28139 , \28140 ,
         \28141 , \28142 , \28143 , \28144 , \28145 , \28146 , \28147 , \28148 , \28149 , \28150 ,
         \28151 , \28152 , \28153 , \28154 , \28155 , \28156 , \28157 , \28158 , \28159 , \28160 ,
         \28161 , \28162 , \28163 , \28164 , \28165 , \28166 , \28167 , \28168 , \28169 , \28170 ,
         \28171 , \28172 , \28173 , \28174 , \28175 , \28176 , \28177 , \28178 , \28179 , \28180 ,
         \28181 , \28182 , \28183 , \28184 , \28185 , \28186 , \28187 , \28188 , \28189 , \28190 ,
         \28191 , \28192 , \28193 , \28194 , \28195 , \28196 , \28197 , \28198 , \28199 , \28200 ,
         \28201 , \28202 , \28203 , \28204 , \28205 , \28206 , \28207 , \28208 , \28209 , \28210 ,
         \28211 , \28212 , \28213 , \28214 , \28215 , \28216 , \28217 , \28218 , \28219 , \28220 ,
         \28221 , \28222 , \28223 , \28224 , \28225 , \28226 , \28227 , \28228 , \28229 , \28230 ,
         \28231 , \28232 , \28233 , \28234 , \28235 , \28236 , \28237 , \28238 , \28239 , \28240 ,
         \28241 , \28242 , \28243 , \28244 , \28245 , \28246 , \28247 , \28248 , \28249 , \28250 ,
         \28251 , \28252 , \28253 , \28254 , \28255 , \28256 , \28257 , \28258 , \28259 , \28260 ,
         \28261 , \28262 , \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 ,
         \28271 , \28272 , \28273 , \28274 , \28275 , \28276 , \28277 , \28278 , \28279 , \28280 ,
         \28281 , \28282 , \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 ,
         \28291 , \28292 , \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 ,
         \28301 , \28302 , \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 ,
         \28311 , \28312 , \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 ,
         \28321 , \28322 , \28323 , \28324 , \28325 , \28326 , \28327 , \28328 , \28329 , \28330 ,
         \28331 , \28332 , \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 ,
         \28341 , \28342 , \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 ,
         \28351 , \28352 , \28353 , \28354 , \28355 , \28356 , \28357 , \28358 , \28359 , \28360 ,
         \28361 , \28362 , \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 ,
         \28371 , \28372 , \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 ,
         \28381 , \28382 , \28383 , \28384 , \28385 , \28386 , \28387 , \28388 , \28389 , \28390 ,
         \28391 , \28392 , \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 ,
         \28401 , \28402 , \28403 , \28404 , \28405 , \28406 , \28407 , \28408 , \28409 , \28410 ,
         \28411 , \28412 , \28413 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 ,
         \28421 , \28422 , \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 ,
         \28431 , \28432 , \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 ,
         \28441 , \28442 , \28443 , \28444 , \28445 , \28446 , \28447 , \28448 , \28449 , \28450 ,
         \28451 , \28452 , \28453 , \28454 , \28455 , \28456 , \28457 , \28458 , \28459 , \28460 ,
         \28461 , \28462 , \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 ,
         \28471 , \28472 , \28473 , \28474 , \28475 , \28476 , \28477 , \28478 , \28479 , \28480 ,
         \28481 , \28482 , \28483 , \28484 , \28485 , \28486 , \28487 , \28488 , \28489 , \28490 ,
         \28491 , \28492 , \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 ,
         \28501 , \28502 , \28503 , \28504 , \28505 , \28506 , \28507 , \28508 , \28509 , \28510 ,
         \28511 , \28512 , \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 ,
         \28521 , \28522 , \28523 , \28524 , \28525 , \28526 , \28527 , \28528 , \28529 , \28530 ,
         \28531 , \28532 , \28533 , \28534 , \28535 , \28536 , \28537 , \28538 , \28539 , \28540 ,
         \28541 , \28542 , \28543 , \28544 , \28545 , \28546 , \28547 , \28548 , \28549 , \28550 ,
         \28551 , \28552 , \28553 , \28554 , \28555 , \28556 , \28557 , \28558 , \28559 , \28560 ,
         \28561 , \28562 , \28563 , \28564 , \28565 , \28566 , \28567 , \28568 , \28569 , \28570 ,
         \28571 , \28572 , \28573 , \28574 , \28575 , \28576 , \28577 , \28578 , \28579 , \28580 ,
         \28581 , \28582 , \28583 , \28584 , \28585 , \28586 , \28587 , \28588 , \28589 , \28590 ,
         \28591 , \28592 , \28593 , \28594 , \28595 , \28596 , \28597 , \28598 , \28599 , \28600 ,
         \28601 , \28602 , \28603 , \28604 , \28605 , \28606 , \28607 , \28608 , \28609 , \28610 ,
         \28611 , \28612 , \28613 , \28614 , \28615 , \28616 , \28617 , \28618 , \28619 , \28620 ,
         \28621 , \28622 , \28623 , \28624 , \28625 , \28626 , \28627 , \28628 , \28629 , \28630 ,
         \28631 , \28632 , \28633 , \28634 , \28635 , \28636 , \28637 , \28638 , \28639 , \28640 ,
         \28641 , \28642 , \28643 , \28644 , \28645 , \28646 , \28647 , \28648 , \28649 , \28650 ,
         \28651 , \28652 , \28653 , \28654 , \28655 , \28656 , \28657 , \28658 , \28659 , \28660 ,
         \28661 , \28662 , \28663 , \28664 , \28665 , \28666 , \28667 , \28668 , \28669 , \28670 ,
         \28671 , \28672 , \28673 , \28674 , \28675 , \28676 , \28677 , \28678 , \28679 , \28680 ,
         \28681 , \28682 , \28683 , \28684 , \28685 , \28686 , \28687 , \28688 , \28689 , \28690 ,
         \28691 , \28692 , \28693 , \28694 , \28695 , \28696 , \28697 , \28698 , \28699 , \28700 ,
         \28701 , \28702 , \28703 , \28704 , \28705 , \28706 , \28707 , \28708 , \28709 , \28710 ,
         \28711 , \28712 , \28713 , \28714 , \28715 , \28716 , \28717 , \28718 , \28719 , \28720 ,
         \28721 , \28722 , \28723 , \28724 , \28725 , \28726 , \28727 , \28728 , \28729 , \28730 ,
         \28731 , \28732 , \28733 , \28734 , \28735 , \28736 , \28737 , \28738 , \28739 , \28740 ,
         \28741 , \28742 , \28743 , \28744 , \28745 , \28746 , \28747 , \28748 , \28749 , \28750 ,
         \28751 , \28752 , \28753 , \28754 , \28755 , \28756 , \28757 , \28758 , \28759 , \28760 ,
         \28761 , \28762 , \28763 , \28764 , \28765 , \28766 , \28767 , \28768 , \28769 , \28770 ,
         \28771 , \28772 , \28773 , \28774 , \28775 , \28776 , \28777 , \28778 , \28779 , \28780 ,
         \28781 , \28782 , \28783 , \28784 , \28785 , \28786 , \28787 , \28788 , \28789 , \28790 ,
         \28791 , \28792 , \28793 , \28794 , \28795 , \28796 , \28797 , \28798 , \28799 , \28800 ,
         \28801 , \28802 , \28803 , \28804 , \28805 , \28806 , \28807 , \28808 , \28809 , \28810 ,
         \28811 , \28812 , \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 ,
         \28821 , \28822 , \28823 , \28824 , \28825 , \28826 , \28827 , \28828 , \28829 , \28830 ,
         \28831 , \28832 , \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 ,
         \28841 , \28842 , \28843 , \28844 , \28845 , \28846 , \28847 , \28848 , \28849 , \28850 ,
         \28851 , \28852 , \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , \28860 ,
         \28861 , \28862 , \28863 , \28864 , \28865 , \28866 , \28867 , \28868 , \28869 , \28870 ,
         \28871 , \28872 , \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , \28880 ,
         \28881 , \28882 , \28883 , \28884 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 ,
         \28891 , \28892 , \28893 , \28894 , \28895 , \28896 , \28897 , \28898 , \28899 , \28900 ,
         \28901 , \28902 , \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 ,
         \28911 , \28912 , \28913 , \28914 , \28915 , \28916 , \28917 , \28918 , \28919 , \28920 ,
         \28921 , \28922 , \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 ,
         \28931 , \28932 , \28933 , \28934 , \28935 , \28936 , \28937 , \28938 , \28939 , \28940 ,
         \28941 , \28942 , \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 ,
         \28951 , \28952 , \28953 , \28954 , \28955 , \28956 , \28957 , \28958 , \28959 , \28960 ,
         \28961 , \28962 , \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , \28969 , \28970 ,
         \28971 , \28972 , \28973 , \28974 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 ,
         \28981 , \28982 , \28983 , \28984 , \28985 , \28986 , \28987 , \28988 , \28989 , \28990 ,
         \28991 , \28992 , \28993 , \28994 , \28995 , \28996 , \28997 , \28998 , \28999 , \29000 ,
         \29001 , \29002 , \29003 , \29004 , \29005 , \29006 , \29007 , \29008 , \29009 , \29010 ,
         \29011 , \29012 , \29013 , \29014 , \29015 , \29016 , \29017 , \29018 , \29019 , \29020 ,
         \29021 , \29022 , \29023 , \29024 , \29025 , \29026 , \29027 , \29028 , \29029 , \29030 ,
         \29031 , \29032 , \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 ,
         \29041 , \29042 , \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 ,
         \29051 , \29052 , \29053 , \29054 , \29055 , \29056 , \29057 , \29058 , \29059 , \29060 ,
         \29061 , \29062 , \29063 , \29064 , \29065 , \29066 , \29067 , \29068 , \29069 , \29070 ,
         \29071 , \29072 , \29073 , \29074 , \29075 , \29076 , \29077 , \29078 , \29079 , \29080 ,
         \29081 , \29082 , \29083 , \29084 , \29085 , \29086 , \29087 , \29088 , \29089 , \29090 ,
         \29091 , \29092 , \29093 , \29094 , \29095 , \29096 , \29097 , \29098 , \29099 , \29100 ,
         \29101 , \29102 , \29103 , \29104 , \29105 , \29106 , \29107 , \29108 , \29109 , \29110 ,
         \29111 , \29112 , \29113 , \29114 , \29115 , \29116 , \29117 , \29118 , \29119 , \29120 ,
         \29121 , \29122 , \29123 , \29124 , \29125 , \29126 , \29127 , \29128 , \29129 , \29130 ,
         \29131 , \29132 , \29133 , \29134 , \29135 , \29136 , \29137 , \29138 , \29139 , \29140 ,
         \29141 , \29142 , \29143 , \29144 , \29145 , \29146 , \29147 , \29148 , \29149 , \29150 ,
         \29151 , \29152 , \29153 , \29154 , \29155 , \29156 , \29157 , \29158 , \29159 , \29160 ,
         \29161 , \29162 , \29163 , \29164 , \29165 , \29166 , \29167 , \29168 , \29169 , \29170 ,
         \29171 , \29172 , \29173 , \29174 , \29175 , \29176 , \29177 , \29178 , \29179 , \29180 ,
         \29181 , \29182 , \29183 , \29184 , \29185 , \29186 , \29187 , \29188 , \29189 , \29190 ,
         \29191 , \29192 , \29193 , \29194 , \29195 , \29196 , \29197 , \29198 , \29199 , \29200 ,
         \29201 , \29202 , \29203 , \29204 , \29205 , \29206 , \29207 , \29208 , \29209 , \29210 ,
         \29211 , \29212 , \29213 , \29214 , \29215 , \29216 , \29217 , \29218 , \29219 , \29220 ,
         \29221 , \29222 , \29223 , \29224 , \29225 , \29226 , \29227 , \29228 , \29229 , \29230 ,
         \29231 , \29232 , \29233 , \29234 , \29235 , \29236 , \29237 , \29238 , \29239 , \29240 ,
         \29241 , \29242 , \29243 , \29244 , \29245 , \29246 , \29247 , \29248 , \29249 , \29250 ,
         \29251 , \29252 , \29253 , \29254 , \29255 , \29256 , \29257 , \29258 , \29259 , \29260 ,
         \29261 , \29262 , \29263 , \29264 , \29265 , \29266 , \29267 , \29268 , \29269 , \29270 ,
         \29271 , \29272 , \29273 , \29274 , \29275 , \29276 , \29277 , \29278 , \29279 , \29280 ,
         \29281 , \29282 , \29283 , \29284 , \29285 , \29286 , \29287 , \29288 , \29289 , \29290 ,
         \29291 , \29292 , \29293 , \29294 , \29295 , \29296 , \29297 , \29298 , \29299 , \29300 ,
         \29301 , \29302 , \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 ,
         \29311 , \29312 , \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 ,
         \29321 , \29322 , \29323 , \29324 , \29325 , \29326 , \29327 , \29328 , \29329 , \29330 ,
         \29331 , \29332 , \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 ,
         \29341 , \29342 , \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 ,
         \29351 , \29352 , \29353 , \29354 , \29355 , \29356 , \29357 , \29358 , \29359 , \29360 ,
         \29361 , \29362 , \29363 , \29364 , \29365 , \29366 , \29367 , \29368 , \29369 , \29370 ,
         \29371 , \29372 , \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 ,
         \29381 , \29382 , \29383 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 ,
         \29391 , \29392 , \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 ,
         \29401 , \29402 , \29403 , \29404 , \29405 , \29406 , \29407 , \29408 , \29409 , \29410 ,
         \29411 , \29412 , \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 ,
         \29421 , \29422 , \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 ,
         \29431 , \29432 , \29433 , \29434 , \29435 , \29436 , \29437 , \29438 , \29439 , \29440 ,
         \29441 , \29442 , \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 ,
         \29451 , \29452 , \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 ,
         \29461 , \29462 , \29463 , \29464 , \29465 , \29466 , \29467 , \29468 , \29469 , \29470 ,
         \29471 , \29472 , \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 ,
         \29481 , \29482 , \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 ,
         \29491 , \29492 , \29493 , \29494 , \29495 , \29496 , \29497 , \29498 , \29499 , \29500 ,
         \29501 , \29502 , \29503 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 ,
         \29511 , \29512 , \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 ,
         \29521 , \29522 , \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29530 ,
         \29531 , \29532 , \29533 , \29534 , \29535 , \29536 , \29537 , \29538 , \29539 , \29540 ,
         \29541 , \29542 , \29543 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 ,
         \29551 , \29552 , \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 ,
         \29561 , \29562 , \29563 , \29564 , \29565 , \29566 , \29567 , \29568 , \29569 , \29570 ,
         \29571 , \29572 , \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 ,
         \29581 , \29582 , \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 ,
         \29591 , \29592 , \29593 , \29594 , \29595 , \29596 , \29597 , \29598 , \29599 , \29600 ,
         \29601 , \29602 , \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 ,
         \29611 , \29612 , \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 ,
         \29621 , \29622 , \29623 , \29624 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 ,
         \29631 , \29632 , \29633 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 ,
         \29641 , \29642 , \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 , \29650 ,
         \29651 , \29652 , \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 ,
         \29661 , \29662 , \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 ,
         \29671 , \29672 , \29673 , \29674 , \29675 , \29676 , \29677 , \29678 , \29679 , \29680 ,
         \29681 , \29682 , \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 ,
         \29691 , \29692 , \29693 , \29694 , \29695 , \29696 , \29697 , \29698 , \29699 , \29700 ,
         \29701 , \29702 , \29703 , \29704 , \29705 , \29706 , \29707 , \29708 , \29709 , \29710 ,
         \29711 , \29712 , \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 ,
         \29721 , \29722 , \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 ,
         \29731 , \29732 , \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 ,
         \29741 , \29742 , \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 ,
         \29751 , \29752 , \29753 , \29754 , \29755 , \29756 , \29757 , \29758 , \29759 , \29760 ,
         \29761 , \29762 , \29763 , \29764 , \29765 , \29766 , \29767 , \29768 , \29769 , \29770 ,
         \29771 , \29772 , \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 ,
         \29781 , \29782 , \29783 , \29784 , \29785 , \29786 , \29787 , \29788 , \29789 , \29790 ,
         \29791 , \29792 , \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 ,
         \29801 , \29802 , \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 ,
         \29811 , \29812 , \29813 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 ,
         \29821 , \29822 , \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 ,
         \29831 , \29832 , \29833 , \29834 , \29835 , \29836 , \29837 , \29838 , \29839 , \29840 ,
         \29841 , \29842 , \29843 , \29844 , \29845 , \29846 , \29847 , \29848 , \29849 , \29850 ,
         \29851 , \29852 , \29853 , \29854 , \29855 , \29856 , \29857 , \29858 , \29859 , \29860 ,
         \29861 , \29862 , \29863 , \29864 , \29865 , \29866 , \29867 , \29868 , \29869 , \29870 ,
         \29871 , \29872 , \29873 , \29874 , \29875 , \29876 , \29877 , \29878 , \29879 , \29880 ,
         \29881 , \29882 , \29883 , \29884 , \29885 , \29886 , \29887 , \29888 , \29889 , \29890 ,
         \29891 , \29892 , \29893 , \29894 , \29895 , \29896 , \29897 , \29898 , \29899 , \29900 ,
         \29901 , \29902 , \29903 , \29904 , \29905 , \29906 , \29907 , \29908 , \29909 , \29910 ,
         \29911 , \29912 , \29913 , \29914 , \29915 , \29916 , \29917 , \29918 , \29919 , \29920 ,
         \29921 , \29922 , \29923 , \29924 , \29925 , \29926 , \29927 , \29928 , \29929 , \29930 ,
         \29931 , \29932 , \29933 , \29934 , \29935 , \29936 , \29937 , \29938 , \29939 , \29940 ,
         \29941 , \29942 , \29943 , \29944 , \29945 , \29946 , \29947 , \29948 , \29949 , \29950 ,
         \29951 , \29952 , \29953 , \29954 , \29955 , \29956 , \29957 , \29958 , \29959 , \29960 ,
         \29961 , \29962 , \29963 , \29964 , \29965 , \29966 , \29967 , \29968 , \29969 , \29970 ,
         \29971 , \29972 , \29973 , \29974 , \29975 , \29976 , \29977 , \29978 , \29979 , \29980 ,
         \29981 , \29982 , \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 ,
         \29991 , \29992 , \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 ,
         \30001 , \30002 , \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 , \30010 ,
         \30011 , \30012 , \30013 , \30014 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 ,
         \30021 , \30022 , \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 ,
         \30031 , \30032 , \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 ,
         \30041 , \30042 , \30043 , \30044 , \30045 , \30046 , \30047 , \30048 , \30049 , \30050 ,
         \30051 , \30052 , \30053 , \30054 , \30055 , \30056 , \30057 , \30058 , \30059 , \30060 ,
         \30061 , \30062 , \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 ,
         \30071 , \30072 , \30073 , \30074 , \30075 , \30076 , \30077 , \30078 , \30079 , \30080 ,
         \30081 , \30082 , \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 ,
         \30091 , \30092 , \30093 , \30094 , \30095 , \30096 , \30097 , \30098 , \30099 , \30100 ,
         \30101 , \30102 , \30103 , \30104 , \30105 , \30106 , \30107 , \30108 , \30109 , \30110 ,
         \30111 , \30112 , \30113 , \30114 , \30115 , \30116 , \30117 , \30118 , \30119 , \30120 ,
         \30121 , \30122 , \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 ,
         \30131 , \30132 , \30133 , \30134 , \30135 , \30136 , \30137 , \30138 , \30139 , \30140 ,
         \30141 , \30142 , \30143 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 ,
         \30151 , \30152 , \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 , \30160 ,
         \30161 , \30162 , \30163 , \30164 , \30165 , \30166 , \30167 , \30168 , \30169 , \30170 ,
         \30171 , \30172 , \30173 , \30174 , \30175 , \30176 , \30177 , \30178 , \30179 , \30180 ,
         \30181 , \30182 , \30183 , \30184 , \30185 , \30186 , \30187 , \30188 , \30189 , \30190 ,
         \30191 , \30192 , \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 ,
         \30201 , \30202 , \30203 , \30204 , \30205 , \30206 , \30207 , \30208 , \30209 , \30210 ,
         \30211 , \30212 , \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 ,
         \30221 , \30222 , \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 ,
         \30231 , \30232 , \30233 , \30234 , \30235 , \30236 , \30237 , \30238 , \30239 , \30240 ,
         \30241 , \30242 , \30243 , \30244 , \30245 , \30246 , \30247 , \30248 , \30249 , \30250 ,
         \30251 , \30252 , \30253 , \30254 , \30255 , \30256 , \30257 , \30258 , \30259 , \30260 ,
         \30261 , \30262 , \30263 , \30264 , \30265 , \30266 , \30267 , \30268 , \30269 , \30270 ,
         \30271 , \30272 , \30273 , \30274 , \30275 , \30276 , \30277 , \30278 , \30279 , \30280 ,
         \30281 , \30282 , \30283 , \30284 , \30285 , \30286 , \30287 , \30288 , \30289 , \30290 ,
         \30291 , \30292 , \30293 , \30294 , \30295 , \30296 , \30297 , \30298 , \30299 , \30300 ,
         \30301 , \30302 , \30303 , \30304 , \30305 , \30306 , \30307 , \30308 , \30309 , \30310 ,
         \30311 , \30312 , \30313 , \30314 , \30315 , \30316 , \30317 , \30318 , \30319 , \30320 ,
         \30321 , \30322 , \30323 , \30324 , \30325 , \30326 , \30327 , \30328 , \30329 , \30330 ,
         \30331 , \30332 , \30333 , \30334 , \30335 , \30336 , \30337 , \30338 , \30339 , \30340 ,
         \30341 , \30342 , \30343 , \30344 , \30345 , \30346 , \30347 , \30348 , \30349 , \30350 ,
         \30351 , \30352 , \30353 , \30354 , \30355 , \30356 , \30357 , \30358 , \30359 , \30360 ,
         \30361 , \30362 , \30363 , \30364 , \30365 , \30366 , \30367 , \30368 , \30369 , \30370 ,
         \30371 , \30372 , \30373 , \30374 , \30375 , \30376 , \30377 , \30378 , \30379 , \30380 ,
         \30381 , \30382 , \30383 , \30384 , \30385 , \30386 , \30387 , \30388 , \30389 , \30390 ,
         \30391 , \30392 , \30393 , \30394 , \30395 , \30396 , \30397 , \30398 , \30399 , \30400 ,
         \30401 , \30402 , \30403 , \30404 , \30405 , \30406 , \30407 , \30408 , \30409 , \30410 ,
         \30411 , \30412 , \30413 , \30414 , \30415 , \30416 , \30417 , \30418 , \30419 , \30420 ,
         \30421 , \30422 , \30423 , \30424 , \30425 , \30426 , \30427 , \30428 , \30429 , \30430 ,
         \30431 , \30432 , \30433 , \30434 , \30435 , \30436 , \30437 , \30438 , \30439 , \30440 ,
         \30441 , \30442 , \30443 , \30444 , \30445 , \30446 , \30447 , \30448 , \30449 , \30450 ,
         \30451 , \30452 , \30453 , \30454 , \30455 , \30456 , \30457 , \30458 , \30459 , \30460 ,
         \30461 , \30462 , \30463 , \30464 , \30465 , \30466 , \30467 , \30468 , \30469 , \30470 ,
         \30471 , \30472 , \30473 , \30474 , \30475 , \30476 , \30477 , \30478 , \30479 , \30480 ,
         \30481 , \30482 , \30483 , \30484 , \30485 , \30486 , \30487 , \30488 , \30489 , \30490 ,
         \30491 , \30492 , \30493 , \30494 , \30495 , \30496 , \30497 , \30498 , \30499 , \30500 ,
         \30501 , \30502 , \30503 , \30504 , \30505 , \30506 , \30507 , \30508 , \30509 , \30510 ,
         \30511 , \30512 , \30513 , \30514 , \30515 , \30516 , \30517 , \30518 , \30519 , \30520 ,
         \30521 , \30522 , \30523 , \30524 , \30525 , \30526 , \30527 , \30528 , \30529 , \30530 ,
         \30531 , \30532 , \30533 , \30534 , \30535 , \30536 , \30537 , \30538 , \30539 , \30540 ,
         \30541 , \30542 , \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 ,
         \30551 , \30552 , \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 ,
         \30561 , \30562 , \30563 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 ,
         \30571 , \30572 , \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 ,
         \30581 , \30582 , \30583 , \30584 , \30585 , \30586 , \30587 , \30588 , \30589 , \30590 ,
         \30591 , \30592 , \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 ,
         \30601 , \30602 , \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 ,
         \30611 , \30612 , \30613 , \30614 , \30615 , \30616 , \30617 , \30618 , \30619 , \30620 ,
         \30621 , \30622 , \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 ,
         \30631 , \30632 , \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 ,
         \30641 , \30642 , \30643 , \30644 , \30645 , \30646 , \30647 , \30648 , \30649 , \30650 ,
         \30651 , \30652 , \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 ,
         \30661 , \30662 , \30663 , \30664 , \30665 , \30666 , \30667 , \30668 , \30669 , \30670 ,
         \30671 , \30672 , \30673 , \30674 , \30675 , \30676 , \30677 , \30678 , \30679 , \30680 ,
         \30681 , \30682 , \30683 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 ,
         \30691 , \30692 , \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 ,
         \30701 , \30702 , \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30710 ,
         \30711 , \30712 , \30713 , \30714 , \30715 , \30716 , \30717 , \30718 , \30719 , \30720 ,
         \30721 , \30722 , \30723 , \30724 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 ,
         \30731 , \30732 , \30733 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 ,
         \30741 , \30742 , \30743 , \30744 , \30745 , \30746 , \30747 , \30748 , \30749 , \30750 ,
         \30751 , \30752 , \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 ,
         \30761 , \30762 , \30763 , \30764 , \30765 , \30766 , \30767 , \30768 , \30769 , \30770 ,
         \30771 , \30772 , \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 ,
         \30781 , \30782 , \30783 , \30784 , \30785 , \30786 , \30787 , \30788 , \30789 , \30790 ,
         \30791 , \30792 , \30793 , \30794 , \30795 , \30796 , \30797 , \30798 , \30799 , \30800 ,
         \30801 , \30802 , \30803 , \30804 , \30805 , \30806 , \30807 , \30808 , \30809 , \30810 ,
         \30811 , \30812 , \30813 , \30814 , \30815 , \30816 , \30817 , \30818 , \30819 , \30820 ,
         \30821 , \30822 , \30823 , \30824 , \30825 , \30826 , \30827 , \30828 , \30829 , \30830 ,
         \30831 , \30832 , \30833 , \30834 , \30835 , \30836 , \30837 , \30838 , \30839 , \30840 ,
         \30841 , \30842 , \30843 , \30844 , \30845 , \30846 , \30847 , \30848 , \30849 , \30850 ,
         \30851 , \30852 , \30853 , \30854 , \30855 , \30856 , \30857 , \30858 , \30859 , \30860 ,
         \30861 , \30862 , \30863 , \30864 , \30865 , \30866 , \30867 , \30868 , \30869 , \30870 ,
         \30871 , \30872 , \30873 , \30874 , \30875 , \30876 , \30877 , \30878 , \30879 , \30880 ,
         \30881 , \30882 , \30883 , \30884 , \30885 , \30886 , \30887 , \30888 , \30889 , \30890 ,
         \30891 , \30892 , \30893 , \30894 , \30895 , \30896 , \30897 , \30898 , \30899 , \30900 ,
         \30901 , \30902 , \30903 , \30904 , \30905 , \30906 , \30907 , \30908 , \30909 , \30910 ,
         \30911 , \30912 , \30913 , \30914 , \30915 , \30916 , \30917 , \30918 , \30919 , \30920 ,
         \30921 , \30922 , \30923 , \30924 , \30925 , \30926 , \30927 , \30928 , \30929 , \30930 ,
         \30931 , \30932 , \30933 , \30934 , \30935 , \30936 , \30937 , \30938 , \30939 , \30940 ,
         \30941 , \30942 , \30943 , \30944 , \30945 , \30946 , \30947 , \30948 , \30949 , \30950 ,
         \30951 , \30952 , \30953 , \30954 , \30955 , \30956 , \30957 , \30958 , \30959 , \30960 ,
         \30961 , \30962 , \30963 , \30964 , \30965 , \30966 , \30967 , \30968 , \30969 , \30970 ,
         \30971 , \30972 , \30973 , \30974 , \30975 , \30976 , \30977 , \30978 , \30979 , \30980 ,
         \30981 , \30982 , \30983 , \30984 , \30985 , \30986 , \30987 , \30988 , \30989 , \30990 ,
         \30991 , \30992 , \30993 , \30994 , \30995 , \30996 , \30997 , \30998 , \30999 , \31000 ,
         \31001 , \31002 , \31003 , \31004 , \31005 , \31006 , \31007 , \31008 , \31009 , \31010 ,
         \31011 , \31012 , \31013 , \31014 , \31015 , \31016 , \31017 , \31018 , \31019 , \31020 ,
         \31021 , \31022 , \31023 , \31024 , \31025 , \31026 , \31027 , \31028 , \31029 , \31030 ,
         \31031 , \31032 , \31033 , \31034 , \31035 , \31036 , \31037 , \31038 , \31039 , \31040 ,
         \31041 , \31042 , \31043 , \31044 , \31045 , \31046 , \31047 , \31048 , \31049 , \31050 ,
         \31051 , \31052 , \31053 , \31054 , \31055 , \31056 , \31057 , \31058 , \31059 , \31060 ,
         \31061 , \31062 , \31063 , \31064 , \31065 , \31066 , \31067 , \31068 , \31069 , \31070 ,
         \31071 , \31072 , \31073 , \31074 , \31075 , \31076 , \31077 , \31078 , \31079 , \31080 ,
         \31081 , \31082 , \31083 , \31084 , \31085 , \31086 , \31087 , \31088 , \31089 , \31090 ,
         \31091 , \31092 , \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , \31100 ,
         \31101 , \31102 , \31103 , \31104 , \31105 , \31106 , \31107 , \31108 , \31109 , \31110 ,
         \31111 , \31112 , \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 ,
         \31121 , \31122 , \31123 , \31124 , \31125 , \31126 , \31127 , \31128 , \31129 , \31130 ,
         \31131 , \31132 , \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , \31139 , \31140 ,
         \31141 , \31142 , \31143 , \31144 , \31145 , \31146 , \31147 , \31148 , \31149 , \31150 ,
         \31151 , \31152 , \31153 , \31154 , \31155 , \31156 , \31157 , \31158 , \31159 , \31160 ,
         \31161 , \31162 , \31163 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 ,
         \31171 , \31172 , \31173 , \31174 , \31175 , \31176 , \31177 , \31178 , \31179 , \31180 ,
         \31181 , \31182 , \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 ,
         \31191 , \31192 , \31193 , \31194 , \31195 , \31196 , \31197 , \31198 , \31199 , \31200 ,
         \31201 , \31202 , \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 ,
         \31211 , \31212 , \31213 , \31214 , \31215 , \31216 , \31217 , \31218 , \31219 , \31220 ,
         \31221 , \31222 , \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 ,
         \31231 , \31232 , \31233 , \31234 , \31235 , \31236 , \31237 , \31238 , \31239 , \31240 ,
         \31241 , \31242 , \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 ,
         \31251 , \31252 , \31253 , \31254 , \31255 , \31256 , \31257 , \31258 , \31259 , \31260 ,
         \31261 , \31262 , \31263 , \31264 , \31265 , \31266 , \31267 , \31268 , \31269 , \31270 ,
         \31271 , \31272 , \31273 , \31274 , \31275 , \31276 , \31277 , \31278 , \31279 , \31280 ,
         \31281 , \31282 , \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 ,
         \31291 , \31292 , \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 ,
         \31301 , \31302 , \31303 , \31304 , \31305 , \31306 , \31307 , \31308 , \31309 , \31310 ,
         \31311 , \31312 , \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 ,
         \31321 , \31322 , \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 ,
         \31331 , \31332 , \31333 , \31334 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 ,
         \31341 , \31342 , \31343 , \31344 , \31345 , \31346 , \31347 , \31348 , \31349 , \31350 ,
         \31351 , \31352 , \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 , \31360 ,
         \31361 , \31362 , \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 ,
         \31371 , \31372 , \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 ,
         \31381 , \31382 , \31383 , \31384 , \31385 , \31386 , \31387 , \31388 , \31389 , \31390 ,
         \31391 , \31392 , \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 ,
         \31401 , \31402 , \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 ,
         \31411 , \31412 , \31413 , \31414 , \31415 , \31416 , \31417 , \31418 , \31419 , \31420 ,
         \31421 , \31422 , \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 ,
         \31431 , \31432 , \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 ,
         \31441 , \31442 , \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 ,
         \31451 , \31452 , \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 ,
         \31461 , \31462 , \31463 , \31464 , \31465 , \31466 , \31467 , \31468 , \31469 , \31470 ,
         \31471 , \31472 , \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 ,
         \31481 , \31482 , \31483 , \31484 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 ,
         \31491 , \31492 , \31493 , \31494 , \31495 , \31496 , \31497 , \31498 , \31499 , \31500 ,
         \31501 , \31502 , \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 ,
         \31511 , \31512 , \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 ,
         \31521 , \31522 , \31523 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 ,
         \31531 , \31532 , \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 ,
         \31541 , \31542 , \31543 , \31544 , \31545 , \31546 , \31547 , \31548 , \31549 , \31550 ,
         \31551 , \31552 , \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 ,
         \31561 , \31562 , \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 ,
         \31571 , \31572 , \31573 , \31574 , \31575 , \31576 , \31577 , \31578 , \31579 , \31580 ,
         \31581 , \31582 , \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 ,
         \31591 , \31592 , \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 ,
         \31601 , \31602 , \31603 , \31604 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 ,
         \31611 , \31612 , \31613 , \31614 , \31615 , \31616 , \31617 , \31618 , \31619 , \31620 ,
         \31621 , \31622 , \31623 , \31624 , \31625 , \31626 , \31627 , \31628 , \31629 , \31630 ,
         \31631 , \31632 , \31633 , \31634 , \31635 , \31636 , \31637 , \31638 , \31639 , \31640 ,
         \31641 , \31642 , \31643 , \31644 , \31645 , \31646 , \31647 , \31648 , \31649 , \31650 ,
         \31651 , \31652 , \31653 , \31654 , \31655 , \31656 , \31657 , \31658 , \31659 , \31660 ,
         \31661 , \31662 , \31663 , \31664 , \31665 , \31666 , \31667 , \31668 , \31669 , \31670 ,
         \31671 , \31672 , \31673 , \31674 , \31675 , \31676 , \31677 , \31678 , \31679 , \31680 ,
         \31681 , \31682 , \31683 , \31684 , \31685 , \31686 , \31687 , \31688 , \31689 , \31690 ,
         \31691 , \31692 , \31693 , \31694 , \31695 , \31696 , \31697 , \31698 , \31699 , \31700 ,
         \31701 , \31702 , \31703 , \31704 , \31705 , \31706 , \31707 , \31708 , \31709 , \31710 ,
         \31711 , \31712 , \31713 , \31714 , \31715 , \31716 , \31717 , \31718 , \31719 , \31720 ,
         \31721 , \31722 , \31723 , \31724 , \31725 , \31726 , \31727 , \31728 , \31729 , \31730 ,
         \31731 , \31732 , \31733 , \31734 , \31735 , \31736 , \31737 , \31738 , \31739 , \31740 ,
         \31741 , \31742 , \31743 , \31744 , \31745 , \31746 , \31747 , \31748 , \31749 , \31750 ,
         \31751 , \31752 , \31753 , \31754 , \31755 , \31756 , \31757 , \31758 , \31759 , \31760 ,
         \31761 , \31762 , \31763 , \31764 , \31765 , \31766 , \31767 , \31768 , \31769 , \31770 ,
         \31771 , \31772 , \31773 , \31774 , \31775 , \31776 , \31777 , \31778 , \31779 , \31780 ,
         \31781 , \31782 , \31783 , \31784 , \31785 , \31786 , \31787 , \31788 , \31789 , \31790 ,
         \31791 , \31792 , \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 ,
         \31801 , \31802 , \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 ,
         \31811 , \31812 , \31813 , \31814 , \31815 , \31816 , \31817 , \31818 , \31819 , \31820 ,
         \31821 , \31822 , \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 ,
         \31831 , \31832 , \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 ,
         \31841 , \31842 , \31843 , \31844 , \31845 , \31846 , \31847 , \31848 , \31849 , \31850 ,
         \31851 , \31852 , \31853 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 ,
         \31861 , \31862 , \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 ,
         \31871 , \31872 , \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 ,
         \31881 , \31882 , \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 ,
         \31891 , \31892 , \31893 , \31894 , \31895 , \31896 , \31897 , \31898 , \31899 , \31900 ,
         \31901 , \31902 , \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 ,
         \31911 , \31912 , \31913 , \31914 , \31915 , \31916 , \31917 , \31918 , \31919 , \31920 ,
         \31921 , \31922 , \31923 , \31924 , \31925 , \31926 , \31927 , \31928 , \31929 , \31930 ,
         \31931 , \31932 , \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 ,
         \31941 , \31942 , \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 ,
         \31951 , \31952 , \31953 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 ,
         \31961 , \31962 , \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 ,
         \31971 , \31972 , \31973 , \31974 , \31975 , \31976 , \31977 , \31978 , \31979 , \31980 ,
         \31981 , \31982 , \31983 , \31984 , \31985 , \31986 , \31987 , \31988 , \31989 , \31990 ,
         \31991 , \31992 , \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 ,
         \32001 , \32002 , \32003 , \32004 , \32005 , \32006 , \32007 , \32008 , \32009 , \32010 ,
         \32011 , \32012 , \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 ,
         \32021 , \32022 , \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 ,
         \32031 , \32032 , \32033 , \32034 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 ,
         \32041 , \32042 , \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 , \32050 ,
         \32051 , \32052 , \32053 , \32054 , \32055 , \32056 , \32057 , \32058 , \32059 , \32060 ,
         \32061 , \32062 , \32063 , \32064 , \32065 , \32066 , \32067 , \32068 , \32069 , \32070 ,
         \32071 , \32072 , \32073 , \32074 , \32075 , \32076 , \32077 , \32078 , \32079 , \32080 ,
         \32081 , \32082 , \32083 , \32084 , \32085 , \32086 , \32087 , \32088 , \32089 , \32090 ,
         \32091 , \32092 , \32093 , \32094 , \32095 , \32096 , \32097 , \32098 , \32099 , \32100 ,
         \32101 , \32102 , \32103 , \32104 , \32105 , \32106 , \32107 , \32108 , \32109 , \32110 ,
         \32111 , \32112 , \32113 , \32114 , \32115 , \32116 , \32117 , \32118 , \32119 , \32120 ,
         \32121 , \32122 , \32123 , \32124 , \32125 , \32126 , \32127 , \32128 , \32129 , \32130 ,
         \32131 , \32132 , \32133 , \32134 , \32135 , \32136 , \32137 , \32138 , \32139 , \32140 ,
         \32141 , \32142 , \32143 , \32144 , \32145 , \32146 , \32147 , \32148 , \32149 , \32150 ,
         \32151 , \32152 , \32153 , \32154 , \32155 , \32156 , \32157 , \32158 , \32159 , \32160 ,
         \32161 , \32162 , \32163 , \32164 , \32165 , \32166 , \32167 , \32168 , \32169 , \32170 ,
         \32171 , \32172 , \32173 , \32174 , \32175 , \32176 , \32177 , \32178 , \32179 , \32180 ,
         \32181 , \32182 , \32183 , \32184 , \32185 , \32186 , \32187 , \32188 , \32189 , \32190 ,
         \32191 , \32192 , \32193 , \32194 , \32195 , \32196 , \32197 , \32198 , \32199 , \32200 ,
         \32201 , \32202 , \32203 , \32204 , \32205 , \32206 , \32207 , \32208 , \32209 , \32210 ,
         \32211 , \32212 , \32213 , \32214 , \32215 , \32216 , \32217 , \32218 , \32219 , \32220 ,
         \32221 , \32222 , \32223 , \32224 , \32225 , \32226 , \32227 , \32228 , \32229 , \32230 ,
         \32231 , \32232 , \32233 , \32234 , \32235 , \32236 , \32237 , \32238 , \32239 , \32240 ,
         \32241 , \32242 , \32243 , \32244 , \32245 , \32246 , \32247 , \32248 , \32249 , \32250 ,
         \32251 , \32252 , \32253 , \32254 , \32255 , \32256 , \32257 , \32258 , \32259 , \32260 ,
         \32261 , \32262 , \32263 , \32264 , \32265 , \32266 , \32267 , \32268 , \32269 , \32270 ,
         \32271 , \32272 , \32273 , \32274 , \32275 , \32276 , \32277 , \32278 , \32279 , \32280 ,
         \32281 , \32282 , \32283 , \32284 , \32285 , \32286 , \32287 , \32288 , \32289 , \32290 ,
         \32291 , \32292 , \32293 , \32294 , \32295 , \32296 , \32297 , \32298 , \32299 , \32300 ,
         \32301 , \32302 , \32303 , \32304 , \32305 , \32306 , \32307 , \32308 , \32309 , \32310 ,
         \32311 , \32312 , \32313 , \32314 , \32315 , \32316 , \32317 , \32318 , \32319 , \32320 ,
         \32321 , \32322 , \32323 , \32324 , \32325 , \32326 , \32327 , \32328 , \32329 , \32330 ,
         \32331 , \32332 , \32333 , \32334 , \32335 , \32336 , \32337 , \32338 , \32339 , \32340 ,
         \32341 , \32342 , \32343 , \32344 , \32345 , \32346 , \32347 , \32348 , \32349 , \32350 ,
         \32351 , \32352 , \32353 , \32354 , \32355 , \32356 , \32357 , \32358 , \32359 , \32360 ,
         \32361 , \32362 , \32363 , \32364 , \32365 , \32366 , \32367 , \32368 , \32369 , \32370 ,
         \32371 , \32372 , \32373 , \32374 , \32375 , \32376 , \32377 , \32378 , \32379 , \32380 ,
         \32381 , \32382 , \32383 , \32384 , \32385 , \32386 , \32387 , \32388 , \32389 , \32390 ,
         \32391 , \32392 , \32393 , \32394 , \32395 , \32396 , \32397 , \32398 , \32399 , \32400 ,
         \32401 , \32402 , \32403 , \32404 , \32405 , \32406 , \32407 , \32408 , \32409 , \32410 ,
         \32411 , \32412 , \32413 , \32414 , \32415 , \32416 , \32417 , \32418 , \32419 , \32420 ,
         \32421 , \32422 , \32423 , \32424 , \32425 , \32426 , \32427 , \32428 , \32429 , \32430 ,
         \32431 , \32432 , \32433 , \32434 , \32435 , \32436 , \32437 , \32438 , \32439 , \32440 ,
         \32441 , \32442 , \32443 , \32444 , \32445 , \32446 , \32447 , \32448 , \32449 , \32450 ,
         \32451 , \32452 , \32453 , \32454 , \32455 , \32456 , \32457 , \32458 , \32459 , \32460 ,
         \32461 , \32462 , \32463 , \32464 , \32465 , \32466 , \32467 , \32468 , \32469 , \32470 ,
         \32471 , \32472 , \32473 , \32474 , \32475 , \32476 , \32477 , \32478 , \32479 , \32480 ,
         \32481 , \32482 , \32483 , \32484 , \32485 , \32486 , \32487 , \32488 , \32489 , \32490 ,
         \32491 , \32492 , \32493 , \32494 , \32495 , \32496 , \32497 , \32498 , \32499 , \32500 ,
         \32501 , \32502 , \32503 , \32504 , \32505 , \32506 , \32507 , \32508 , \32509 , \32510 ,
         \32511 , \32512 , \32513 , \32514 , \32515 , \32516 , \32517 , \32518 , \32519 , \32520 ,
         \32521 , \32522 , \32523 , \32524 , \32525 , \32526 , \32527 , \32528 , \32529 , \32530 ,
         \32531 , \32532 , \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 , \32540 ,
         \32541 , \32542 , \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 ,
         \32551 , \32552 , \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 ,
         \32561 , \32562 , \32563 , \32564 , \32565 , \32566 , \32567 , \32568 , \32569 , \32570 ,
         \32571 , \32572 , \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 ,
         \32581 , \32582 , \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 ,
         \32591 , \32592 , \32593 , \32594 , \32595 , \32596 , \32597 , \32598 , \32599 , \32600 ,
         \32601 , \32602 , \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 ,
         \32611 , \32612 , \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 ,
         \32621 , \32622 , \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 ,
         \32631 , \32632 , \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 ,
         \32641 , \32642 , \32643 , \32644 , \32645 , \32646 , \32647 , \32648 , \32649 , \32650 ,
         \32651 , \32652 , \32653 , \32654 , \32655 , \32656 , \32657 , \32658 , \32659 , \32660 ,
         \32661 , \32662 , \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 ,
         \32671 , \32672 , \32673 , \32674 , \32675 , \32676 , \32677 , \32678 , \32679 , \32680 ,
         \32681 , \32682 , \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 ,
         \32691 , \32692 , \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 ,
         \32701 , \32702 , \32703 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 ,
         \32711 , \32712 , \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 ,
         \32721 , \32722 , \32723 , \32724 , \32725 , \32726 , \32727 , \32728 , \32729 , \32730 ,
         \32731 , \32732 , \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 ,
         \32741 , \32742 , \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 ,
         \32751 , \32752 , \32753 , \32754 , \32755 , \32756 , \32757 , \32758 , \32759 , \32760 ,
         \32761 , \32762 , \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 ,
         \32771 , \32772 , \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 ,
         \32781 , \32782 , \32783 , \32784 , \32785 , \32786 , \32787 , \32788 , \32789 , \32790 ,
         \32791 , \32792 , \32793 , \32794 , \32795 , \32796 , \32797 , \32798 , \32799 , \32800 ,
         \32801 , \32802 , \32803 , \32804 , \32805 , \32806 , \32807 , \32808 , \32809 , \32810 ,
         \32811 , \32812 , \32813 , \32814 , \32815 , \32816 , \32817 , \32818 , \32819 , \32820 ,
         \32821 , \32822 , \32823 , \32824 , \32825 , \32826 , \32827 , \32828 , \32829 , \32830 ,
         \32831 , \32832 , \32833 , \32834 , \32835 , \32836 , \32837 , \32838 , \32839 , \32840 ,
         \32841 , \32842 , \32843 , \32844 , \32845 , \32846 , \32847 , \32848 , \32849 , \32850 ,
         \32851 , \32852 , \32853 , \32854 , \32855 , \32856 , \32857 , \32858 , \32859 , \32860 ,
         \32861 , \32862 , \32863 , \32864 , \32865 , \32866 , \32867 , \32868 , \32869 , \32870 ,
         \32871 , \32872 , \32873 , \32874 , \32875 , \32876 , \32877 , \32878 , \32879 , \32880 ,
         \32881 , \32882 , \32883 , \32884 , \32885 , \32886 , \32887 , \32888 , \32889 , \32890 ,
         \32891 , \32892 , \32893 , \32894 , \32895 , \32896 , \32897 , \32898 , \32899 , \32900 ,
         \32901 , \32902 , \32903 , \32904 , \32905 , \32906 , \32907 , \32908 , \32909 , \32910 ,
         \32911 , \32912 , \32913 , \32914 , \32915 , \32916 , \32917 , \32918 , \32919 , \32920 ,
         \32921 , \32922 , \32923 , \32924 , \32925 , \32926 , \32927 , \32928 , \32929 , \32930 ,
         \32931 , \32932 , \32933 , \32934 , \32935 , \32936 , \32937 , \32938 , \32939 , \32940 ,
         \32941 , \32942 , \32943 , \32944 , \32945 , \32946 , \32947 , \32948 , \32949 , \32950 ,
         \32951 , \32952 , \32953 , \32954 , \32955 , \32956 , \32957 , \32958 , \32959 , \32960 ,
         \32961 , \32962 , \32963 , \32964 , \32965 , \32966 , \32967 , \32968 , \32969 , \32970 ,
         \32971 , \32972 , \32973 , \32974 , \32975 , \32976 , \32977 , \32978 , \32979 , \32980 ,
         \32981 , \32982 , \32983 , \32984 , \32985 , \32986 , \32987 , \32988 , \32989 , \32990 ,
         \32991 , \32992 , \32993 , \32994 , \32995 , \32996 , \32997 , \32998 , \32999 , \33000 ,
         \33001 , \33002 , \33003 , \33004 , \33005 , \33006 , \33007 , \33008 , \33009 , \33010 ,
         \33011 , \33012 , \33013 , \33014 , \33015 , \33016 , \33017 , \33018 , \33019 , \33020 ,
         \33021 , \33022 , \33023 , \33024 , \33025 , \33026 , \33027 , \33028 , \33029 , \33030 ,
         \33031 , \33032 , \33033 , \33034 , \33035 , \33036 , \33037 , \33038 , \33039 , \33040 ,
         \33041 , \33042 , \33043 , \33044 , \33045 , \33046 , \33047 , \33048 , \33049 , \33050 ,
         \33051 , \33052 , \33053 , \33054 , \33055 , \33056 , \33057 , \33058 , \33059 , \33060 ,
         \33061 , \33062 , \33063 , \33064 , \33065 , \33066 , \33067 , \33068 , \33069 , \33070 ,
         \33071 , \33072 , \33073 , \33074 , \33075 , \33076 , \33077 , \33078 , \33079 , \33080 ,
         \33081 , \33082 , \33083 , \33084 , \33085 , \33086 , \33087 , \33088 , \33089 , \33090 ,
         \33091 , \33092 , \33093 , \33094 , \33095 , \33096 , \33097 , \33098 , \33099 , \33100 ,
         \33101 , \33102 , \33103 , \33104 , \33105 , \33106 , \33107 , \33108 , \33109 , \33110 ,
         \33111 , \33112 , \33113 , \33114 , \33115 , \33116 , \33117 , \33118 , \33119 , \33120 ,
         \33121 , \33122 , \33123 , \33124 , \33125 , \33126 , \33127 , \33128 , \33129 , \33130 ,
         \33131 , \33132 , \33133 , \33134 , \33135 , \33136 , \33137 , \33138 , \33139 , \33140 ,
         \33141 , \33142 , \33143 , \33144 , \33145 , \33146 , \33147 , \33148 , \33149 , \33150 ,
         \33151 , \33152 , \33153 , \33154 , \33155 , \33156 , \33157 , \33158 , \33159 , \33160 ,
         \33161 , \33162 , \33163 , \33164 , \33165 , \33166 , \33167 , \33168 , \33169 , \33170 ,
         \33171 , \33172 , \33173 , \33174 , \33175 , \33176 , \33177 , \33178 , \33179 , \33180 ,
         \33181 , \33182 , \33183 , \33184 , \33185 , \33186 , \33187 , \33188 , \33189 , \33190 ,
         \33191 , \33192 , \33193 , \33194 , \33195 , \33196 , \33197 , \33198 , \33199 , \33200 ,
         \33201 , \33202 , \33203 , \33204 , \33205 , \33206 , \33207 , \33208 , \33209 , \33210 ,
         \33211 , \33212 , \33213 , \33214 , \33215 , \33216 , \33217 , \33218 , \33219 , \33220 ,
         \33221 , \33222 , \33223 , \33224 , \33225 , \33226 , \33227 , \33228 , \33229 , \33230 ,
         \33231 , \33232 , \33233 , \33234 , \33235 , \33236 , \33237 , \33238 , \33239 , \33240 ,
         \33241 , \33242 , \33243 , \33244 , \33245 , \33246 , \33247 , \33248 , \33249 , \33250 ,
         \33251 , \33252 , \33253 , \33254 , \33255 , \33256 , \33257 , \33258 , \33259 , \33260 ,
         \33261 , \33262 , \33263 , \33264 , \33265 , \33266 , \33267 , \33268 , \33269 , \33270 ,
         \33271 , \33272 , \33273 , \33274 , \33275 , \33276 , \33277 , \33278 , \33279 , \33280 ,
         \33281 , \33282 , \33283 , \33284 , \33285 , \33286 , \33287 , \33288 , \33289 , \33290 ,
         \33291 , \33292 , \33293 , \33294 , \33295 , \33296 , \33297 , \33298 , \33299 , \33300 ,
         \33301 , \33302 , \33303 , \33304 , \33305 , \33306 , \33307 , \33308 , \33309 , \33310 ,
         \33311 , \33312 , \33313 , \33314 , \33315 , \33316 , \33317 , \33318 , \33319 , \33320 ,
         \33321 , \33322 , \33323 , \33324 , \33325 , \33326 , \33327 , \33328 , \33329 , \33330 ,
         \33331 , \33332 , \33333 , \33334 , \33335 , \33336 , \33337 , \33338 , \33339 , \33340 ,
         \33341 , \33342 , \33343 , \33344 , \33345 , \33346 , \33347 , \33348 , \33349 , \33350 ,
         \33351 , \33352 , \33353 , \33354 , \33355 , \33356 , \33357 , \33358 , \33359 , \33360 ,
         \33361 , \33362 , \33363 , \33364 , \33365 , \33366 , \33367 , \33368 , \33369 , \33370 ,
         \33371 , \33372 , \33373 , \33374 , \33375 , \33376 , \33377 , \33378 , \33379 , \33380 ,
         \33381 , \33382 , \33383 , \33384 , \33385 , \33386 , \33387 , \33388 , \33389 , \33390 ,
         \33391 , \33392 , \33393 , \33394 , \33395 , \33396 , \33397 , \33398 , \33399 , \33400 ,
         \33401 , \33402 , \33403 , \33404 , \33405 , \33406 , \33407 , \33408 , \33409 , \33410 ,
         \33411 , \33412 , \33413 , \33414 , \33415 , \33416 , \33417 , \33418 , \33419 , \33420 ,
         \33421 , \33422 , \33423 , \33424 , \33425 , \33426 , \33427 , \33428 , \33429 , \33430 ,
         \33431 , \33432 , \33433 , \33434 , \33435 , \33436 , \33437 , \33438 , \33439 , \33440 ,
         \33441 , \33442 , \33443 , \33444 , \33445 , \33446 , \33447 , \33448 , \33449 , \33450 ,
         \33451 , \33452 , \33453 , \33454 , \33455 , \33456 , \33457 , \33458 , \33459 , \33460 ,
         \33461 , \33462 , \33463 , \33464 , \33465 , \33466 , \33467 , \33468 , \33469 , \33470 ,
         \33471 , \33472 , \33473 , \33474 , \33475 , \33476 , \33477 , \33478 , \33479 , \33480 ,
         \33481 , \33482 , \33483 , \33484 , \33485 , \33486 , \33487 , \33488 , \33489 , \33490 ,
         \33491 , \33492 , \33493 , \33494 , \33495 , \33496 , \33497 , \33498 , \33499 , \33500 ,
         \33501 , \33502 , \33503 , \33504 , \33505 , \33506 , \33507 , \33508 , \33509 , \33510 ,
         \33511 , \33512 , \33513 , \33514 , \33515 , \33516 , \33517 , \33518 , \33519 , \33520 ,
         \33521 , \33522 , \33523 , \33524 , \33525 , \33526 , \33527 , \33528 , \33529 , \33530 ,
         \33531 , \33532 , \33533 , \33534 , \33535 , \33536 , \33537 , \33538 , \33539 , \33540 ,
         \33541 , \33542 , \33543 , \33544 , \33545 , \33546 , \33547 , \33548 , \33549 , \33550 ,
         \33551 , \33552 , \33553 , \33554 , \33555 , \33556 , \33557 , \33558 , \33559 , \33560 ,
         \33561 , \33562 , \33563 , \33564 , \33565 , \33566 , \33567 , \33568 , \33569 , \33570 ,
         \33571 , \33572 , \33573 , \33574 , \33575 , \33576 , \33577 , \33578 , \33579 , \33580 ,
         \33581 , \33582 , \33583 , \33584 , \33585 , \33586 , \33587 , \33588 , \33589 , \33590 ,
         \33591 , \33592 , \33593 , \33594 , \33595 , \33596 , \33597 , \33598 , \33599 , \33600 ,
         \33601 , \33602 , \33603 , \33604 , \33605 , \33606 , \33607 , \33608 , \33609 , \33610 ,
         \33611 , \33612 , \33613 , \33614 , \33615 , \33616 , \33617 , \33618 , \33619 , \33620 ,
         \33621 , \33622 , \33623 , \33624 , \33625 , \33626 , \33627 , \33628 , \33629 , \33630 ,
         \33631 , \33632 , \33633 , \33634 , \33635 , \33636 , \33637 , \33638 , \33639 , \33640 ,
         \33641 , \33642 , \33643 , \33644 , \33645 , \33646 , \33647 , \33648 , \33649 , \33650 ,
         \33651 , \33652 , \33653 , \33654 , \33655 , \33656 , \33657 , \33658 , \33659 , \33660 ,
         \33661 , \33662 , \33663 , \33664 , \33665 , \33666 , \33667 , \33668 , \33669 , \33670 ,
         \33671 , \33672 , \33673 , \33674 , \33675 , \33676 , \33677 , \33678 , \33679 , \33680 ,
         \33681 , \33682 , \33683 , \33684 , \33685 , \33686 , \33687 , \33688 , \33689 , \33690 ,
         \33691 , \33692 , \33693 , \33694 , \33695 , \33696 , \33697 , \33698 , \33699 , \33700 ,
         \33701 , \33702 , \33703 , \33704 , \33705 , \33706 , \33707 , \33708 , \33709 , \33710 ,
         \33711 , \33712 , \33713 , \33714 , \33715 , \33716 , \33717 , \33718 , \33719 , \33720 ,
         \33721 , \33722 , \33723 , \33724 , \33725 , \33726 , \33727 , \33728 , \33729 , \33730 ,
         \33731 , \33732 , \33733 , \33734 , \33735 , \33736 , \33737 , \33738 , \33739 , \33740 ,
         \33741 , \33742 , \33743 , \33744 , \33745 , \33746 , \33747 , \33748 , \33749 , \33750 ,
         \33751 , \33752 , \33753 , \33754 , \33755 , \33756 , \33757 , \33758 , \33759 , \33760 ,
         \33761 , \33762 , \33763 , \33764 , \33765 , \33766 , \33767 , \33768 , \33769 , \33770 ,
         \33771 , \33772 , \33773 , \33774 , \33775 , \33776 , \33777 , \33778 , \33779 , \33780 ,
         \33781 , \33782 , \33783 , \33784 , \33785 , \33786 , \33787 , \33788 , \33789 , \33790 ,
         \33791 , \33792 , \33793 , \33794 , \33795 , \33796 , \33797 , \33798 , \33799 , \33800 ,
         \33801 , \33802 , \33803 , \33804 , \33805 , \33806 , \33807 , \33808 , \33809 , \33810 ,
         \33811 , \33812 , \33813 , \33814 , \33815 , \33816 , \33817 , \33818 , \33819 , \33820 ,
         \33821 , \33822 , \33823 , \33824 , \33825 , \33826 , \33827 , \33828 , \33829 , \33830 ,
         \33831 , \33832 , \33833 , \33834 , \33835 , \33836 , \33837 , \33838 , \33839 , \33840 ,
         \33841 , \33842 , \33843 , \33844 , \33845 , \33846 , \33847 , \33848 , \33849 , \33850 ,
         \33851 , \33852 , \33853 , \33854 , \33855 , \33856 , \33857 , \33858 , \33859 , \33860 ,
         \33861 , \33862 , \33863 , \33864 , \33865 , \33866 , \33867 , \33868 , \33869 , \33870 ,
         \33871 , \33872 , \33873 , \33874 , \33875 , \33876 , \33877 , \33878 , \33879 , \33880 ,
         \33881 , \33882 , \33883 , \33884 , \33885 , \33886 , \33887 , \33888 , \33889 , \33890 ,
         \33891 , \33892 , \33893 , \33894 , \33895 , \33896 , \33897 , \33898 , \33899 , \33900 ,
         \33901 , \33902 , \33903 , \33904 , \33905 , \33906 , \33907 , \33908 , \33909 , \33910 ,
         \33911 , \33912 , \33913 , \33914 , \33915 , \33916 , \33917 , \33918 , \33919 , \33920 ,
         \33921 , \33922 , \33923 , \33924 , \33925 , \33926 , \33927 , \33928 , \33929 , \33930 ,
         \33931 , \33932 , \33933 , \33934 , \33935 , \33936 , \33937 , \33938 , \33939 , \33940 ,
         \33941 , \33942 , \33943 , \33944 , \33945 , \33946 , \33947 , \33948 , \33949 , \33950 ,
         \33951 , \33952 , \33953 , \33954 , \33955 , \33956 , \33957 , \33958 , \33959 , \33960 ,
         \33961 , \33962 , \33963 , \33964 , \33965 , \33966 , \33967 , \33968 , \33969 , \33970 ,
         \33971 , \33972 , \33973 , \33974 , \33975 , \33976 , \33977 , \33978 , \33979 , \33980 ,
         \33981 , \33982 , \33983 , \33984 , \33985 , \33986 , \33987 , \33988 , \33989 , \33990 ,
         \33991 , \33992 , \33993 , \33994 , \33995 , \33996 , \33997 , \33998 , \33999 , \34000 ,
         \34001 , \34002 , \34003 , \34004 , \34005 , \34006 , \34007 , \34008 , \34009 , \34010 ,
         \34011 , \34012 , \34013 , \34014 , \34015 , \34016 , \34017 , \34018 , \34019 , \34020 ,
         \34021 , \34022 , \34023 , \34024 , \34025 , \34026 , \34027 , \34028 , \34029 , \34030 ,
         \34031 , \34032 , \34033 , \34034 , \34035 , \34036 , \34037 , \34038 , \34039 , \34040 ,
         \34041 , \34042 , \34043 , \34044 , \34045 , \34046 , \34047 , \34048 , \34049 , \34050 ,
         \34051 , \34052 , \34053 , \34054 , \34055 , \34056 , \34057 , \34058 , \34059 , \34060 ,
         \34061 , \34062 , \34063 , \34064 , \34065 , \34066 , \34067 , \34068 , \34069 , \34070 ,
         \34071 , \34072 , \34073 , \34074 , \34075 , \34076 , \34077 , \34078 , \34079 , \34080 ,
         \34081 , \34082 , \34083 , \34084 , \34085 , \34086 , \34087 , \34088 , \34089 , \34090 ,
         \34091 , \34092 , \34093 , \34094 , \34095 , \34096 , \34097 , \34098 , \34099 , \34100 ,
         \34101 , \34102 , \34103 , \34104 , \34105 , \34106 , \34107 , \34108 , \34109 , \34110 ,
         \34111 , \34112 , \34113 , \34114 , \34115 , \34116 , \34117 , \34118 , \34119 , \34120 ,
         \34121 , \34122 , \34123 , \34124 , \34125 , \34126 , \34127 , \34128 , \34129 , \34130 ,
         \34131 , \34132 , \34133 , \34134 , \34135 , \34136 , \34137 , \34138 , \34139 , \34140 ,
         \34141 , \34142 , \34143 , \34144 , \34145 , \34146 , \34147 , \34148 , \34149 , \34150 ,
         \34151 , \34152 , \34153 , \34154 , \34155 , \34156 , \34157 , \34158 , \34159 , \34160 ,
         \34161 , \34162 , \34163 , \34164 , \34165 , \34166 , \34167 , \34168 , \34169 , \34170 ,
         \34171 , \34172 , \34173 , \34174 , \34175 , \34176 , \34177 , \34178 , \34179 , \34180 ,
         \34181 , \34182 , \34183 , \34184 , \34185 , \34186 , \34187 , \34188 , \34189 , \34190 ,
         \34191 , \34192 , \34193 , \34194 , \34195 , \34196 , \34197 , \34198 , \34199 , \34200 ,
         \34201 , \34202 , \34203 , \34204 , \34205 , \34206 , \34207 , \34208 , \34209 , \34210 ,
         \34211 , \34212 , \34213 , \34214 , \34215 , \34216 , \34217 , \34218 , \34219 , \34220 ,
         \34221 , \34222 , \34223 , \34224 , \34225 , \34226 , \34227 , \34228 , \34229 , \34230 ,
         \34231 , \34232 , \34233 , \34234 , \34235 , \34236 , \34237 , \34238 , \34239 , \34240 ,
         \34241 , \34242 , \34243 , \34244 , \34245 , \34246 , \34247 , \34248 , \34249 , \34250 ,
         \34251 , \34252 , \34253 , \34254 , \34255 , \34256 , \34257 , \34258 , \34259 , \34260 ,
         \34261 , \34262 , \34263 , \34264 , \34265 , \34266 , \34267 , \34268 , \34269 , \34270 ,
         \34271 , \34272 , \34273 , \34274 , \34275 , \34276 , \34277 , \34278 , \34279 , \34280 ,
         \34281 , \34282 , \34283 , \34284 , \34285 , \34286 , \34287 , \34288 , \34289 , \34290 ,
         \34291 , \34292 , \34293 , \34294 , \34295 , \34296 , \34297 , \34298 , \34299 , \34300 ,
         \34301 , \34302 , \34303 , \34304 , \34305 , \34306 , \34307 , \34308 , \34309 , \34310 ,
         \34311 , \34312 , \34313 , \34314 , \34315 , \34316 , \34317 , \34318 , \34319 , \34320 ,
         \34321 , \34322 , \34323 , \34324 , \34325 , \34326 , \34327 , \34328 , \34329 , \34330 ,
         \34331 , \34332 , \34333 , \34334 , \34335 , \34336 , \34337 , \34338 , \34339 , \34340 ,
         \34341 , \34342 , \34343 , \34344 , \34345 , \34346 , \34347 , \34348 , \34349 , \34350 ,
         \34351 , \34352 , \34353 , \34354 , \34355 , \34356 , \34357 , \34358 , \34359 , \34360 ,
         \34361 , \34362 , \34363 , \34364 , \34365 , \34366 , \34367 , \34368 , \34369 , \34370 ,
         \34371 , \34372 , \34373 , \34374 , \34375 , \34376 , \34377 , \34378 , \34379 , \34380 ,
         \34381 , \34382 , \34383 , \34384 , \34385 , \34386 , \34387 , \34388 , \34389 , \34390 ,
         \34391 , \34392 , \34393 , \34394 , \34395 , \34396 , \34397 , \34398 , \34399 , \34400 ,
         \34401 , \34402 , \34403 , \34404 , \34405 , \34406 , \34407 , \34408 , \34409 , \34410 ,
         \34411 , \34412 , \34413 , \34414 , \34415 , \34416 , \34417 , \34418 , \34419 , \34420 ,
         \34421 , \34422 , \34423 , \34424 , \34425 , \34426 , \34427 , \34428 , \34429 , \34430 ,
         \34431 , \34432 , \34433 , \34434 , \34435 , \34436 , \34437 , \34438 , \34439 , \34440 ,
         \34441 , \34442 , \34443 , \34444 , \34445 , \34446 , \34447 , \34448 , \34449 , \34450 ,
         \34451 , \34452 , \34453 , \34454 , \34455 , \34456 , \34457 , \34458 , \34459 , \34460 ,
         \34461 , \34462 , \34463 , \34464 , \34465 , \34466 , \34467 , \34468 , \34469 , \34470 ,
         \34471 , \34472 , \34473 , \34474 , \34475 , \34476 , \34477 , \34478 , \34479 , \34480 ,
         \34481 , \34482 , \34483 , \34484 , \34485 , \34486 , \34487 , \34488 , \34489 , \34490 ,
         \34491 , \34492 , \34493 , \34494 , \34495 , \34496 , \34497 , \34498 , \34499 , \34500 ,
         \34501 , \34502 , \34503 , \34504 , \34505 , \34506 , \34507 , \34508 , \34509 , \34510 ,
         \34511 , \34512 , \34513 , \34514 , \34515 , \34516 , \34517 , \34518 , \34519 , \34520 ,
         \34521 , \34522 , \34523 , \34524 , \34525 , \34526 , \34527 , \34528 , \34529 , \34530 ,
         \34531 , \34532 , \34533 , \34534 , \34535 , \34536 , \34537 , \34538 , \34539 , \34540 ,
         \34541 , \34542 , \34543 , \34544 , \34545 , \34546 , \34547 , \34548 , \34549 , \34550 ,
         \34551 , \34552 , \34553 , \34554 , \34555 , \34556 , \34557 , \34558 , \34559 , \34560 ,
         \34561 , \34562 , \34563 , \34564 , \34565 , \34566 , \34567 , \34568 , \34569 , \34570 ,
         \34571 , \34572 , \34573 , \34574 , \34575 , \34576 , \34577 , \34578 , \34579 , \34580 ,
         \34581 , \34582 , \34583 , \34584 , \34585 , \34586 , \34587 , \34588 , \34589 , \34590 ,
         \34591 , \34592 , \34593 , \34594 , \34595 , \34596 , \34597 , \34598 , \34599 , \34600 ,
         \34601 , \34602 , \34603 , \34604 , \34605 , \34606 , \34607 , \34608 , \34609 , \34610 ,
         \34611 , \34612 , \34613 , \34614 , \34615 , \34616 , \34617 , \34618 , \34619 , \34620 ,
         \34621 , \34622 , \34623 , \34624 , \34625 , \34626 , \34627 , \34628 , \34629 , \34630 ,
         \34631 , \34632 , \34633 , \34634 , \34635 , \34636 , \34637 , \34638 , \34639 , \34640 ,
         \34641 , \34642 , \34643 , \34644 , \34645 , \34646 , \34647 , \34648 , \34649 , \34650 ,
         \34651 , \34652 , \34653 , \34654 , \34655 , \34656 , \34657 , \34658 , \34659 , \34660 ,
         \34661 , \34662 , \34663 , \34664 , \34665 , \34666 , \34667 , \34668 , \34669 , \34670 ,
         \34671 , \34672 , \34673 , \34674 , \34675 , \34676 , \34677 , \34678 , \34679 , \34680 ,
         \34681 , \34682 , \34683 , \34684 , \34685 , \34686 , \34687 , \34688 , \34689 , \34690 ,
         \34691 , \34692 , \34693 , \34694 , \34695 , \34696 , \34697 , \34698 , \34699 , \34700 ,
         \34701 , \34702 , \34703 , \34704 , \34705 , \34706 , \34707 , \34708 , \34709 , \34710 ,
         \34711 , \34712 , \34713 , \34714 , \34715 , \34716 , \34717 , \34718 , \34719 , \34720 ,
         \34721 , \34722 , \34723 , \34724 , \34725 , \34726 , \34727 , \34728 , \34729 , \34730 ,
         \34731 , \34732 , \34733 , \34734 , \34735 , \34736 , \34737 , \34738 , \34739 , \34740 ,
         \34741 , \34742 , \34743 , \34744 , \34745 , \34746 , \34747 , \34748 , \34749 , \34750 ,
         \34751 , \34752 , \34753 , \34754 , \34755 , \34756 , \34757 , \34758 , \34759 , \34760 ,
         \34761 , \34762 , \34763 , \34764 , \34765 , \34766 , \34767 , \34768 , \34769 , \34770 ,
         \34771 , \34772 , \34773 , \34774 , \34775 , \34776 , \34777 , \34778 , \34779 , \34780 ,
         \34781 , \34782 , \34783 , \34784 , \34785 , \34786 , \34787 , \34788 , \34789 , \34790 ,
         \34791 , \34792 , \34793 , \34794 , \34795 , \34796 , \34797 , \34798 , \34799 , \34800 ,
         \34801 , \34802 , \34803 , \34804 , \34805 , \34806 , \34807 , \34808 , \34809 , \34810 ,
         \34811 , \34812 , \34813 , \34814 , \34815 , \34816 , \34817 , \34818 , \34819 , \34820 ,
         \34821 , \34822 , \34823 , \34824 , \34825 , \34826 , \34827 , \34828 , \34829 , \34830 ,
         \34831 , \34832 , \34833 , \34834 , \34835 , \34836 , \34837 , \34838 , \34839 , \34840 ,
         \34841 , \34842 , \34843 , \34844 , \34845 , \34846 , \34847 , \34848 , \34849 , \34850 ,
         \34851 , \34852 , \34853 , \34854 , \34855 , \34856 , \34857 , \34858 , \34859 , \34860 ,
         \34861 , \34862 , \34863 , \34864 , \34865 , \34866 , \34867 , \34868 , \34869 , \34870 ,
         \34871 , \34872 , \34873 , \34874 , \34875 , \34876 , \34877 , \34878 , \34879 , \34880 ,
         \34881 , \34882 , \34883 , \34884 , \34885 , \34886 , \34887 , \34888 , \34889 , \34890 ,
         \34891 , \34892 , \34893 , \34894 , \34895 , \34896 , \34897 , \34898 , \34899 , \34900 ,
         \34901 , \34902 , \34903 , \34904 , \34905 , \34906 , \34907 , \34908 , \34909 , \34910 ,
         \34911 , \34912 , \34913 , \34914 , \34915 , \34916 , \34917 , \34918 , \34919 , \34920 ,
         \34921 , \34922 , \34923 , \34924 , \34925 , \34926 , \34927 , \34928 , \34929 , \34930 ,
         \34931 , \34932 , \34933 , \34934 , \34935 , \34936 , \34937 , \34938 , \34939 , \34940 ,
         \34941 , \34942 , \34943 , \34944 , \34945 , \34946 , \34947 , \34948 , \34949 , \34950 ,
         \34951 , \34952 , \34953 , \34954 , \34955 , \34956 , \34957 , \34958 , \34959 , \34960 ,
         \34961 , \34962 , \34963 , \34964 , \34965 , \34966 , \34967 , \34968 , \34969 , \34970 ,
         \34971 , \34972 , \34973 , \34974 , \34975 , \34976 , \34977 , \34978 , \34979 , \34980 ,
         \34981 , \34982 , \34983 , \34984 , \34985 , \34986 , \34987 , \34988 , \34989 , \34990 ,
         \34991 , \34992 , \34993 , \34994 , \34995 , \34996 , \34997 , \34998 , \34999 , \35000 ,
         \35001 , \35002 , \35003 , \35004 , \35005 , \35006 , \35007 , \35008 , \35009 , \35010 ,
         \35011 , \35012 , \35013 , \35014 , \35015 , \35016 , \35017 , \35018 , \35019 , \35020 ,
         \35021 , \35022 , \35023 , \35024 , \35025 , \35026 , \35027 , \35028 , \35029 , \35030 ,
         \35031 , \35032 , \35033 , \35034 , \35035 , \35036 , \35037 , \35038 , \35039 , \35040 ,
         \35041 , \35042 , \35043 , \35044 , \35045 , \35046 , \35047 , \35048 , \35049 , \35050 ,
         \35051 , \35052 , \35053 , \35054 , \35055 , \35056 , \35057 , \35058 , \35059 , \35060 ,
         \35061 , \35062 , \35063 , \35064 , \35065 , \35066 , \35067 , \35068 , \35069 , \35070 ,
         \35071 , \35072 , \35073 , \35074 , \35075 , \35076 , \35077 , \35078 , \35079 , \35080 ,
         \35081 , \35082 , \35083 , \35084 , \35085 , \35086 , \35087 , \35088 , \35089 , \35090 ,
         \35091 , \35092 , \35093 , \35094 , \35095 , \35096 , \35097 , \35098 , \35099 , \35100 ,
         \35101 , \35102 , \35103 , \35104 , \35105 , \35106 , \35107 , \35108 , \35109 , \35110 ,
         \35111 , \35112 , \35113 , \35114 , \35115 , \35116 , \35117 , \35118 , \35119 , \35120 ,
         \35121 , \35122 , \35123 , \35124 , \35125 , \35126 , \35127 , \35128 , \35129 , \35130 ,
         \35131 , \35132 , \35133 , \35134 , \35135 , \35136 , \35137 , \35138 , \35139 , \35140 ,
         \35141 , \35142 , \35143 , \35144 , \35145 , \35146 , \35147 , \35148 , \35149 , \35150 ,
         \35151 , \35152 , \35153 , \35154 , \35155 , \35156 , \35157 , \35158 , \35159 , \35160 ,
         \35161 , \35162 , \35163 , \35164 , \35165 , \35166 , \35167 , \35168 , \35169 , \35170 ,
         \35171 , \35172 , \35173 , \35174 , \35175 , \35176 , \35177 , \35178 , \35179 , \35180 ,
         \35181 , \35182 , \35183 , \35184 , \35185 , \35186 , \35187 , \35188 , \35189 , \35190 ,
         \35191 , \35192 , \35193 , \35194 , \35195 , \35196 , \35197 , \35198 , \35199 , \35200 ,
         \35201 , \35202 , \35203 , \35204 , \35205 , \35206 , \35207 , \35208 , \35209 , \35210 ,
         \35211 , \35212 , \35213 , \35214 , \35215 , \35216 , \35217 , \35218 , \35219 , \35220 ,
         \35221 , \35222 , \35223 , \35224 , \35225 , \35226 , \35227 , \35228 , \35229 , \35230 ,
         \35231 , \35232 , \35233 , \35234 , \35235 , \35236 , \35237 , \35238 , \35239 , \35240 ,
         \35241 , \35242 , \35243 , \35244 , \35245 , \35246 , \35247 , \35248 , \35249 , \35250 ,
         \35251 , \35252 , \35253 , \35254 , \35255 , \35256 , \35257 , \35258 , \35259 , \35260 ,
         \35261 , \35262 , \35263 , \35264 , \35265 , \35266 , \35267 , \35268 , \35269 , \35270 ,
         \35271 , \35272 , \35273 , \35274 , \35275 , \35276 , \35277 , \35278 , \35279 , \35280 ,
         \35281 , \35282 , \35283 , \35284 , \35285 , \35286 , \35287 , \35288 , \35289 , \35290 ,
         \35291 , \35292 , \35293 , \35294 , \35295 , \35296 , \35297 , \35298 , \35299 , \35300 ,
         \35301 , \35302 , \35303 , \35304 , \35305 , \35306 , \35307 , \35308 , \35309 , \35310 ,
         \35311 , \35312 , \35313 , \35314 , \35315 , \35316 , \35317 , \35318 , \35319 , \35320 ,
         \35321 , \35322 , \35323 , \35324 , \35325 , \35326 , \35327 , \35328 , \35329 , \35330 ,
         \35331 , \35332 , \35333 , \35334 , \35335 , \35336 , \35337 , \35338 , \35339 , \35340 ,
         \35341 , \35342 , \35343 , \35344 , \35345 , \35346 , \35347 , \35348 , \35349 , \35350 ,
         \35351 , \35352 , \35353 , \35354 , \35355 , \35356 , \35357 , \35358 , \35359 , \35360 ,
         \35361 , \35362 , \35363 , \35364 , \35365 , \35366 , \35367 , \35368 , \35369 , \35370 ,
         \35371 , \35372 , \35373 , \35374 , \35375 , \35376 , \35377 , \35378 , \35379 , \35380 ,
         \35381 , \35382 , \35383 , \35384 , \35385 , \35386 , \35387 , \35388 , \35389 , \35390 ,
         \35391 , \35392 , \35393 , \35394 , \35395 , \35396 , \35397 , \35398 , \35399 , \35400 ,
         \35401 , \35402 , \35403 , \35404 , \35405 , \35406 , \35407 , \35408 , \35409 , \35410 ,
         \35411 , \35412 , \35413 , \35414 , \35415 , \35416 , \35417 , \35418 , \35419 , \35420 ,
         \35421 , \35422 , \35423 , \35424 , \35425 , \35426 , \35427 , \35428 , \35429 , \35430 ,
         \35431 , \35432 , \35433 , \35434 , \35435 , \35436 , \35437 , \35438 , \35439 , \35440 ,
         \35441 , \35442 , \35443 , \35444 , \35445 , \35446 , \35447 , \35448 , \35449 , \35450 ,
         \35451 , \35452 , \35453 , \35454 , \35455 , \35456 , \35457 , \35458 , \35459 , \35460 ,
         \35461 , \35462 , \35463 , \35464 , \35465 , \35466 , \35467 , \35468 , \35469 , \35470 ,
         \35471 , \35472 , \35473 , \35474 , \35475 , \35476 , \35477 , \35478 , \35479 , \35480 ,
         \35481 , \35482 , \35483 , \35484 , \35485 , \35486 , \35487 , \35488 , \35489 , \35490 ,
         \35491 , \35492 , \35493 , \35494 , \35495 , \35496 , \35497 , \35498 , \35499 , \35500 ,
         \35501 , \35502 , \35503 , \35504 , \35505 , \35506 , \35507 , \35508 , \35509 , \35510 ,
         \35511 , \35512 , \35513 , \35514 , \35515 , \35516 , \35517 , \35518 , \35519 , \35520 ,
         \35521 , \35522 , \35523 , \35524 , \35525 , \35526 , \35527 , \35528 , \35529 , \35530 ,
         \35531 , \35532 , \35533 , \35534 , \35535 , \35536 , \35537 , \35538 , \35539 , \35540 ,
         \35541 , \35542 , \35543 , \35544 , \35545 , \35546 , \35547 , \35548 , \35549 , \35550 ,
         \35551 , \35552 , \35553 , \35554 , \35555 , \35556 , \35557 , \35558 , \35559 , \35560 ,
         \35561 , \35562 , \35563 , \35564 , \35565 , \35566 , \35567 , \35568 , \35569 , \35570 ,
         \35571 , \35572 , \35573 , \35574 , \35575 , \35576 , \35577 , \35578 , \35579 , \35580 ,
         \35581 , \35582 , \35583 , \35584 , \35585 , \35586 , \35587 , \35588 , \35589 , \35590 ,
         \35591 , \35592 , \35593 , \35594 , \35595 , \35596 , \35597 , \35598 , \35599 , \35600 ,
         \35601 , \35602 , \35603 , \35604 , \35605 , \35606 , \35607 , \35608 , \35609 , \35610 ,
         \35611 , \35612 , \35613 , \35614 , \35615 , \35616 , \35617 , \35618 , \35619 , \35620 ,
         \35621 , \35622 , \35623 , \35624 , \35625 , \35626 , \35627 , \35628 , \35629 , \35630 ,
         \35631 , \35632 , \35633 , \35634 , \35635 , \35636 , \35637 , \35638 , \35639 , \35640 ,
         \35641 , \35642 , \35643 , \35644 , \35645 , \35646 , \35647 , \35648 , \35649 , \35650 ,
         \35651 , \35652 , \35653 , \35654 , \35655 , \35656 , \35657 , \35658 , \35659 , \35660 ,
         \35661 , \35662 , \35663 , \35664 , \35665 , \35666 , \35667 , \35668 , \35669 , \35670 ,
         \35671 , \35672 , \35673 , \35674 , \35675 , \35676 , \35677 , \35678 , \35679 , \35680 ,
         \35681 , \35682 , \35683 , \35684 , \35685 , \35686 , \35687 , \35688 , \35689 , \35690 ,
         \35691 , \35692 , \35693 , \35694 , \35695 , \35696 , \35697 , \35698 , \35699 , \35700 ,
         \35701 , \35702 , \35703 , \35704 , \35705 , \35706 , \35707 , \35708 , \35709 , \35710 ,
         \35711 , \35712 , \35713 , \35714 , \35715 , \35716 , \35717 , \35718 , \35719 , \35720 ,
         \35721 , \35722 , \35723 , \35724 , \35725 , \35726 , \35727 , \35728 , \35729 , \35730 ,
         \35731 , \35732 , \35733 , \35734 , \35735 , \35736 , \35737 , \35738 , \35739 , \35740 ,
         \35741 , \35742 , \35743 , \35744 , \35745 , \35746 , \35747 , \35748 , \35749 , \35750 ,
         \35751 , \35752 , \35753 , \35754 , \35755 , \35756 , \35757 , \35758 , \35759 , \35760 ,
         \35761 , \35762 , \35763 , \35764 , \35765 , \35766 , \35767 , \35768 , \35769 , \35770 ,
         \35771 , \35772 , \35773 , \35774 , \35775 , \35776 , \35777 , \35778 , \35779 , \35780 ,
         \35781 , \35782 , \35783 , \35784 , \35785 , \35786 , \35787 , \35788 , \35789 , \35790 ,
         \35791 , \35792 , \35793 , \35794 , \35795 , \35796 , \35797 , \35798 , \35799 , \35800 ,
         \35801 , \35802 , \35803 , \35804 , \35805 , \35806 , \35807 , \35808 , \35809 , \35810 ,
         \35811 , \35812 , \35813 , \35814 , \35815 , \35816 , \35817 , \35818 , \35819 , \35820 ,
         \35821 , \35822 , \35823 , \35824 , \35825 , \35826 , \35827 , \35828 , \35829 , \35830 ,
         \35831 , \35832 , \35833 , \35834 , \35835 , \35836 , \35837 , \35838 , \35839 , \35840 ,
         \35841 , \35842 , \35843 , \35844 , \35845 , \35846 , \35847 , \35848 , \35849 , \35850 ,
         \35851 , \35852 , \35853 , \35854 , \35855 , \35856 , \35857 , \35858 , \35859 , \35860 ,
         \35861 , \35862 , \35863 , \35864 , \35865 , \35866 , \35867 , \35868 , \35869 , \35870 ,
         \35871 , \35872 , \35873 , \35874 , \35875 , \35876 , \35877 , \35878 , \35879 , \35880 ,
         \35881 , \35882 , \35883 , \35884 , \35885 , \35886 , \35887 , \35888 , \35889 , \35890 ,
         \35891 , \35892 , \35893 , \35894 , \35895 , \35896 , \35897 , \35898 , \35899 , \35900 ,
         \35901 , \35902 , \35903 , \35904 , \35905 , \35906 , \35907 , \35908 , \35909 , \35910 ,
         \35911 , \35912 , \35913 , \35914 , \35915 , \35916 , \35917 , \35918 , \35919 , \35920 ,
         \35921 , \35922 , \35923 , \35924 , \35925 , \35926 , \35927 , \35928 , \35929 , \35930 ,
         \35931 , \35932 , \35933 , \35934 , \35935 , \35936 , \35937 , \35938 , \35939 , \35940 ,
         \35941 , \35942 , \35943 , \35944 , \35945 , \35946 , \35947 , \35948 , \35949 , \35950 ,
         \35951 , \35952 , \35953 , \35954 , \35955 , \35956 , \35957 , \35958 , \35959 , \35960 ,
         \35961 , \35962 , \35963 , \35964 , \35965 , \35966 , \35967 , \35968 , \35969 , \35970 ,
         \35971 , \35972 , \35973 , \35974 , \35975 , \35976 , \35977 , \35978 , \35979 , \35980 ,
         \35981 , \35982 , \35983 , \35984 , \35985 , \35986 , \35987 , \35988 , \35989 , \35990 ,
         \35991 , \35992 , \35993 , \35994 , \35995 , \35996 , \35997 , \35998 , \35999 , \36000 ,
         \36001 , \36002 , \36003 , \36004 , \36005 , \36006 , \36007 , \36008 , \36009 , \36010 ,
         \36011 , \36012 , \36013 , \36014 , \36015 , \36016 , \36017 , \36018 , \36019 , \36020 ,
         \36021 , \36022 , \36023 , \36024 , \36025 , \36026 , \36027 , \36028 , \36029 , \36030 ,
         \36031 , \36032 , \36033 , \36034 , \36035 , \36036 , \36037 , \36038 , \36039 , \36040 ,
         \36041 , \36042 , \36043 , \36044 , \36045 , \36046 , \36047 , \36048 , \36049 , \36050 ,
         \36051 , \36052 , \36053 , \36054 , \36055 , \36056 , \36057 , \36058 , \36059 , \36060 ,
         \36061 , \36062 , \36063 , \36064 , \36065 , \36066 , \36067 , \36068 , \36069 , \36070 ,
         \36071 , \36072 , \36073 , \36074 , \36075 , \36076 , \36077 , \36078 , \36079 , \36080 ,
         \36081 , \36082 , \36083 , \36084 , \36085 , \36086 , \36087 , \36088 , \36089 , \36090 ,
         \36091 , \36092 , \36093 , \36094 , \36095 , \36096 , \36097 , \36098 , \36099 , \36100 ,
         \36101 , \36102 , \36103 , \36104 , \36105 , \36106 , \36107 , \36108 , \36109 , \36110 ,
         \36111 , \36112 , \36113 , \36114 , \36115 , \36116 , \36117 , \36118 , \36119 , \36120 ,
         \36121 , \36122 , \36123 , \36124 , \36125 , \36126 , \36127 , \36128 , \36129 , \36130 ,
         \36131 , \36132 , \36133 , \36134 , \36135 , \36136 , \36137 , \36138 , \36139 , \36140 ,
         \36141 , \36142 , \36143 , \36144 , \36145 , \36146 , \36147 , \36148 , \36149 , \36150 ,
         \36151 , \36152 , \36153 , \36154 , \36155 , \36156 , \36157 , \36158 , \36159 , \36160 ,
         \36161 , \36162 , \36163 , \36164 , \36165 , \36166 , \36167 , \36168 , \36169 , \36170 ,
         \36171 , \36172 , \36173 , \36174 , \36175 , \36176 , \36177 , \36178 , \36179 , \36180 ,
         \36181 , \36182 , \36183 , \36184 , \36185 , \36186 , \36187 , \36188 , \36189 , \36190 ,
         \36191 , \36192 , \36193 , \36194 , \36195 , \36196 , \36197 , \36198 , \36199 , \36200 ,
         \36201 , \36202 , \36203 , \36204 , \36205 , \36206 , \36207 , \36208 , \36209 , \36210 ,
         \36211 , \36212 , \36213 , \36214 , \36215 , \36216 , \36217 , \36218 , \36219 , \36220 ,
         \36221 , \36222 , \36223 , \36224 , \36225 , \36226 , \36227 , \36228 , \36229 , \36230 ,
         \36231 , \36232 , \36233 , \36234 , \36235 , \36236 , \36237 , \36238 , \36239 , \36240 ,
         \36241 , \36242 , \36243 , \36244 , \36245 , \36246 , \36247 , \36248 , \36249 , \36250 ,
         \36251 , \36252 , \36253 , \36254 , \36255 , \36256 , \36257 , \36258 , \36259 , \36260 ,
         \36261 , \36262 , \36263 , \36264 , \36265 , \36266 , \36267 , \36268 , \36269 , \36270 ,
         \36271 , \36272 , \36273 , \36274 , \36275 , \36276 , \36277 , \36278 , \36279 , \36280 ,
         \36281 , \36282 , \36283 , \36284 , \36285 , \36286 , \36287 , \36288 , \36289 , \36290 ,
         \36291 , \36292 , \36293 , \36294 , \36295 , \36296 , \36297 , \36298 , \36299 , \36300 ,
         \36301 , \36302 , \36303 , \36304 , \36305 , \36306 , \36307 , \36308 , \36309 , \36310 ,
         \36311 , \36312 , \36313 , \36314 , \36315 , \36316 , \36317 , \36318 , \36319 , \36320 ,
         \36321 , \36322 , \36323 , \36324 , \36325 , \36326 , \36327 , \36328 , \36329 , \36330 ,
         \36331 , \36332 , \36333 , \36334 , \36335 , \36336 , \36337 , \36338 , \36339 , \36340 ,
         \36341 , \36342 , \36343 , \36344 , \36345 , \36346 , \36347 , \36348 , \36349 , \36350 ,
         \36351 , \36352 , \36353 , \36354 , \36355 , \36356 , \36357 , \36358 , \36359 , \36360 ,
         \36361 , \36362 , \36363 , \36364 , \36365 , \36366 , \36367 , \36368 , \36369 , \36370 ,
         \36371 , \36372 , \36373 , \36374 , \36375 , \36376 , \36377 , \36378 , \36379 , \36380 ,
         \36381 , \36382 , \36383 , \36384 , \36385 , \36386 , \36387 , \36388 , \36389 , \36390 ,
         \36391 , \36392 , \36393 , \36394 , \36395 , \36396 , \36397 , \36398 , \36399 , \36400 ,
         \36401 , \36402 , \36403 , \36404 , \36405 , \36406 , \36407 , \36408 , \36409 , \36410 ,
         \36411 , \36412 , \36413 , \36414 , \36415 , \36416 , \36417 , \36418 , \36419 , \36420 ,
         \36421 , \36422 , \36423 , \36424 , \36425 , \36426 , \36427 , \36428 , \36429 , \36430 ,
         \36431 , \36432 , \36433 , \36434 , \36435 , \36436 , \36437 , \36438 , \36439 , \36440 ,
         \36441 , \36442 , \36443 , \36444 , \36445 , \36446 , \36447 , \36448 , \36449 , \36450 ,
         \36451 , \36452 , \36453 , \36454 , \36455 , \36456 , \36457 , \36458 , \36459 , \36460 ,
         \36461 , \36462 , \36463 , \36464 , \36465 , \36466 , \36467 , \36468 , \36469 , \36470 ,
         \36471 , \36472 , \36473 , \36474 , \36475 , \36476 , \36477 , \36478 , \36479 , \36480 ,
         \36481 , \36482 , \36483 , \36484 , \36485 , \36486 , \36487 , \36488 , \36489 , \36490 ,
         \36491 , \36492 , \36493 , \36494 , \36495 , \36496 , \36497 , \36498 , \36499 , \36500 ,
         \36501 , \36502 , \36503 , \36504 , \36505 , \36506 , \36507 , \36508 , \36509 , \36510 ,
         \36511 , \36512 , \36513 , \36514 , \36515 , \36516 , \36517 , \36518 , \36519 , \36520 ,
         \36521 , \36522 , \36523 , \36524 , \36525 , \36526 , \36527 , \36528 , \36529 , \36530 ,
         \36531 , \36532 , \36533 , \36534 , \36535 , \36536 , \36537 , \36538 , \36539 , \36540 ,
         \36541 , \36542 , \36543 , \36544 , \36545 , \36546 , \36547 , \36548 , \36549 , \36550 ,
         \36551 , \36552 , \36553 , \36554 , \36555 , \36556 , \36557 , \36558 , \36559 , \36560 ,
         \36561 , \36562 , \36563 , \36564 , \36565 , \36566 , \36567 , \36568 , \36569 , \36570 ,
         \36571 , \36572 , \36573 , \36574 , \36575 , \36576 , \36577 , \36578 , \36579 , \36580 ,
         \36581 , \36582 , \36583 , \36584 , \36585 , \36586 , \36587 , \36588 , \36589 , \36590 ,
         \36591 , \36592 , \36593 , \36594 , \36595 , \36596 , \36597 , \36598 , \36599 , \36600 ,
         \36601 , \36602 , \36603 , \36604 , \36605 , \36606 , \36607 , \36608 , \36609 , \36610 ,
         \36611 , \36612 , \36613 , \36614 , \36615 , \36616 , \36617 , \36618 , \36619 , \36620 ,
         \36621 , \36622 , \36623 , \36624 , \36625 , \36626 , \36627 , \36628 , \36629 , \36630 ,
         \36631 , \36632 , \36633 , \36634 , \36635 , \36636 , \36637 , \36638 , \36639 , \36640 ,
         \36641 , \36642 , \36643 , \36644 , \36645 , \36646 , \36647 , \36648 , \36649 , \36650 ,
         \36651 , \36652 , \36653 , \36654 , \36655 , \36656 , \36657 , \36658 , \36659 , \36660 ,
         \36661 , \36662 , \36663 , \36664 , \36665 , \36666 , \36667 , \36668 , \36669 , \36670 ,
         \36671 , \36672 , \36673 , \36674 , \36675 , \36676 , \36677 , \36678 , \36679 , \36680 ,
         \36681 , \36682 , \36683 , \36684 , \36685 , \36686 , \36687 , \36688 , \36689 , \36690 ,
         \36691 , \36692 , \36693 , \36694 , \36695 , \36696 , \36697 , \36698 , \36699 , \36700 ,
         \36701 , \36702 , \36703 , \36704 , \36705 , \36706 , \36707 , \36708 , \36709 , \36710 ,
         \36711 , \36712 , \36713 , \36714 , \36715 , \36716 , \36717 , \36718 , \36719 , \36720 ,
         \36721 , \36722 , \36723 , \36724 , \36725 , \36726 , \36727 , \36728 , \36729 , \36730 ,
         \36731 , \36732 , \36733 , \36734 , \36735 , \36736 , \36737 , \36738 , \36739 , \36740 ,
         \36741 , \36742 , \36743 , \36744 , \36745 , \36746 , \36747 , \36748 , \36749 , \36750 ,
         \36751 , \36752 , \36753 , \36754 , \36755 , \36756 , \36757 , \36758 , \36759 , \36760 ,
         \36761 , \36762 , \36763 , \36764 , \36765 , \36766 , \36767 , \36768 , \36769 , \36770 ,
         \36771 , \36772 , \36773 , \36774 , \36775 , \36776 , \36777 , \36778 , \36779 , \36780 ,
         \36781 , \36782 , \36783 , \36784 , \36785 , \36786 , \36787 , \36788 , \36789 , \36790 ,
         \36791 , \36792 , \36793 , \36794 , \36795 , \36796 , \36797 , \36798 , \36799 , \36800 ,
         \36801 , \36802 , \36803 , \36804 , \36805 , \36806 , \36807 , \36808 , \36809 , \36810 ,
         \36811 , \36812 , \36813 , \36814 , \36815 , \36816 , \36817 , \36818 , \36819 , \36820 ,
         \36821 , \36822 , \36823 , \36824 , \36825 , \36826 , \36827 , \36828 , \36829 , \36830 ,
         \36831 , \36832 , \36833 , \36834 , \36835 , \36836 , \36837 , \36838 , \36839 , \36840 ,
         \36841 , \36842 , \36843 , \36844 , \36845 , \36846 , \36847 , \36848 , \36849 , \36850 ,
         \36851 , \36852 , \36853 , \36854 , \36855 , \36856 , \36857 , \36858 , \36859 , \36860 ,
         \36861 , \36862 , \36863 , \36864 , \36865 , \36866 , \36867 , \36868 , \36869 , \36870 ,
         \36871 , \36872 , \36873 , \36874 , \36875 , \36876 , \36877 , \36878 , \36879 , \36880 ,
         \36881 , \36882 , \36883 , \36884 , \36885 , \36886 , \36887 , \36888 , \36889 , \36890 ,
         \36891 , \36892 , \36893 , \36894 , \36895 , \36896 , \36897 , \36898 , \36899 , \36900 ,
         \36901 , \36902 , \36903 , \36904 , \36905 , \36906 , \36907 , \36908 , \36909 , \36910 ,
         \36911 , \36912 , \36913 , \36914 , \36915 , \36916 , \36917 , \36918 , \36919 , \36920 ,
         \36921 , \36922 , \36923 , \36924 , \36925 , \36926 , \36927 , \36928 , \36929 , \36930 ,
         \36931 , \36932 , \36933 , \36934 , \36935 , \36936 , \36937 , \36938 , \36939 , \36940 ,
         \36941 , \36942 , \36943 , \36944 , \36945 , \36946 , \36947 , \36948 , \36949 , \36950 ,
         \36951 , \36952 , \36953 , \36954 , \36955 , \36956 , \36957 , \36958 , \36959 , \36960 ,
         \36961 , \36962 , \36963 , \36964 , \36965 , \36966 , \36967 , \36968 , \36969 , \36970 ,
         \36971 , \36972 , \36973 , \36974 , \36975 , \36976 , \36977 , \36978 , \36979 , \36980 ,
         \36981 , \36982 , \36983 , \36984 , \36985 , \36986 , \36987 , \36988 , \36989 , \36990 ,
         \36991 , \36992 , \36993 , \36994 , \36995 , \36996 , \36997 , \36998 , \36999 , \37000 ,
         \37001 , \37002 , \37003 , \37004 , \37005 , \37006 , \37007 , \37008 , \37009 , \37010 ,
         \37011 , \37012 , \37013 , \37014 , \37015 , \37016 , \37017 , \37018 , \37019 , \37020 ,
         \37021 , \37022 , \37023 , \37024 , \37025 , \37026 , \37027 , \37028 , \37029 , \37030 ,
         \37031 , \37032 , \37033 , \37034 , \37035 , \37036 , \37037 , \37038 , \37039 , \37040 ,
         \37041 , \37042 , \37043 , \37044 , \37045 , \37046 , \37047 , \37048 , \37049 , \37050 ,
         \37051 , \37052 , \37053 , \37054 , \37055 , \37056 , \37057 , \37058 , \37059 , \37060 ,
         \37061 , \37062 , \37063 , \37064 , \37065 , \37066 , \37067 , \37068 , \37069 , \37070 ,
         \37071 , \37072 , \37073 , \37074 , \37075 , \37076 , \37077 , \37078 , \37079 , \37080 ,
         \37081 , \37082 , \37083 , \37084 , \37085 , \37086 , \37087 , \37088 , \37089 , \37090 ,
         \37091 , \37092 , \37093 , \37094 , \37095 , \37096 , \37097 , \37098 , \37099 , \37100 ,
         \37101 , \37102 , \37103 , \37104 , \37105 , \37106 , \37107 , \37108 , \37109 , \37110 ,
         \37111 , \37112 , \37113 , \37114 , \37115 , \37116 , \37117 , \37118 , \37119 , \37120 ,
         \37121 , \37122 , \37123 , \37124 , \37125 , \37126 , \37127 , \37128 , \37129 , \37130 ,
         \37131 , \37132 , \37133 , \37134 , \37135 , \37136 , \37137 , \37138 , \37139 , \37140 ,
         \37141 , \37142 , \37143 , \37144 , \37145 , \37146 , \37147 , \37148 , \37149 , \37150 ,
         \37151 , \37152 , \37153 , \37154 , \37155 , \37156 , \37157 , \37158 , \37159 , \37160 ,
         \37161 , \37162 , \37163 , \37164 , \37165 , \37166 , \37167 , \37168 , \37169 , \37170 ,
         \37171 , \37172 , \37173 , \37174 , \37175 , \37176 , \37177 , \37178 , \37179 , \37180 ,
         \37181 , \37182 , \37183 , \37184 , \37185 , \37186 , \37187 , \37188 , \37189 , \37190 ,
         \37191 , \37192 , \37193 , \37194 , \37195 , \37196 , \37197 , \37198 , \37199 , \37200 ,
         \37201 , \37202 , \37203 , \37204 , \37205 , \37206 , \37207 , \37208 , \37209 , \37210 ,
         \37211 , \37212 , \37213 , \37214 , \37215 , \37216 , \37217 , \37218 , \37219 , \37220 ,
         \37221 , \37222 , \37223 , \37224 , \37225 , \37226 , \37227 , \37228 , \37229 , \37230 ,
         \37231 , \37232 , \37233 , \37234 , \37235 , \37236 , \37237 , \37238 , \37239 , \37240 ,
         \37241 , \37242 , \37243 , \37244 , \37245 , \37246 , \37247 , \37248 , \37249 , \37250 ,
         \37251 , \37252 , \37253 , \37254 , \37255 , \37256 , \37257 , \37258 , \37259 , \37260 ,
         \37261 , \37262 , \37263 , \37264 , \37265 , \37266 , \37267 , \37268 , \37269 , \37270 ,
         \37271 , \37272 , \37273 , \37274 , \37275 , \37276 , \37277 , \37278 , \37279 , \37280 ,
         \37281 , \37282 , \37283 , \37284 , \37285 , \37286 , \37287 , \37288 , \37289 , \37290 ,
         \37291 , \37292 , \37293 , \37294 , \37295 , \37296 , \37297 , \37298 , \37299 , \37300 ,
         \37301 , \37302 , \37303 , \37304 , \37305 , \37306 , \37307 , \37308 , \37309 , \37310 ,
         \37311 , \37312 , \37313 , \37314 , \37315 , \37316 , \37317 , \37318 , \37319 , \37320 ,
         \37321 , \37322 , \37323 , \37324 , \37325 , \37326 , \37327 , \37328 , \37329 , \37330 ,
         \37331 , \37332 , \37333 , \37334 , \37335 , \37336 , \37337 , \37338 , \37339 , \37340 ,
         \37341 , \37342 , \37343 , \37344 , \37345 , \37346 , \37347 , \37348 , \37349 , \37350 ,
         \37351 , \37352 , \37353 , \37354 , \37355 , \37356 , \37357 , \37358 , \37359 , \37360 ,
         \37361 , \37362 , \37363 , \37364 , \37365 , \37366 , \37367 , \37368 , \37369 , \37370 ,
         \37371 , \37372 , \37373 , \37374 , \37375 , \37376 , \37377 , \37378 , \37379 , \37380 ,
         \37381 , \37382 , \37383 , \37384 , \37385 , \37386 , \37387 , \37388 , \37389 , \37390 ,
         \37391 , \37392 , \37393 , \37394 , \37395 , \37396 , \37397 , \37398 , \37399 , \37400 ,
         \37401 , \37402 , \37403 , \37404 , \37405 , \37406 , \37407 , \37408 , \37409 , \37410 ,
         \37411 , \37412 , \37413 , \37414 , \37415 , \37416 , \37417 , \37418 , \37419 , \37420 ,
         \37421 , \37422 , \37423 , \37424 , \37425 , \37426 , \37427 , \37428 , \37429 , \37430 ,
         \37431 , \37432 , \37433 , \37434 , \37435 , \37436 , \37437 , \37438 , \37439 , \37440 ,
         \37441 , \37442 , \37443 , \37444 , \37445 , \37446 , \37447 , \37448 , \37449 , \37450 ,
         \37451 , \37452 , \37453 , \37454 , \37455 , \37456 , \37457 , \37458 , \37459 , \37460 ,
         \37461 , \37462 , \37463 , \37464 , \37465 , \37466 , \37467 , \37468 , \37469 , \37470 ,
         \37471 , \37472 , \37473 , \37474 , \37475 , \37476 , \37477 , \37478 , \37479 , \37480 ,
         \37481 , \37482 , \37483 , \37484 , \37485 , \37486 , \37487 , \37488 , \37489 , \37490 ,
         \37491 , \37492 , \37493 , \37494 , \37495 , \37496 , \37497 , \37498 , \37499 , \37500 ,
         \37501 , \37502 , \37503 , \37504 , \37505 , \37506 , \37507 , \37508 , \37509 , \37510 ,
         \37511 , \37512 , \37513 , \37514 , \37515 , \37516 , \37517 , \37518 , \37519 , \37520 ,
         \37521 , \37522 , \37523 , \37524 , \37525 , \37526 , \37527 , \37528 , \37529 , \37530 ,
         \37531 , \37532 , \37533 , \37534 , \37535 , \37536 , \37537 , \37538 , \37539 , \37540 ,
         \37541 , \37542 , \37543 , \37544 , \37545 , \37546 , \37547 , \37548 , \37549 , \37550 ,
         \37551 , \37552 , \37553 , \37554 , \37555 , \37556 , \37557 , \37558 , \37559 , \37560 ,
         \37561 , \37562 , \37563 , \37564 , \37565 , \37566 , \37567 , \37568 , \37569 , \37570 ,
         \37571 , \37572 , \37573 , \37574 , \37575 , \37576 , \37577 , \37578 , \37579 , \37580 ,
         \37581 , \37582 , \37583 , \37584 , \37585 , \37586 , \37587 , \37588 , \37589 , \37590 ,
         \37591 , \37592 , \37593 , \37594 , \37595 , \37596 , \37597 , \37598 , \37599 , \37600 ,
         \37601 , \37602 , \37603 , \37604 , \37605 , \37606 , \37607 , \37608 , \37609 , \37610 ,
         \37611 , \37612 , \37613 , \37614 , \37615 , \37616 , \37617 , \37618 , \37619 , \37620 ,
         \37621 , \37622 , \37623 , \37624 , \37625 , \37626 , \37627 , \37628 , \37629 , \37630 ,
         \37631 , \37632 , \37633 , \37634 , \37635 , \37636 , \37637 , \37638 , \37639 , \37640 ,
         \37641 , \37642 , \37643 , \37644 , \37645 , \37646 , \37647 , \37648 , \37649 , \37650 ,
         \37651 , \37652 , \37653 , \37654 , \37655 , \37656 , \37657 , \37658 , \37659 , \37660 ,
         \37661 , \37662 , \37663 , \37664 , \37665 , \37666 , \37667 , \37668 , \37669 , \37670 ,
         \37671 , \37672 , \37673 , \37674 , \37675 , \37676 , \37677 , \37678 , \37679 , \37680 ,
         \37681 , \37682 , \37683 , \37684 , \37685 , \37686 , \37687 , \37688 , \37689 , \37690 ,
         \37691 , \37692 , \37693 , \37694 , \37695 , \37696 , \37697 , \37698 , \37699 , \37700 ,
         \37701 , \37702 , \37703 , \37704 , \37705 , \37706 , \37707 , \37708 , \37709 , \37710 ,
         \37711 , \37712 , \37713 , \37714 , \37715 , \37716 , \37717 , \37718 , \37719 , \37720 ,
         \37721 , \37722 , \37723 , \37724 , \37725 , \37726 , \37727 , \37728 , \37729 , \37730 ,
         \37731 , \37732 , \37733 , \37734 , \37735 , \37736 , \37737 , \37738 , \37739 , \37740 ,
         \37741 , \37742 , \37743 , \37744 , \37745 , \37746 , \37747 , \37748 , \37749 , \37750 ,
         \37751 , \37752 , \37753 , \37754 , \37755 , \37756 , \37757 , \37758 , \37759 , \37760 ,
         \37761 , \37762 , \37763 , \37764 , \37765 , \37766 , \37767 , \37768 , \37769 , \37770 ,
         \37771 , \37772 , \37773 , \37774 , \37775 , \37776 , \37777 , \37778 , \37779 , \37780 ,
         \37781 , \37782 , \37783 , \37784 , \37785 , \37786 , \37787 , \37788 , \37789 , \37790 ,
         \37791 , \37792 , \37793 , \37794 , \37795 , \37796 , \37797 , \37798 , \37799 , \37800 ,
         \37801 , \37802 , \37803 , \37804 , \37805 , \37806 , \37807 , \37808 , \37809 , \37810 ,
         \37811 , \37812 , \37813 , \37814 , \37815 , \37816 , \37817 , \37818 , \37819 , \37820 ,
         \37821 , \37822 , \37823 , \37824 , \37825 , \37826 , \37827 , \37828 , \37829 , \37830 ,
         \37831 , \37832 , \37833 , \37834 , \37835 , \37836 , \37837 , \37838 , \37839 , \37840 ,
         \37841 , \37842 , \37843 , \37844 , \37845 , \37846 , \37847 , \37848 , \37849 , \37850 ,
         \37851 , \37852 , \37853 , \37854 , \37855 , \37856 , \37857 , \37858 , \37859 , \37860 ,
         \37861 , \37862 , \37863 , \37864 , \37865 , \37866 , \37867 , \37868 , \37869 , \37870 ,
         \37871 , \37872 , \37873 , \37874 , \37875 , \37876 , \37877 , \37878 , \37879 , \37880 ,
         \37881 , \37882 , \37883 , \37884 , \37885 , \37886 , \37887 , \37888 , \37889 , \37890 ,
         \37891 , \37892 , \37893 , \37894 , \37895 , \37896 , \37897 , \37898 , \37899 , \37900 ,
         \37901 , \37902 , \37903 , \37904 , \37905 , \37906 , \37907 , \37908 , \37909 , \37910 ,
         \37911 , \37912 , \37913 , \37914 , \37915 , \37916 , \37917 , \37918 , \37919 , \37920 ,
         \37921 , \37922 , \37923 , \37924 , \37925 , \37926 , \37927 , \37928 , \37929 , \37930 ,
         \37931 , \37932 , \37933 , \37934 , \37935 , \37936 , \37937 , \37938 , \37939 , \37940 ,
         \37941 , \37942 , \37943 , \37944 , \37945 , \37946 , \37947 , \37948 , \37949 , \37950 ,
         \37951 , \37952 , \37953 , \37954 , \37955 , \37956 , \37957 , \37958 , \37959 , \37960 ,
         \37961 , \37962 , \37963 , \37964 , \37965 , \37966 , \37967 , \37968 , \37969 , \37970 ,
         \37971 , \37972 , \37973 , \37974 , \37975 , \37976 , \37977 , \37978 , \37979 , \37980 ,
         \37981 , \37982 , \37983 , \37984 , \37985 , \37986 , \37987 , \37988 , \37989 , \37990 ,
         \37991 , \37992 , \37993 , \37994 , \37995 , \37996 , \37997 , \37998 , \37999 , \38000 ,
         \38001 , \38002 , \38003 , \38004 , \38005 , \38006 , \38007 , \38008 , \38009 , \38010 ,
         \38011 , \38012 , \38013 , \38014 , \38015 , \38016 , \38017 , \38018 , \38019 , \38020 ,
         \38021 , \38022 , \38023 , \38024 , \38025 , \38026 , \38027 , \38028 , \38029 , \38030 ,
         \38031 , \38032 , \38033 , \38034 , \38035 , \38036 , \38037 , \38038 , \38039 , \38040 ,
         \38041 , \38042 , \38043 , \38044 , \38045 , \38046 , \38047 , \38048 , \38049 , \38050 ,
         \38051 , \38052 , \38053 , \38054 , \38055 , \38056 , \38057 , \38058 , \38059 , \38060 ,
         \38061 , \38062 , \38063 , \38064 , \38065 , \38066 , \38067 , \38068 , \38069 , \38070 ,
         \38071 , \38072 , \38073 , \38074 , \38075 , \38076 , \38077 , \38078 , \38079 , \38080 ,
         \38081 , \38082 , \38083 , \38084 , \38085 , \38086 , \38087 , \38088 , \38089 , \38090 ,
         \38091 , \38092 , \38093 , \38094 , \38095 , \38096 , \38097 , \38098 , \38099 , \38100 ,
         \38101 , \38102 , \38103 , \38104 , \38105 , \38106 , \38107 , \38108 , \38109 , \38110 ,
         \38111 , \38112 , \38113 , \38114 , \38115 , \38116 , \38117 , \38118 , \38119 , \38120 ,
         \38121 , \38122 , \38123 , \38124 , \38125 , \38126 , \38127 , \38128 , \38129 , \38130 ,
         \38131 , \38132 , \38133 , \38134 , \38135 , \38136 , \38137 , \38138 , \38139 , \38140 ,
         \38141 , \38142 , \38143 , \38144 , \38145 , \38146 , \38147 , \38148 , \38149 , \38150 ,
         \38151 , \38152 , \38153 , \38154 , \38155 , \38156 , \38157 , \38158 , \38159 , \38160 ,
         \38161 , \38162 , \38163 , \38164 , \38165 , \38166 , \38167 , \38168 , \38169 , \38170 ,
         \38171 , \38172 , \38173 , \38174 , \38175 , \38176 , \38177 , \38178 , \38179 , \38180 ,
         \38181 , \38182 , \38183 , \38184 , \38185 , \38186 , \38187 , \38188 , \38189 , \38190 ,
         \38191 , \38192 , \38193 , \38194 , \38195 , \38196 , \38197 , \38198 , \38199 , \38200 ,
         \38201 , \38202 , \38203 , \38204 , \38205 , \38206 , \38207 , \38208 , \38209 , \38210 ,
         \38211 , \38212 , \38213 , \38214 , \38215 , \38216 , \38217 , \38218 , \38219 , \38220 ,
         \38221 , \38222 , \38223 , \38224 , \38225 , \38226 , \38227 , \38228 , \38229 , \38230 ,
         \38231 , \38232 , \38233 , \38234 , \38235 , \38236 , \38237 , \38238 , \38239 , \38240 ,
         \38241 , \38242 , \38243 , \38244 , \38245 , \38246 , \38247 , \38248 , \38249 , \38250 ,
         \38251 , \38252 , \38253 , \38254 , \38255 , \38256 , \38257 , \38258 , \38259 , \38260 ,
         \38261 , \38262 , \38263 , \38264 , \38265 , \38266 , \38267 , \38268 , \38269 , \38270 ,
         \38271 , \38272 , \38273 , \38274 , \38275 , \38276 , \38277 , \38278 , \38279 , \38280 ,
         \38281 , \38282 , \38283 , \38284 , \38285 , \38286 , \38287 , \38288 , \38289 , \38290 ,
         \38291 , \38292 , \38293 , \38294 , \38295 , \38296 , \38297 , \38298 , \38299 , \38300 ,
         \38301 , \38302 , \38303 , \38304 , \38305 , \38306 , \38307 , \38308 , \38309 , \38310 ,
         \38311 , \38312 , \38313 , \38314 , \38315 , \38316 , \38317 , \38318 , \38319 , \38320 ,
         \38321 , \38322 , \38323 , \38324 , \38325 , \38326 , \38327 , \38328 , \38329 , \38330 ,
         \38331 , \38332 , \38333 , \38334 , \38335 , \38336 , \38337 , \38338 , \38339 , \38340 ,
         \38341 , \38342 , \38343 , \38344 , \38345 , \38346 , \38347 , \38348 , \38349 , \38350 ,
         \38351 , \38352 , \38353 , \38354 , \38355 , \38356 , \38357 , \38358 , \38359 , \38360 ,
         \38361 , \38362 , \38363 , \38364 , \38365 , \38366 , \38367 , \38368 , \38369 , \38370 ,
         \38371 , \38372 , \38373 , \38374 , \38375 , \38376 , \38377 , \38378 , \38379 , \38380 ,
         \38381 , \38382 , \38383 , \38384 , \38385 , \38386 , \38387 , \38388 , \38389 , \38390 ,
         \38391 , \38392 , \38393 , \38394 , \38395 , \38396 , \38397 , \38398 , \38399 , \38400 ,
         \38401 , \38402 , \38403 , \38404 , \38405 , \38406 , \38407 , \38408 , \38409 , \38410 ,
         \38411 , \38412 , \38413 , \38414 , \38415 , \38416 , \38417 , \38418 , \38419 , \38420 ,
         \38421 , \38422 , \38423 , \38424 , \38425 , \38426 , \38427 , \38428 , \38429 , \38430 ,
         \38431 , \38432 , \38433 , \38434 , \38435 , \38436 , \38437 , \38438 , \38439 , \38440 ,
         \38441 , \38442 , \38443 , \38444 , \38445 , \38446 , \38447 , \38448 , \38449 , \38450 ,
         \38451 , \38452 , \38453 , \38454 , \38455 , \38456 , \38457 , \38458 , \38459 , \38460 ,
         \38461 , \38462 , \38463 , \38464 , \38465 , \38466 , \38467 , \38468 , \38469 , \38470 ,
         \38471 , \38472 , \38473 , \38474 , \38475 , \38476 , \38477 , \38478 , \38479 , \38480 ,
         \38481 , \38482 , \38483 , \38484 , \38485 , \38486 , \38487 , \38488 , \38489 , \38490 ,
         \38491 , \38492 , \38493 , \38494 , \38495 , \38496 , \38497 , \38498 , \38499 , \38500 ,
         \38501 , \38502 , \38503 , \38504 , \38505 , \38506 , \38507 , \38508 , \38509 , \38510 ,
         \38511 , \38512 , \38513 , \38514 , \38515 , \38516 , \38517 , \38518 , \38519 , \38520 ,
         \38521 , \38522 , \38523 , \38524 , \38525 , \38526 , \38527 , \38528 , \38529 , \38530 ,
         \38531 , \38532 , \38533 , \38534 , \38535 , \38536 , \38537 , \38538 , \38539 , \38540 ,
         \38541 , \38542 , \38543 , \38544 , \38545 , \38546 , \38547 , \38548 , \38549 , \38550 ,
         \38551 , \38552 , \38553 , \38554 , \38555 , \38556 , \38557 , \38558 , \38559 , \38560 ,
         \38561 , \38562 , \38563 , \38564 , \38565 , \38566 , \38567 , \38568 , \38569 , \38570 ,
         \38571 , \38572 , \38573 , \38574 , \38575 , \38576 , \38577 , \38578 , \38579 , \38580 ,
         \38581 , \38582 , \38583 , \38584 , \38585 , \38586 , \38587 , \38588 , \38589 , \38590 ,
         \38591 , \38592 , \38593 , \38594 , \38595 , \38596 , \38597 , \38598 , \38599 , \38600 ,
         \38601 , \38602 , \38603 , \38604 , \38605 , \38606 , \38607 , \38608 , \38609 , \38610 ,
         \38611 , \38612 , \38613 , \38614 , \38615 , \38616 , \38617 , \38618 , \38619 , \38620 ,
         \38621 , \38622 , \38623 , \38624 , \38625 , \38626 , \38627 , \38628 , \38629 , \38630 ,
         \38631 , \38632 , \38633 , \38634 , \38635 , \38636 , \38637 , \38638 , \38639 , \38640 ,
         \38641 , \38642 , \38643 , \38644 , \38645 , \38646 , \38647 , \38648 , \38649 , \38650 ,
         \38651 , \38652 , \38653 , \38654 , \38655 , \38656 , \38657 , \38658 , \38659 , \38660 ,
         \38661 , \38662 , \38663 , \38664 , \38665 , \38666 , \38667 , \38668 , \38669 , \38670 ,
         \38671 , \38672 , \38673 , \38674 , \38675 , \38676 , \38677 , \38678 , \38679 , \38680 ,
         \38681 , \38682 , \38683 , \38684 , \38685 , \38686 , \38687 , \38688 , \38689 , \38690 ,
         \38691 , \38692 , \38693 , \38694 , \38695 , \38696 , \38697 , \38698 , \38699 , \38700 ,
         \38701 , \38702 , \38703 , \38704 , \38705 , \38706 , \38707 , \38708 , \38709 , \38710 ,
         \38711 , \38712 , \38713 , \38714 , \38715 , \38716 , \38717 , \38718 , \38719 , \38720 ,
         \38721 , \38722 , \38723 , \38724 , \38725 , \38726 , \38727 , \38728 , \38729 , \38730 ,
         \38731 , \38732 , \38733 , \38734 , \38735 , \38736 , \38737 , \38738 , \38739 , \38740 ,
         \38741 , \38742 , \38743 , \38744 , \38745 , \38746 , \38747 , \38748 , \38749 , \38750 ,
         \38751 , \38752 , \38753 , \38754 , \38755 , \38756 , \38757 , \38758 , \38759 , \38760 ,
         \38761 , \38762 , \38763 , \38764 , \38765 , \38766 , \38767 , \38768 , \38769 , \38770 ,
         \38771 , \38772 , \38773 , \38774 , \38775 , \38776 , \38777 , \38778 , \38779 , \38780 ,
         \38781 , \38782 , \38783 , \38784 , \38785 , \38786 , \38787 , \38788 , \38789 , \38790 ,
         \38791 , \38792 , \38793 , \38794 , \38795 , \38796 , \38797 , \38798 , \38799 , \38800 ,
         \38801 , \38802 , \38803 , \38804 , \38805 , \38806 , \38807 , \38808 , \38809 , \38810 ,
         \38811 , \38812 , \38813 , \38814 , \38815 , \38816 , \38817 , \38818 , \38819 , \38820 ,
         \38821 , \38822 , \38823 , \38824 , \38825 , \38826 , \38827 , \38828 , \38829 , \38830 ,
         \38831 , \38832 , \38833 , \38834 , \38835 , \38836 , \38837 , \38838 , \38839 , \38840 ,
         \38841 , \38842 , \38843 , \38844 , \38845 , \38846 , \38847 , \38848 , \38849 , \38850 ,
         \38851 , \38852 , \38853 , \38854 , \38855 , \38856 , \38857 , \38858 , \38859 , \38860 ,
         \38861 , \38862 , \38863 , \38864 , \38865 , \38866 , \38867 , \38868 , \38869 , \38870 ,
         \38871 , \38872 , \38873 , \38874 , \38875 , \38876 , \38877 , \38878 , \38879 , \38880 ,
         \38881 , \38882 , \38883 , \38884 , \38885 , \38886 , \38887 , \38888 , \38889 , \38890 ,
         \38891 , \38892 , \38893 , \38894 , \38895 , \38896 , \38897 , \38898 , \38899 , \38900 ,
         \38901 , \38902 , \38903 , \38904 , \38905 , \38906 , \38907 , \38908 , \38909 , \38910 ,
         \38911 , \38912 , \38913 , \38914 , \38915 , \38916 , \38917 , \38918 , \38919 , \38920 ,
         \38921 , \38922 , \38923 , \38924 , \38925 , \38926 , \38927 , \38928 , \38929 , \38930 ,
         \38931 , \38932 , \38933 , \38934 , \38935 , \38936 , \38937 , \38938 , \38939 , \38940 ,
         \38941 , \38942 , \38943 , \38944 , \38945 , \38946 , \38947 , \38948 , \38949 , \38950 ,
         \38951 , \38952 , \38953 , \38954 , \38955 , \38956 , \38957 , \38958 , \38959 , \38960 ,
         \38961 , \38962 , \38963 , \38964 , \38965 , \38966 , \38967 , \38968 , \38969 , \38970 ,
         \38971 , \38972 , \38973 , \38974 , \38975 , \38976 , \38977 , \38978 , \38979 , \38980 ,
         \38981 , \38982 , \38983 , \38984 , \38985 , \38986 , \38987 , \38988 , \38989 , \38990 ,
         \38991 , \38992 , \38993 , \38994 , \38995 , \38996 , \38997 , \38998 , \38999 , \39000 ,
         \39001 , \39002 , \39003 , \39004 , \39005 , \39006 , \39007 , \39008 , \39009 , \39010 ,
         \39011 , \39012 , \39013 , \39014 , \39015 , \39016 , \39017 , \39018 , \39019 , \39020 ,
         \39021 , \39022 , \39023 , \39024 , \39025 , \39026 , \39027 , \39028 , \39029 , \39030 ,
         \39031 , \39032 , \39033 , \39034 , \39035 , \39036 , \39037 , \39038 , \39039 , \39040 ,
         \39041 , \39042 , \39043 , \39044 , \39045 , \39046 , \39047 , \39048 , \39049 , \39050 ,
         \39051 , \39052 , \39053 , \39054 , \39055 , \39056 , \39057 , \39058 , \39059 , \39060 ,
         \39061 , \39062 , \39063 , \39064 , \39065 , \39066 , \39067 , \39068 , \39069 , \39070 ,
         \39071 , \39072 , \39073 , \39074 , \39075 , \39076 , \39077 , \39078 , \39079 , \39080 ,
         \39081 , \39082 , \39083 , \39084 , \39085 , \39086 , \39087 , \39088 , \39089 , \39090 ,
         \39091 , \39092 , \39093 , \39094 , \39095 , \39096 , \39097 , \39098 , \39099 , \39100 ,
         \39101 , \39102 , \39103 , \39104 , \39105 , \39106 , \39107 , \39108 , \39109 , \39110 ,
         \39111 , \39112 , \39113 , \39114 , \39115 , \39116 , \39117 , \39118 , \39119 , \39120 ,
         \39121 , \39122 , \39123 , \39124 , \39125 , \39126 , \39127 , \39128 , \39129 , \39130 ,
         \39131 , \39132 , \39133 , \39134 , \39135 , \39136 , \39137 , \39138 , \39139 , \39140 ,
         \39141 , \39142 , \39143 , \39144 , \39145 , \39146 , \39147 , \39148 , \39149 , \39150 ,
         \39151 , \39152 , \39153 , \39154 , \39155 , \39156 , \39157 , \39158 , \39159 , \39160 ,
         \39161 , \39162 , \39163 , \39164 , \39165 , \39166 , \39167 , \39168 , \39169 , \39170 ,
         \39171 , \39172 , \39173 , \39174 , \39175 , \39176 , \39177 , \39178 , \39179 , \39180 ,
         \39181 , \39182 , \39183 , \39184 , \39185 , \39186 , \39187 , \39188 , \39189 , \39190 ,
         \39191 , \39192 , \39193 , \39194 , \39195 , \39196 , \39197 , \39198 , \39199 , \39200 ,
         \39201 , \39202 , \39203 , \39204 , \39205 , \39206 , \39207 , \39208 , \39209 , \39210 ,
         \39211 , \39212 , \39213 , \39214 , \39215 , \39216 , \39217 , \39218 , \39219 , \39220 ,
         \39221 , \39222 , \39223 , \39224 , \39225 , \39226 , \39227 , \39228 , \39229 , \39230 ,
         \39231 , \39232 , \39233 , \39234 , \39235 , \39236 , \39237 , \39238 , \39239 , \39240 ,
         \39241 , \39242 , \39243 , \39244 , \39245 , \39246 , \39247 , \39248 , \39249 , \39250 ,
         \39251 , \39252 , \39253 , \39254 , \39255 , \39256 , \39257 , \39258 , \39259 , \39260 ,
         \39261 , \39262 , \39263 , \39264 , \39265 , \39266 , \39267 , \39268 , \39269 , \39270 ,
         \39271 , \39272 , \39273 , \39274 , \39275 , \39276 , \39277 , \39278 , \39279 , \39280 ,
         \39281 , \39282 , \39283 , \39284 , \39285 , \39286 , \39287 , \39288 , \39289 , \39290 ,
         \39291 , \39292 , \39293 , \39294 , \39295 , \39296 , \39297 , \39298 , \39299 , \39300 ,
         \39301 , \39302 , \39303 , \39304 , \39305 , \39306 , \39307 , \39308 , \39309 , \39310 ,
         \39311 , \39312 , \39313 , \39314 , \39315 , \39316 , \39317 , \39318 , \39319 , \39320 ,
         \39321 , \39322 , \39323 , \39324 , \39325 , \39326 , \39327 , \39328 , \39329 , \39330 ,
         \39331 , \39332 , \39333 , \39334 , \39335 , \39336 , \39337 , \39338 , \39339 , \39340 ,
         \39341 , \39342 , \39343 , \39344 , \39345 , \39346 , \39347 , \39348 , \39349 , \39350 ,
         \39351 , \39352 , \39353 , \39354 , \39355 , \39356 , \39357 , \39358 , \39359 , \39360 ,
         \39361 , \39362 , \39363 , \39364 , \39365 , \39366 , \39367 , \39368 , \39369 , \39370 ,
         \39371 , \39372 , \39373 , \39374 , \39375 , \39376 , \39377 , \39378 , \39379 , \39380 ,
         \39381 , \39382 , \39383 , \39384 , \39385 , \39386 , \39387 , \39388 , \39389 , \39390 ,
         \39391 , \39392 , \39393 , \39394 , \39395 , \39396 , \39397 , \39398 , \39399 , \39400 ,
         \39401 , \39402 , \39403 , \39404 , \39405 , \39406 , \39407 , \39408 , \39409 , \39410 ,
         \39411 , \39412 , \39413 , \39414 , \39415 , \39416 , \39417 , \39418 , \39419 , \39420 ,
         \39421 , \39422 , \39423 , \39424 , \39425 , \39426 , \39427 , \39428 , \39429 , \39430 ,
         \39431 , \39432 , \39433 , \39434 , \39435 , \39436 , \39437 , \39438 , \39439 , \39440 ,
         \39441 , \39442 , \39443 , \39444 , \39445 , \39446 , \39447 , \39448 , \39449 , \39450 ,
         \39451 , \39452 , \39453 , \39454 , \39455 , \39456 , \39457 , \39458 , \39459 , \39460 ,
         \39461 , \39462 , \39463 , \39464 , \39465 , \39466 , \39467 , \39468 , \39469 , \39470 ,
         \39471 , \39472 , \39473 , \39474 , \39475 , \39476 , \39477 , \39478 , \39479 , \39480 ,
         \39481 , \39482 , \39483 , \39484 , \39485 , \39486 , \39487 , \39488 , \39489 , \39490 ,
         \39491 , \39492 , \39493 , \39494 , \39495 , \39496 , \39497 , \39498 , \39499 , \39500 ,
         \39501 , \39502 , \39503 , \39504 , \39505 , \39506 , \39507 , \39508 , \39509 , \39510 ,
         \39511 , \39512 , \39513 , \39514 , \39515 , \39516 , \39517 , \39518 , \39519 , \39520 ,
         \39521 , \39522 , \39523 , \39524 , \39525 , \39526 , \39527 , \39528 , \39529 , \39530 ,
         \39531 , \39532 , \39533 , \39534 , \39535 , \39536 , \39537 , \39538 , \39539 , \39540 ,
         \39541 , \39542 , \39543 , \39544 , \39545 , \39546 , \39547 , \39548 , \39549 , \39550 ,
         \39551 , \39552 , \39553 , \39554 , \39555 , \39556 , \39557 , \39558 , \39559 , \39560 ,
         \39561 , \39562 , \39563 , \39564 , \39565 , \39566 , \39567 , \39568 , \39569 , \39570 ,
         \39571 , \39572 , \39573 , \39574 , \39575 , \39576 , \39577 , \39578 , \39579 , \39580 ,
         \39581 , \39582 , \39583 , \39584 , \39585 , \39586 , \39587 , \39588 , \39589 , \39590 ,
         \39591 , \39592 , \39593 , \39594 , \39595 , \39596 , \39597 , \39598 , \39599 , \39600 ,
         \39601 , \39602 , \39603 , \39604 , \39605 , \39606 , \39607 , \39608 , \39609 , \39610 ,
         \39611 , \39612 , \39613 , \39614 , \39615 , \39616 , \39617 , \39618 , \39619 , \39620 ,
         \39621 , \39622 , \39623 , \39624 , \39625 , \39626 , \39627 , \39628 , \39629 , \39630 ,
         \39631 , \39632 , \39633 , \39634 , \39635 , \39636 , \39637 , \39638 , \39639 , \39640 ,
         \39641 , \39642 , \39643 , \39644 , \39645 , \39646 , \39647 , \39648 , \39649 , \39650 ,
         \39651 , \39652 , \39653 , \39654 , \39655 , \39656 , \39657 , \39658 , \39659 , \39660 ,
         \39661 , \39662 , \39663 , \39664 , \39665 , \39666 , \39667 , \39668 , \39669 , \39670 ,
         \39671 , \39672 , \39673 , \39674 , \39675 , \39676 , \39677 , \39678 , \39679 , \39680 ,
         \39681 , \39682 , \39683 , \39684 , \39685 , \39686 , \39687 , \39688 , \39689 , \39690 ,
         \39691 , \39692 , \39693 , \39694 , \39695 , \39696 , \39697 , \39698 , \39699 , \39700 ,
         \39701 , \39702 , \39703 , \39704 , \39705 , \39706 , \39707 , \39708 , \39709 , \39710 ,
         \39711 , \39712 , \39713 , \39714 , \39715 , \39716 , \39717 , \39718 , \39719 , \39720 ,
         \39721 , \39722 , \39723 , \39724 , \39725 , \39726 , \39727 , \39728 , \39729 , \39730 ,
         \39731 , \39732 , \39733 , \39734 , \39735 , \39736 , \39737 , \39738 , \39739 , \39740 ,
         \39741 , \39742 , \39743 , \39744 , \39745 , \39746 , \39747 , \39748 , \39749 , \39750 ,
         \39751 , \39752 , \39753 , \39754 , \39755 , \39756 , \39757 , \39758 , \39759 , \39760 ,
         \39761 , \39762 , \39763 , \39764 , \39765 , \39766 , \39767 , \39768 , \39769 , \39770 ,
         \39771 , \39772 , \39773 , \39774 , \39775 , \39776 , \39777 , \39778 , \39779 , \39780 ,
         \39781 , \39782 , \39783 , \39784 , \39785 , \39786 , \39787 , \39788 , \39789 , \39790 ,
         \39791 , \39792 , \39793 , \39794 , \39795 , \39796 , \39797 , \39798 , \39799 , \39800 ,
         \39801 , \39802 , \39803 , \39804 , \39805 , \39806 , \39807 , \39808 , \39809 , \39810 ,
         \39811 , \39812 , \39813 , \39814 , \39815 , \39816 , \39817 , \39818 , \39819 , \39820 ,
         \39821 , \39822 , \39823 , \39824 , \39825 , \39826 , \39827 , \39828 , \39829 , \39830 ,
         \39831 , \39832 , \39833 , \39834 , \39835 , \39836 , \39837 , \39838 , \39839 , \39840 ,
         \39841 , \39842 , \39843 , \39844 , \39845 , \39846 , \39847 , \39848 , \39849 , \39850 ,
         \39851 , \39852 , \39853 , \39854 , \39855 , \39856 , \39857 , \39858 , \39859 , \39860 ,
         \39861 , \39862 , \39863 , \39864 , \39865 , \39866 , \39867 , \39868 , \39869 , \39870 ,
         \39871 , \39872 , \39873 , \39874 , \39875 , \39876 , \39877 , \39878 , \39879 , \39880 ,
         \39881 , \39882 , \39883 , \39884 , \39885 , \39886 , \39887 , \39888 , \39889 , \39890 ,
         \39891 , \39892 , \39893 , \39894 , \39895 , \39896 , \39897 , \39898 , \39899 , \39900 ,
         \39901 , \39902 , \39903 , \39904 , \39905 , \39906 , \39907 , \39908 , \39909 , \39910 ,
         \39911 , \39912 , \39913 , \39914 , \39915 , \39916 , \39917 , \39918 , \39919 , \39920 ,
         \39921 , \39922 , \39923 , \39924 , \39925 , \39926 , \39927 , \39928 , \39929 , \39930 ,
         \39931 , \39932 , \39933 , \39934 , \39935 , \39936 , \39937 , \39938 , \39939 , \39940 ,
         \39941 , \39942 , \39943 , \39944 , \39945 , \39946 , \39947 , \39948 , \39949 , \39950 ,
         \39951 , \39952 , \39953 , \39954 , \39955 , \39956 , \39957 , \39958 , \39959 , \39960 ,
         \39961 , \39962 , \39963 , \39964 , \39965 , \39966 , \39967 , \39968 , \39969 , \39970 ,
         \39971 , \39972 , \39973 , \39974 , \39975 , \39976 , \39977 , \39978 , \39979 , \39980 ,
         \39981 , \39982 , \39983 , \39984 , \39985 , \39986 , \39987 , \39988 , \39989 , \39990 ,
         \39991 , \39992 , \39993 , \39994 , \39995 , \39996 , \39997 , \39998 , \39999 , \40000 ,
         \40001 , \40002 , \40003 , \40004 , \40005 , \40006 , \40007 , \40008 , \40009 , \40010 ,
         \40011 , \40012 , \40013 , \40014 , \40015 , \40016 , \40017 , \40018 , \40019 , \40020 ,
         \40021 , \40022 , \40023 , \40024 , \40025 , \40026 , \40027 , \40028 , \40029 , \40030 ,
         \40031 , \40032 , \40033 , \40034 , \40035 , \40036 , \40037 , \40038 , \40039 , \40040 ,
         \40041 , \40042 , \40043 , \40044 , \40045 , \40046 , \40047 , \40048 , \40049 , \40050 ,
         \40051 , \40052 , \40053 , \40054 , \40055 , \40056 , \40057 , \40058 , \40059 , \40060 ,
         \40061 , \40062 , \40063 , \40064 , \40065 , \40066 , \40067 , \40068 , \40069 , \40070 ,
         \40071 , \40072 , \40073 , \40074 , \40075 , \40076 , \40077 , \40078 , \40079 , \40080 ,
         \40081 , \40082 , \40083 , \40084 , \40085 , \40086 , \40087 , \40088 , \40089 , \40090 ,
         \40091 , \40092 , \40093 , \40094 , \40095 , \40096 , \40097 , \40098 , \40099 , \40100 ,
         \40101 , \40102 , \40103 , \40104 , \40105 , \40106 , \40107 , \40108 , \40109 , \40110 ,
         \40111 , \40112 , \40113 , \40114 , \40115 , \40116 , \40117 , \40118 , \40119 , \40120 ,
         \40121 , \40122 , \40123 , \40124 , \40125 , \40126 , \40127 , \40128 , \40129 , \40130 ,
         \40131 , \40132 , \40133 , \40134 , \40135 , \40136 , \40137 , \40138 , \40139 , \40140 ,
         \40141 , \40142 , \40143 , \40144 , \40145 , \40146 , \40147 , \40148 , \40149 , \40150 ,
         \40151 , \40152 , \40153 , \40154 , \40155 , \40156 , \40157 , \40158 , \40159 , \40160 ,
         \40161 , \40162 , \40163 , \40164 , \40165 , \40166 , \40167 , \40168 , \40169 , \40170 ,
         \40171 , \40172 , \40173 , \40174 , \40175 , \40176 , \40177 , \40178 , \40179 , \40180 ,
         \40181 , \40182 , \40183 , \40184 , \40185 , \40186 , \40187 , \40188 , \40189 , \40190 ,
         \40191 , \40192 , \40193 , \40194 , \40195 , \40196 , \40197 , \40198 , \40199 , \40200 ,
         \40201 , \40202 , \40203 , \40204 , \40205 , \40206 , \40207 , \40208 , \40209 , \40210 ,
         \40211 , \40212 , \40213 , \40214 , \40215 , \40216 , \40217 , \40218 , \40219 , \40220 ,
         \40221 , \40222 , \40223 , \40224 , \40225 , \40226 , \40227 , \40228 , \40229 , \40230 ,
         \40231 , \40232 , \40233 , \40234 , \40235 , \40236 , \40237 , \40238 , \40239 , \40240 ,
         \40241 , \40242 , \40243 , \40244 , \40245 , \40246 , \40247 , \40248 , \40249 , \40250 ,
         \40251 , \40252 , \40253 , \40254 , \40255 , \40256 , \40257 , \40258 , \40259 , \40260 ,
         \40261 , \40262 , \40263 , \40264 , \40265 , \40266 , \40267 , \40268 , \40269 , \40270 ,
         \40271 , \40272 , \40273 , \40274 , \40275 , \40276 , \40277 , \40278 , \40279 , \40280 ,
         \40281 , \40282 , \40283 , \40284 , \40285 , \40286 , \40287 , \40288 , \40289 , \40290 ,
         \40291 , \40292 , \40293 , \40294 , \40295 , \40296 , \40297 , \40298 , \40299 , \40300 ,
         \40301 , \40302 , \40303 , \40304 , \40305 , \40306 , \40307 , \40308 , \40309 , \40310 ,
         \40311 , \40312 , \40313 , \40314 , \40315 , \40316 , \40317 , \40318 , \40319 , \40320 ,
         \40321 , \40322 , \40323 , \40324 , \40325 , \40326 , \40327 , \40328 , \40329 , \40330 ,
         \40331 , \40332 , \40333 , \40334 , \40335 , \40336 , \40337 , \40338 , \40339 , \40340 ,
         \40341 , \40342 , \40343 , \40344 , \40345 , \40346 , \40347 , \40348 , \40349 , \40350 ,
         \40351 , \40352 , \40353 , \40354 , \40355 , \40356 , \40357 , \40358 , \40359 , \40360 ,
         \40361 , \40362 , \40363 , \40364 , \40365 , \40366 , \40367 , \40368 , \40369 , \40370 ,
         \40371 , \40372 , \40373 , \40374 , \40375 , \40376 , \40377 , \40378 , \40379 , \40380 ,
         \40381 , \40382 , \40383 , \40384 , \40385 , \40386 , \40387 , \40388 , \40389 , \40390 ,
         \40391 , \40392 , \40393 , \40394 , \40395 , \40396 , \40397 , \40398 , \40399 , \40400 ,
         \40401 , \40402 , \40403 , \40404 , \40405 , \40406 , \40407 , \40408 , \40409 , \40410 ,
         \40411 , \40412 , \40413 , \40414 , \40415 , \40416 , \40417 , \40418 , \40419 , \40420 ,
         \40421 , \40422 , \40423 , \40424 , \40425 , \40426 , \40427 , \40428 , \40429 , \40430 ,
         \40431 , \40432 , \40433 , \40434 , \40435 , \40436 , \40437 , \40438 , \40439 , \40440 ,
         \40441 , \40442 , \40443 , \40444 , \40445 , \40446 , \40447 , \40448 , \40449 , \40450 ,
         \40451 , \40452 , \40453 , \40454 , \40455 , \40456 , \40457 , \40458 , \40459 , \40460 ,
         \40461 , \40462 , \40463 , \40464 , \40465 , \40466 , \40467 , \40468 , \40469 , \40470 ,
         \40471 , \40472 , \40473 , \40474 , \40475 , \40476 , \40477 , \40478 , \40479 , \40480 ,
         \40481 , \40482 , \40483 , \40484 , \40485 , \40486 , \40487 , \40488 , \40489 , \40490 ,
         \40491 , \40492 , \40493 , \40494 , \40495 , \40496 , \40497 , \40498 , \40499 , \40500 ,
         \40501 , \40502 , \40503 , \40504 , \40505 , \40506 , \40507 , \40508 , \40509 , \40510 ,
         \40511 , \40512 , \40513 , \40514 , \40515 , \40516 , \40517 , \40518 , \40519 , \40520 ,
         \40521 , \40522 , \40523 , \40524 , \40525 , \40526 , \40527 , \40528 , \40529 , \40530 ,
         \40531 , \40532 , \40533 , \40534 , \40535 , \40536 , \40537 , \40538 , \40539 , \40540 ,
         \40541 , \40542 , \40543 , \40544 , \40545 , \40546 , \40547 , \40548 , \40549 , \40550 ,
         \40551 , \40552 , \40553 , \40554 , \40555 , \40556 , \40557 , \40558 , \40559 , \40560 ,
         \40561 , \40562 , \40563 , \40564 , \40565 , \40566 , \40567 , \40568 , \40569 , \40570 ,
         \40571 , \40572 , \40573 , \40574 , \40575 , \40576 , \40577 , \40578 , \40579 , \40580 ,
         \40581 , \40582 , \40583 , \40584 , \40585 , \40586 , \40587 , \40588 , \40589 , \40590 ,
         \40591 , \40592 , \40593 , \40594 , \40595 , \40596 , \40597 , \40598 , \40599 , \40600 ,
         \40601 , \40602 , \40603 , \40604 , \40605 , \40606 , \40607 , \40608 , \40609 , \40610 ,
         \40611 , \40612 , \40613 , \40614 , \40615 , \40616 , \40617 , \40618 , \40619 , \40620 ,
         \40621 , \40622 , \40623 , \40624 , \40625 , \40626 , \40627 , \40628 , \40629 , \40630 ,
         \40631 , \40632 , \40633 , \40634 , \40635 , \40636 , \40637 , \40638 , \40639 , \40640 ,
         \40641 , \40642 , \40643 , \40644 , \40645 , \40646 , \40647 , \40648 , \40649 , \40650 ,
         \40651 , \40652 , \40653 , \40654 , \40655 , \40656 , \40657 , \40658 , \40659 , \40660 ,
         \40661 , \40662 , \40663 , \40664 , \40665 , \40666 , \40667 , \40668 , \40669 , \40670 ,
         \40671 , \40672 , \40673 , \40674 , \40675 , \40676 , \40677 , \40678 , \40679 , \40680 ,
         \40681 , \40682 , \40683 , \40684 , \40685 , \40686 , \40687 , \40688 , \40689 , \40690 ,
         \40691 , \40692 , \40693 , \40694 , \40695 , \40696 , \40697 , \40698 , \40699 , \40700 ,
         \40701 , \40702 , \40703 , \40704 , \40705 , \40706 , \40707 , \40708 , \40709 , \40710 ,
         \40711 , \40712 , \40713 , \40714 , \40715 , \40716 , \40717 , \40718 , \40719 , \40720 ,
         \40721 , \40722 , \40723 , \40724 , \40725 , \40726 , \40727 , \40728 , \40729 , \40730 ,
         \40731 , \40732 , \40733 , \40734 , \40735 , \40736 , \40737 , \40738 , \40739 , \40740 ,
         \40741 , \40742 , \40743 , \40744 , \40745 , \40746 , \40747 , \40748 , \40749 , \40750 ,
         \40751 , \40752 , \40753 , \40754 , \40755 , \40756 , \40757 , \40758 , \40759 , \40760 ,
         \40761 , \40762 , \40763 , \40764 , \40765 , \40766 , \40767 , \40768 , \40769 , \40770 ,
         \40771 , \40772 , \40773 , \40774 , \40775 , \40776 , \40777 , \40778 , \40779 , \40780 ,
         \40781 , \40782 , \40783 , \40784 , \40785 , \40786 , \40787 , \40788 , \40789 , \40790 ,
         \40791 , \40792 , \40793 , \40794 , \40795 , \40796 , \40797 , \40798 , \40799 , \40800 ,
         \40801 , \40802 , \40803 , \40804 , \40805 , \40806 , \40807 , \40808 , \40809 , \40810 ,
         \40811 , \40812 , \40813 , \40814 , \40815 , \40816 , \40817 , \40818 , \40819 , \40820 ,
         \40821 , \40822 , \40823 , \40824 , \40825 , \40826 , \40827 , \40828 , \40829 , \40830 ,
         \40831 , \40832 , \40833 , \40834 , \40835 , \40836 , \40837 , \40838 , \40839 , \40840 ,
         \40841 , \40842 , \40843 , \40844 , \40845 , \40846 , \40847 , \40848 , \40849 , \40850 ,
         \40851 , \40852 , \40853 , \40854 , \40855 , \40856 , \40857 , \40858 , \40859 , \40860 ,
         \40861 , \40862 , \40863 , \40864 , \40865 , \40866 , \40867 , \40868 , \40869 , \40870 ,
         \40871 , \40872 , \40873 , \40874 , \40875 , \40876 , \40877 , \40878 , \40879 , \40880 ,
         \40881 , \40882 , \40883 , \40884 , \40885 , \40886 , \40887 , \40888 , \40889 , \40890 ,
         \40891 , \40892 , \40893 , \40894 , \40895 , \40896 , \40897 , \40898 , \40899 , \40900 ,
         \40901 , \40902 , \40903 , \40904 , \40905 , \40906 , \40907 , \40908 , \40909 , \40910 ,
         \40911 , \40912 , \40913 , \40914 , \40915 , \40916 , \40917 , \40918 , \40919 , \40920 ,
         \40921 , \40922 , \40923 , \40924 , \40925 , \40926 , \40927 , \40928 , \40929 , \40930 ,
         \40931 , \40932 , \40933 , \40934 , \40935 , \40936 , \40937 , \40938 , \40939 , \40940 ,
         \40941 , \40942 , \40943 , \40944 , \40945 , \40946 , \40947 , \40948 , \40949 , \40950 ,
         \40951 , \40952 , \40953 , \40954 , \40955 , \40956 , \40957 , \40958 , \40959 , \40960 ,
         \40961 , \40962 , \40963 , \40964 , \40965 , \40966 , \40967 , \40968 , \40969 , \40970 ,
         \40971 , \40972 , \40973 , \40974 , \40975 , \40976 , \40977 , \40978 , \40979 , \40980 ,
         \40981 , \40982 , \40983 , \40984 , \40985 , \40986 , \40987 , \40988 , \40989 , \40990 ,
         \40991 , \40992 , \40993 , \40994 , \40995 , \40996 , \40997 , \40998 , \40999 , \41000 ,
         \41001 , \41002 , \41003 , \41004 , \41005 , \41006 , \41007 , \41008 , \41009 , \41010 ,
         \41011 , \41012 , \41013 , \41014 , \41015 , \41016 , \41017 , \41018 , \41019 , \41020 ,
         \41021 , \41022 , \41023 , \41024 , \41025 , \41026 , \41027 , \41028 , \41029 , \41030 ,
         \41031 , \41032 , \41033 , \41034 , \41035 , \41036 , \41037 , \41038 , \41039 , \41040 ,
         \41041 , \41042 , \41043 , \41044 , \41045 , \41046 , \41047 , \41048 , \41049 , \41050 ,
         \41051 , \41052 , \41053 , \41054 , \41055 , \41056 , \41057 , \41058 , \41059 , \41060 ,
         \41061 , \41062 , \41063 , \41064 , \41065 , \41066 , \41067 , \41068 , \41069 , \41070 ,
         \41071 , \41072 , \41073 , \41074 , \41075 , \41076 , \41077 , \41078 , \41079 , \41080 ,
         \41081 , \41082 , \41083 , \41084 , \41085 , \41086 , \41087 , \41088 , \41089 , \41090 ,
         \41091 , \41092 , \41093 , \41094 , \41095 , \41096 , \41097 , \41098 , \41099 , \41100 ,
         \41101 , \41102 , \41103 , \41104 , \41105 , \41106 , \41107 , \41108 , \41109 , \41110 ,
         \41111 , \41112 , \41113 , \41114 , \41115 , \41116 , \41117 , \41118 , \41119 , \41120 ,
         \41121 , \41122 , \41123 , \41124 , \41125 , \41126 , \41127 , \41128 , \41129 , \41130 ,
         \41131 , \41132 , \41133 , \41134 , \41135 , \41136 , \41137 , \41138 , \41139 , \41140 ,
         \41141 , \41142 , \41143 , \41144 , \41145 , \41146 , \41147 , \41148 , \41149 , \41150 ,
         \41151 , \41152 , \41153 , \41154 , \41155 , \41156 , \41157 , \41158 , \41159 , \41160 ,
         \41161 , \41162 , \41163 , \41164 , \41165 , \41166 , \41167 , \41168 , \41169 , \41170 ,
         \41171 , \41172 , \41173 , \41174 , \41175 , \41176 , \41177 , \41178 , \41179 , \41180 ,
         \41181 , \41182 , \41183 , \41184 , \41185 , \41186 , \41187 , \41188 , \41189 , \41190 ,
         \41191 , \41192 , \41193 , \41194 , \41195 , \41196 , \41197 , \41198 , \41199 , \41200 ,
         \41201 , \41202 , \41203 , \41204 , \41205 , \41206 , \41207 , \41208 , \41209 , \41210 ,
         \41211 , \41212 , \41213 , \41214 , \41215 , \41216 , \41217 , \41218 , \41219 , \41220 ,
         \41221 , \41222 , \41223 , \41224 , \41225 , \41226 , \41227 , \41228 , \41229 , \41230 ,
         \41231 , \41232 , \41233 , \41234 , \41235 , \41236 , \41237 , \41238 , \41239 , \41240 ,
         \41241 , \41242 , \41243 , \41244 , \41245 , \41246 , \41247 , \41248 , \41249 , \41250 ,
         \41251 , \41252 , \41253 , \41254 , \41255 , \41256 , \41257 , \41258 , \41259 , \41260 ,
         \41261 , \41262 , \41263 , \41264 , \41265 , \41266 , \41267 , \41268 , \41269 , \41270 ,
         \41271 , \41272 , \41273 , \41274 , \41275 , \41276 , \41277 , \41278 , \41279 , \41280 ,
         \41281 , \41282 , \41283 , \41284 , \41285 , \41286 , \41287 , \41288 , \41289 , \41290 ,
         \41291 , \41292 , \41293 , \41294 , \41295 , \41296 , \41297 , \41298 , \41299 , \41300 ,
         \41301 , \41302 , \41303 , \41304 , \41305 , \41306 , \41307 , \41308 , \41309 , \41310 ,
         \41311 , \41312 , \41313 , \41314 , \41315 , \41316 , \41317 , \41318 , \41319 , \41320 ,
         \41321 , \41322 , \41323 , \41324 , \41325 , \41326 , \41327 , \41328 , \41329 , \41330 ,
         \41331 , \41332 , \41333 , \41334 , \41335 , \41336 , \41337 , \41338 , \41339 , \41340 ,
         \41341 , \41342 , \41343 , \41344 , \41345 , \41346 , \41347 , \41348 , \41349 , \41350 ,
         \41351 , \41352 , \41353 , \41354 , \41355 , \41356 , \41357 , \41358 , \41359 , \41360 ,
         \41361 , \41362 , \41363 , \41364 , \41365 , \41366 , \41367 , \41368 , \41369 , \41370 ,
         \41371 , \41372 , \41373 , \41374 , \41375 , \41376 , \41377 , \41378 , \41379 , \41380 ,
         \41381 , \41382 , \41383 , \41384 , \41385 , \41386 , \41387 , \41388 , \41389 , \41390 ,
         \41391 , \41392 , \41393 , \41394 , \41395 , \41396 , \41397 , \41398 , \41399 , \41400 ,
         \41401 , \41402 , \41403 , \41404 , \41405 , \41406 , \41407 , \41408 , \41409 , \41410 ,
         \41411 , \41412 , \41413 , \41414 , \41415 , \41416 , \41417 , \41418 , \41419 , \41420 ,
         \41421 , \41422 , \41423 , \41424 , \41425 , \41426 , \41427 , \41428 , \41429 , \41430 ,
         \41431 , \41432 , \41433 , \41434 , \41435 , \41436 , \41437 , \41438 , \41439 , \41440 ,
         \41441 , \41442 , \41443 , \41444 , \41445 , \41446 , \41447 , \41448 , \41449 , \41450 ,
         \41451 , \41452 , \41453 , \41454 , \41455 , \41456 , \41457 , \41458 , \41459 , \41460 ,
         \41461 , \41462 , \41463 , \41464 , \41465 , \41466 , \41467 , \41468 , \41469 , \41470 ,
         \41471 , \41472 , \41473 , \41474 , \41475 , \41476 , \41477 , \41478 , \41479 , \41480 ,
         \41481 , \41482 , \41483 , \41484 , \41485 , \41486 , \41487 , \41488 , \41489 , \41490 ,
         \41491 , \41492 , \41493 , \41494 , \41495 , \41496 , \41497 , \41498 , \41499 , \41500 ,
         \41501 , \41502 , \41503 , \41504 , \41505 , \41506 , \41507 , \41508 , \41509 , \41510 ,
         \41511 , \41512 , \41513 , \41514 , \41515 , \41516 , \41517 , \41518 , \41519 , \41520 ,
         \41521 , \41522 , \41523 , \41524 , \41525 , \41526 , \41527 , \41528 , \41529 , \41530 ,
         \41531 , \41532 , \41533 , \41534 , \41535 , \41536 , \41537 , \41538 , \41539 , \41540 ,
         \41541 , \41542 , \41543 , \41544 , \41545 , \41546 , \41547 , \41548 , \41549 , \41550 ,
         \41551 , \41552 , \41553 , \41554 , \41555 , \41556 , \41557 , \41558 , \41559 , \41560 ,
         \41561 , \41562 , \41563 , \41564 , \41565 , \41566 , \41567 , \41568 , \41569 , \41570 ,
         \41571 , \41572 , \41573 , \41574 , \41575 , \41576 , \41577 , \41578 , \41579 , \41580 ,
         \41581 , \41582 , \41583 , \41584 , \41585 , \41586 , \41587 , \41588 , \41589 , \41590 ,
         \41591 , \41592 , \41593 , \41594 , \41595 , \41596 , \41597 , \41598 , \41599 , \41600 ,
         \41601 , \41602 , \41603 , \41604 , \41605 , \41606 , \41607 , \41608 , \41609 , \41610 ,
         \41611 , \41612 , \41613 , \41614 , \41615 , \41616 , \41617 , \41618 , \41619 , \41620 ,
         \41621 , \41622 , \41623 , \41624 , \41625 , \41626 , \41627 , \41628 , \41629 , \41630 ,
         \41631 , \41632 , \41633 , \41634 , \41635 , \41636 , \41637 , \41638 , \41639 , \41640 ,
         \41641 , \41642 , \41643 , \41644 , \41645 , \41646 , \41647 , \41648 , \41649 , \41650 ,
         \41651 , \41652 , \41653 , \41654 , \41655 , \41656 , \41657 , \41658 , \41659 , \41660 ,
         \41661 , \41662 , \41663 , \41664 , \41665 , \41666 , \41667 , \41668 , \41669 , \41670 ,
         \41671 , \41672 , \41673 , \41674 , \41675 , \41676 , \41677 , \41678 , \41679 , \41680 ,
         \41681 , \41682 , \41683 , \41684 , \41685 , \41686 , \41687 , \41688 , \41689 , \41690 ,
         \41691 , \41692 , \41693 , \41694 , \41695 , \41696 , \41697 , \41698 , \41699 , \41700 ,
         \41701 , \41702 , \41703 , \41704 , \41705 , \41706 , \41707 , \41708 , \41709 , \41710 ,
         \41711 , \41712 , \41713 , \41714 , \41715 , \41716 , \41717 , \41718 , \41719 , \41720 ,
         \41721 , \41722 , \41723 , \41724 , \41725 , \41726 , \41727 , \41728 , \41729 , \41730 ,
         \41731 , \41732 , \41733 , \41734 , \41735 , \41736 , \41737 , \41738 , \41739 , \41740 ,
         \41741 , \41742 , \41743 , \41744 , \41745 , \41746 , \41747 , \41748 , \41749 , \41750 ,
         \41751 , \41752 , \41753 , \41754 , \41755 , \41756 , \41757 , \41758 , \41759 , \41760 ,
         \41761 , \41762 , \41763 , \41764 , \41765 , \41766 , \41767 , \41768 , \41769 , \41770 ,
         \41771 , \41772 , \41773 , \41774 , \41775 , \41776 , \41777 , \41778 , \41779 , \41780 ,
         \41781 , \41782 , \41783 , \41784 , \41785 , \41786 , \41787 , \41788 , \41789 , \41790 ,
         \41791 , \41792 , \41793 , \41794 , \41795 , \41796 , \41797 , \41798 , \41799 , \41800 ,
         \41801 , \41802 , \41803 , \41804 , \41805 , \41806 , \41807 , \41808 , \41809 , \41810 ,
         \41811 , \41812 , \41813 , \41814 , \41815 , \41816 , \41817 , \41818 , \41819 , \41820 ,
         \41821 , \41822 , \41823 , \41824 , \41825 , \41826 , \41827 , \41828 , \41829 , \41830 ,
         \41831 , \41832 , \41833 , \41834 , \41835 , \41836 , \41837 , \41838 , \41839 , \41840 ,
         \41841 , \41842 , \41843 , \41844 , \41845 , \41846 , \41847 , \41848 , \41849 , \41850 ,
         \41851 , \41852 , \41853 , \41854 , \41855 , \41856 , \41857 , \41858 , \41859 , \41860 ,
         \41861 , \41862 , \41863 , \41864 , \41865 , \41866 , \41867 , \41868 , \41869 , \41870 ,
         \41871 , \41872 , \41873 , \41874 , \41875 , \41876 , \41877 , \41878 , \41879 , \41880 ,
         \41881 , \41882 , \41883 , \41884 , \41885 , \41886 , \41887 , \41888 , \41889 , \41890 ,
         \41891 , \41892 , \41893 , \41894 , \41895 , \41896 , \41897 , \41898 , \41899 , \41900 ,
         \41901 , \41902 , \41903 , \41904 , \41905 , \41906 , \41907 , \41908 , \41909 , \41910 ,
         \41911 , \41912 , \41913 , \41914 , \41915 , \41916 , \41917 , \41918 , \41919 , \41920 ,
         \41921 , \41922 , \41923 , \41924 , \41925 , \41926 , \41927 , \41928 , \41929 , \41930 ,
         \41931 , \41932 , \41933 , \41934 , \41935 , \41936 , \41937 , \41938 , \41939 , \41940 ,
         \41941 , \41942 , \41943 , \41944 , \41945 , \41946 , \41947 , \41948 , \41949 , \41950 ,
         \41951 , \41952 , \41953 , \41954 , \41955 , \41956 , \41957 , \41958 , \41959 , \41960 ,
         \41961 , \41962 , \41963 , \41964 , \41965 , \41966 , \41967 , \41968 , \41969 , \41970 ,
         \41971 , \41972 , \41973 , \41974 , \41975 , \41976 , \41977 , \41978 , \41979 , \41980 ,
         \41981 , \41982 , \41983 , \41984 , \41985 , \41986 , \41987 , \41988 , \41989 , \41990 ,
         \41991 , \41992 , \41993 , \41994 , \41995 , \41996 , \41997 , \41998 , \41999 , \42000 ,
         \42001 , \42002 , \42003 , \42004 , \42005 , \42006 , \42007 , \42008 , \42009 , \42010 ,
         \42011 , \42012 , \42013 , \42014 , \42015 , \42016 , \42017 , \42018 , \42019 , \42020 ,
         \42021 , \42022 , \42023 , \42024 , \42025 , \42026 , \42027 , \42028 , \42029 , \42030 ,
         \42031 , \42032 , \42033 , \42034 , \42035 , \42036 , \42037 , \42038 , \42039 , \42040 ,
         \42041 , \42042 , \42043 , \42044 , \42045 , \42046 , \42047 , \42048 , \42049 , \42050 ,
         \42051 , \42052 , \42053 , \42054 , \42055 , \42056 , \42057 , \42058 , \42059 , \42060 ,
         \42061 , \42062 , \42063 , \42064 , \42065 , \42066 , \42067 , \42068 , \42069 , \42070 ,
         \42071 , \42072 , \42073 , \42074 , \42075 , \42076 , \42077 , \42078 , \42079 , \42080 ,
         \42081 , \42082 , \42083 , \42084 , \42085 , \42086 , \42087 , \42088 , \42089 , \42090 ,
         \42091 , \42092 , \42093 , \42094 , \42095 , \42096 , \42097 , \42098 , \42099 , \42100 ,
         \42101 , \42102 , \42103 , \42104 , \42105 , \42106 , \42107 , \42108 , \42109 , \42110 ,
         \42111 , \42112 , \42113 , \42114 , \42115 , \42116 , \42117 , \42118 , \42119 , \42120 ,
         \42121 , \42122 , \42123 , \42124 , \42125 , \42126 , \42127 , \42128 , \42129 , \42130 ,
         \42131 , \42132 , \42133 , \42134 , \42135 , \42136 , \42137 , \42138 , \42139 , \42140 ,
         \42141 , \42142 , \42143 , \42144 , \42145 , \42146 , \42147 , \42148 , \42149 , \42150 ,
         \42151 , \42152 , \42153 , \42154 , \42155 , \42156 , \42157 , \42158 , \42159 , \42160 ,
         \42161 , \42162 , \42163 , \42164 , \42165 , \42166 , \42167 , \42168 , \42169 , \42170 ,
         \42171 , \42172 , \42173 , \42174 , \42175 , \42176 , \42177 , \42178 , \42179 , \42180 ,
         \42181 , \42182 , \42183 , \42184 , \42185 , \42186 , \42187 , \42188 , \42189 , \42190 ,
         \42191 , \42192 , \42193 , \42194 , \42195 , \42196 , \42197 , \42198 , \42199 , \42200 ,
         \42201 , \42202 , \42203 , \42204 , \42205 , \42206 , \42207 , \42208 , \42209 , \42210 ,
         \42211 , \42212 , \42213 , \42214 , \42215 , \42216 , \42217 , \42218 , \42219 , \42220 ,
         \42221 , \42222 , \42223 , \42224 , \42225 , \42226 , \42227 , \42228 , \42229 , \42230 ,
         \42231 , \42232 , \42233 , \42234 , \42235 , \42236 , \42237 , \42238 , \42239 , \42240 ,
         \42241 , \42242 , \42243 , \42244 , \42245 , \42246 , \42247 , \42248 , \42249 , \42250 ,
         \42251 , \42252 , \42253 , \42254 , \42255 , \42256 , \42257 , \42258 , \42259 , \42260 ,
         \42261 , \42262 , \42263 , \42264 , \42265 , \42266 , \42267 , \42268 , \42269 , \42270 ,
         \42271 , \42272 , \42273 , \42274 , \42275 , \42276 , \42277 , \42278 , \42279 , \42280 ,
         \42281 , \42282 , \42283 , \42284 , \42285 , \42286 , \42287 , \42288 , \42289 , \42290 ,
         \42291 , \42292 , \42293 , \42294 , \42295 , \42296 , \42297 , \42298 , \42299 , \42300 ,
         \42301 , \42302 , \42303 , \42304 , \42305 , \42306 , \42307 , \42308 , \42309 , \42310 ,
         \42311 , \42312 , \42313 , \42314 , \42315 , \42316 , \42317 , \42318 , \42319 , \42320 ,
         \42321 , \42322 , \42323 , \42324 , \42325 , \42326 , \42327 , \42328 , \42329 , \42330 ,
         \42331 , \42332 , \42333 , \42334 , \42335 , \42336 , \42337 , \42338 , \42339 , \42340 ,
         \42341 , \42342 , \42343 , \42344 , \42345 , \42346 , \42347 , \42348 , \42349 , \42350 ,
         \42351 , \42352 , \42353 , \42354 , \42355 , \42356 , \42357 , \42358 , \42359 , \42360 ,
         \42361 , \42362 , \42363 , \42364 , \42365 , \42366 , \42367 , \42368 , \42369 , \42370 ,
         \42371 , \42372 , \42373 , \42374 , \42375 , \42376 , \42377 , \42378 , \42379 , \42380 ,
         \42381 , \42382 , \42383 , \42384 , \42385 , \42386 , \42387 , \42388 , \42389 , \42390 ,
         \42391 , \42392 , \42393 , \42394 , \42395 , \42396 , \42397 , \42398 , \42399 , \42400 ,
         \42401 , \42402 , \42403 , \42404 , \42405 , \42406 , \42407 , \42408 , \42409 , \42410 ,
         \42411 , \42412 , \42413 , \42414 , \42415 , \42416 , \42417 , \42418 , \42419 , \42420 ,
         \42421 , \42422 , \42423 , \42424 , \42425 , \42426 , \42427 , \42428 , \42429 , \42430 ,
         \42431 , \42432 , \42433 , \42434 , \42435 , \42436 , \42437 , \42438 , \42439 , \42440 ,
         \42441 , \42442 , \42443 , \42444 , \42445 , \42446 , \42447 , \42448 , \42449 , \42450 ,
         \42451 , \42452 , \42453 , \42454 , \42455 , \42456 , \42457 , \42458 , \42459 , \42460 ,
         \42461 , \42462 , \42463 , \42464 , \42465 , \42466 , \42467 , \42468 , \42469 , \42470 ,
         \42471 , \42472 , \42473 , \42474 , \42475 , \42476 , \42477 , \42478 , \42479 , \42480 ,
         \42481 , \42482 , \42483 , \42484 , \42485 , \42486 , \42487 , \42488 , \42489 , \42490 ,
         \42491 , \42492 , \42493 , \42494 , \42495 , \42496 , \42497 , \42498 , \42499 , \42500 ,
         \42501 , \42502 , \42503 , \42504 , \42505 , \42506 , \42507 , \42508 , \42509 , \42510 ,
         \42511 , \42512 , \42513 , \42514 , \42515 , \42516 , \42517 , \42518 , \42519 , \42520 ,
         \42521 , \42522 , \42523 , \42524 , \42525 , \42526 , \42527 , \42528 , \42529 , \42530 ,
         \42531 , \42532 , \42533 , \42534 , \42535 , \42536 , \42537 , \42538 , \42539 , \42540 ,
         \42541 , \42542 , \42543 , \42544 , \42545 , \42546 , \42547 , \42548 , \42549 , \42550 ,
         \42551 , \42552 , \42553 , \42554 , \42555 , \42556 , \42557 , \42558 , \42559 , \42560 ,
         \42561 , \42562 , \42563 , \42564 , \42565 , \42566 , \42567 , \42568 , \42569 , \42570 ,
         \42571 , \42572 , \42573 , \42574 , \42575 , \42576 , \42577 , \42578 , \42579 , \42580 ,
         \42581 , \42582 , \42583 , \42584 , \42585 , \42586 , \42587 , \42588 , \42589 , \42590 ,
         \42591 , \42592 , \42593 , \42594 , \42595 , \42596 , \42597 , \42598 , \42599 , \42600 ,
         \42601 , \42602 , \42603 , \42604 , \42605 , \42606 , \42607 , \42608 , \42609 , \42610 ,
         \42611 , \42612 , \42613 , \42614 , \42615 , \42616 , \42617 , \42618 , \42619 , \42620 ,
         \42621 , \42622 , \42623 , \42624 , \42625 , \42626 , \42627 , \42628 , \42629 , \42630 ,
         \42631 , \42632 , \42633 , \42634 , \42635 , \42636 , \42637 , \42638 , \42639 , \42640 ,
         \42641 , \42642 , \42643 , \42644 , \42645 , \42646 , \42647 , \42648 , \42649 , \42650 ,
         \42651 , \42652 , \42653 , \42654 , \42655 , \42656 , \42657 , \42658 , \42659 , \42660 ,
         \42661 , \42662 , \42663 , \42664 , \42665 , \42666 , \42667 , \42668 , \42669 , \42670 ,
         \42671 , \42672 , \42673 , \42674 , \42675 , \42676 , \42677 , \42678 , \42679 , \42680 ,
         \42681 , \42682 , \42683 , \42684 , \42685 , \42686 , \42687 , \42688 , \42689 , \42690 ,
         \42691 , \42692 , \42693 , \42694 , \42695 , \42696 , \42697 , \42698 , \42699 , \42700 ,
         \42701 , \42702 , \42703 , \42704 , \42705 , \42706 , \42707 , \42708 , \42709 , \42710 ,
         \42711 , \42712 , \42713 , \42714 , \42715 , \42716 , \42717 , \42718 , \42719 , \42720 ,
         \42721 , \42722 , \42723 , \42724 , \42725 , \42726 , \42727 , \42728 , \42729 , \42730 ,
         \42731 , \42732 , \42733 , \42734 , \42735 , \42736 , \42737 , \42738 , \42739 , \42740 ,
         \42741 , \42742 , \42743 , \42744 , \42745 , \42746 , \42747 , \42748 , \42749 , \42750 ,
         \42751 , \42752 , \42753 , \42754 , \42755 , \42756 , \42757 , \42758 , \42759 , \42760 ,
         \42761 , \42762 , \42763 , \42764 , \42765 , \42766 , \42767 , \42768 , \42769 , \42770 ,
         \42771 , \42772 , \42773 , \42774 , \42775 , \42776 , \42777 , \42778 , \42779 , \42780 ,
         \42781 , \42782 , \42783 , \42784 , \42785 , \42786 , \42787 , \42788 , \42789 , \42790 ,
         \42791 , \42792 , \42793 , \42794 , \42795 , \42796 , \42797 , \42798 , \42799 , \42800 ,
         \42801 , \42802 , \42803 , \42804 , \42805 , \42806 , \42807 , \42808 , \42809 , \42810 ,
         \42811 , \42812 , \42813 , \42814 , \42815 , \42816 , \42817 , \42818 , \42819 , \42820 ,
         \42821 , \42822 , \42823 , \42824 , \42825 , \42826 , \42827 , \42828 , \42829 , \42830 ,
         \42831 , \42832 , \42833 , \42834 , \42835 , \42836 , \42837 , \42838 , \42839 , \42840 ,
         \42841 , \42842 , \42843 , \42844 , \42845 , \42846 , \42847 , \42848 , \42849 , \42850 ,
         \42851 , \42852 , \42853 , \42854 , \42855 , \42856 , \42857 , \42858 , \42859 , \42860 ,
         \42861 , \42862 , \42863 , \42864 , \42865 , \42866 , \42867 , \42868 , \42869 , \42870 ,
         \42871 , \42872 , \42873 , \42874 , \42875 , \42876 , \42877 , \42878 , \42879 , \42880 ,
         \42881 , \42882 , \42883 , \42884 , \42885 , \42886 , \42887 , \42888 , \42889 , \42890 ,
         \42891 , \42892 , \42893 , \42894 , \42895 , \42896 , \42897 , \42898 , \42899 , \42900 ,
         \42901 , \42902 , \42903 , \42904 , \42905 , \42906 , \42907 , \42908 , \42909 , \42910 ,
         \42911 , \42912 , \42913 , \42914 , \42915 , \42916 , \42917 , \42918 , \42919 , \42920 ,
         \42921 , \42922 , \42923 , \42924 , \42925 , \42926 , \42927 , \42928 , \42929 , \42930 ,
         \42931 , \42932 , \42933 , \42934 , \42935 , \42936 , \42937 , \42938 , \42939 , \42940 ,
         \42941 , \42942 , \42943 , \42944 , \42945 , \42946 , \42947 , \42948 , \42949 , \42950 ,
         \42951 , \42952 , \42953 , \42954 , \42955 , \42956 , \42957 , \42958 , \42959 , \42960 ,
         \42961 , \42962 , \42963 , \42964 , \42965 , \42966 , \42967 , \42968 , \42969 , \42970 ,
         \42971 , \42972 , \42973 , \42974 , \42975 , \42976 , \42977 , \42978 , \42979 , \42980 ,
         \42981 , \42982 , \42983 , \42984 , \42985 , \42986 , \42987 , \42988 , \42989 , \42990 ,
         \42991 , \42992 , \42993 , \42994 , \42995 , \42996 , \42997 , \42998 , \42999 , \43000 ,
         \43001 , \43002 , \43003 , \43004 , \43005 , \43006 , \43007 , \43008 , \43009 , \43010 ,
         \43011 , \43012 , \43013 , \43014 , \43015 , \43016 , \43017 , \43018 , \43019 , \43020 ,
         \43021 , \43022 , \43023 , \43024 , \43025 , \43026 , \43027 , \43028 , \43029 , \43030 ,
         \43031 , \43032 , \43033 , \43034 , \43035 , \43036 , \43037 , \43038 , \43039 , \43040 ,
         \43041 , \43042 , \43043 , \43044 , \43045 , \43046 , \43047 , \43048 , \43049 , \43050 ,
         \43051 , \43052 , \43053 , \43054 , \43055 , \43056 , \43057 , \43058 , \43059 , \43060 ,
         \43061 , \43062 , \43063 , \43064 , \43065 , \43066 , \43067 , \43068 , \43069 , \43070 ,
         \43071 , \43072 , \43073 , \43074 , \43075 , \43076 , \43077 , \43078 , \43079 , \43080 ,
         \43081 , \43082 , \43083 , \43084 , \43085 , \43086 , \43087 , \43088 , \43089 , \43090 ,
         \43091 , \43092 , \43093 , \43094 , \43095 , \43096 , \43097 , \43098 , \43099 , \43100 ,
         \43101 , \43102 , \43103 , \43104 , \43105 , \43106 , \43107 , \43108 , \43109 , \43110 ,
         \43111 , \43112 , \43113 , \43114 , \43115 , \43116 , \43117 , \43118 , \43119 , \43120 ,
         \43121 , \43122 , \43123 , \43124 , \43125 , \43126 , \43127 , \43128 , \43129 , \43130 ,
         \43131 , \43132 , \43133 , \43134 , \43135 , \43136 , \43137 , \43138 , \43139 , \43140 ,
         \43141 , \43142 , \43143 , \43144 , \43145 , \43146 , \43147 , \43148 , \43149 , \43150 ,
         \43151 , \43152 , \43153 , \43154 , \43155 , \43156 , \43157 , \43158 , \43159 , \43160 ,
         \43161 , \43162 , \43163 , \43164 , \43165 , \43166 , \43167 , \43168 , \43169 , \43170 ,
         \43171 , \43172 , \43173 , \43174 , \43175 , \43176 , \43177 , \43178 , \43179 , \43180 ,
         \43181 , \43182 , \43183 , \43184 , \43185 , \43186 , \43187 , \43188 , \43189 , \43190 ,
         \43191 , \43192 , \43193 , \43194 , \43195 , \43196 , \43197 , \43198 , \43199 , \43200 ,
         \43201 , \43202 , \43203 , \43204 , \43205 , \43206 , \43207 , \43208 , \43209 , \43210 ,
         \43211 , \43212 , \43213 , \43214 , \43215 , \43216 , \43217 , \43218 , \43219 , \43220 ,
         \43221 , \43222 , \43223 , \43224 , \43225 , \43226 , \43227 , \43228 , \43229 , \43230 ,
         \43231 , \43232 , \43233 , \43234 , \43235 , \43236 , \43237 , \43238 , \43239 , \43240 ,
         \43241 , \43242 , \43243 , \43244 , \43245 , \43246 , \43247 , \43248 , \43249 , \43250 ,
         \43251 , \43252 , \43253 , \43254 , \43255 , \43256 , \43257 , \43258 , \43259 , \43260 ,
         \43261 , \43262 , \43263 , \43264 , \43265 , \43266 , \43267 , \43268 , \43269 , \43270 ,
         \43271 , \43272 , \43273 , \43274 , \43275 , \43276 , \43277 , \43278 , \43279 , \43280 ,
         \43281 , \43282 , \43283 , \43284 , \43285 , \43286 , \43287 , \43288 , \43289 , \43290 ,
         \43291 , \43292 , \43293 , \43294 , \43295 , \43296 , \43297 , \43298 , \43299 , \43300 ,
         \43301 , \43302 , \43303 , \43304 , \43305 , \43306 , \43307 , \43308 , \43309 , \43310 ,
         \43311 , \43312 , \43313 , \43314 , \43315 , \43316 , \43317 , \43318 , \43319 , \43320 ,
         \43321 , \43322 , \43323 , \43324 , \43325 , \43326 , \43327 , \43328 , \43329 , \43330 ,
         \43331 , \43332 , \43333 , \43334 , \43335 , \43336 , \43337 , \43338 , \43339 , \43340 ,
         \43341 , \43342 , \43343 , \43344 , \43345 , \43346 , \43347 , \43348 , \43349 , \43350 ,
         \43351 , \43352 , \43353 , \43354 , \43355 , \43356 , \43357 , \43358 , \43359 , \43360 ,
         \43361 , \43362 , \43363 , \43364 , \43365 , \43366 , \43367 , \43368 , \43369 , \43370 ,
         \43371 , \43372 , \43373 , \43374 , \43375 , \43376 , \43377 , \43378 , \43379 , \43380 ,
         \43381 , \43382 , \43383 , \43384 , \43385 , \43386 , \43387 , \43388 , \43389 , \43390 ,
         \43391 , \43392 , \43393 , \43394 , \43395 , \43396 , \43397 , \43398 , \43399 , \43400 ,
         \43401 , \43402 , \43403 , \43404 , \43405 , \43406 , \43407 , \43408 , \43409 , \43410 ,
         \43411 , \43412 , \43413 , \43414 , \43415 , \43416 , \43417 , \43418 , \43419 , \43420 ,
         \43421 , \43422 , \43423 , \43424 , \43425 , \43426 , \43427 , \43428 , \43429 , \43430 ,
         \43431 , \43432 , \43433 , \43434 , \43435 , \43436 , \43437 , \43438 , \43439 , \43440 ,
         \43441 , \43442 , \43443 , \43444 , \43445 , \43446 , \43447 , \43448 , \43449 , \43450 ,
         \43451 , \43452 , \43453 , \43454 , \43455 , \43456 , \43457 , \43458 , \43459 , \43460 ,
         \43461 , \43462 , \43463 , \43464 , \43465 , \43466 , \43467 , \43468 , \43469 , \43470 ,
         \43471 , \43472 , \43473 , \43474 , \43475 , \43476 , \43477 , \43478 , \43479 , \43480 ,
         \43481 , \43482 , \43483 , \43484 , \43485 , \43486 , \43487 , \43488 , \43489 , \43490 ,
         \43491 , \43492 , \43493 , \43494 , \43495 , \43496 , \43497 , \43498 , \43499 , \43500 ,
         \43501 , \43502 , \43503 , \43504 , \43505 , \43506 , \43507 , \43508 , \43509 , \43510 ,
         \43511 , \43512 , \43513 , \43514 , \43515 , \43516 , \43517 , \43518 , \43519 , \43520 ,
         \43521 , \43522 , \43523 , \43524 , \43525 , \43526 , \43527 , \43528 , \43529 , \43530 ,
         \43531 , \43532 , \43533 , \43534 , \43535 , \43536 , \43537 , \43538 , \43539 , \43540 ,
         \43541 , \43542 , \43543 , \43544 , \43545 , \43546 , \43547 , \43548 , \43549 , \43550 ,
         \43551 , \43552 , \43553 , \43554 , \43555 , \43556 , \43557 , \43558 , \43559 , \43560 ,
         \43561 , \43562 , \43563 , \43564 , \43565 , \43566 , \43567 , \43568 , \43569 , \43570 ,
         \43571 , \43572 , \43573 , \43574 , \43575 , \43576 , \43577 , \43578 , \43579 , \43580 ,
         \43581 , \43582 , \43583 , \43584 , \43585 , \43586 , \43587 , \43588 , \43589 , \43590 ,
         \43591 , \43592 , \43593 , \43594 , \43595 , \43596 , \43597 , \43598 , \43599 , \43600 ,
         \43601 , \43602 , \43603 , \43604 , \43605 , \43606 , \43607 , \43608 , \43609 , \43610 ,
         \43611 , \43612 , \43613 , \43614 , \43615 , \43616 , \43617 , \43618 , \43619 , \43620 ,
         \43621 , \43622 , \43623 , \43624 , \43625 , \43626 , \43627 , \43628 , \43629 , \43630 ,
         \43631 , \43632 , \43633 , \43634 , \43635 , \43636 , \43637 , \43638 , \43639 , \43640 ,
         \43641 , \43642 , \43643 , \43644 , \43645 , \43646 , \43647 , \43648 , \43649 , \43650 ,
         \43651 , \43652 , \43653 , \43654 , \43655 , \43656 , \43657 , \43658 , \43659 , \43660 ,
         \43661 , \43662 , \43663 , \43664 , \43665 , \43666 , \43667 , \43668 , \43669 , \43670 ,
         \43671 , \43672 , \43673 , \43674 , \43675 , \43676 , \43677 , \43678 , \43679 , \43680 ,
         \43681 , \43682 , \43683 , \43684 , \43685 , \43686 , \43687 , \43688 , \43689 , \43690 ,
         \43691 , \43692 , \43693 , \43694 , \43695 , \43696 , \43697 , \43698 , \43699 , \43700 ,
         \43701 , \43702 , \43703 , \43704 , \43705 , \43706 , \43707 , \43708 , \43709 , \43710 ,
         \43711 , \43712 , \43713 , \43714 , \43715 , \43716 , \43717 , \43718 , \43719 , \43720 ,
         \43721 , \43722 , \43723 , \43724 , \43725 , \43726 , \43727 , \43728 , \43729 , \43730 ,
         \43731 , \43732 , \43733 , \43734 , \43735 , \43736 , \43737 , \43738 , \43739 , \43740 ,
         \43741 , \43742 , \43743 , \43744 , \43745 , \43746 , \43747 , \43748 , \43749 , \43750 ,
         \43751 , \43752 , \43753 , \43754 , \43755 , \43756 , \43757 , \43758 , \43759 , \43760 ,
         \43761 , \43762 , \43763 , \43764 , \43765 , \43766 , \43767 , \43768 , \43769 , \43770 ,
         \43771 , \43772 , \43773 , \43774 , \43775 , \43776 , \43777 , \43778 , \43779 , \43780 ,
         \43781 , \43782 , \43783 , \43784 , \43785 , \43786 , \43787 , \43788 , \43789 , \43790 ,
         \43791 , \43792 , \43793 , \43794 , \43795 , \43796 , \43797 , \43798 , \43799 , \43800 ,
         \43801 , \43802 , \43803 , \43804 , \43805 , \43806 , \43807 , \43808 , \43809 , \43810 ,
         \43811 , \43812 , \43813 , \43814 , \43815 , \43816 , \43817 , \43818 , \43819 , \43820 ,
         \43821 , \43822 , \43823 , \43824 , \43825 , \43826 , \43827 , \43828 , \43829 , \43830 ,
         \43831 , \43832 , \43833 , \43834 , \43835 , \43836 , \43837 , \43838 , \43839 , \43840 ,
         \43841 , \43842 , \43843 , \43844 , \43845 , \43846 , \43847 , \43848 , \43849 , \43850 ,
         \43851 , \43852 , \43853 , \43854 , \43855 , \43856 , \43857 , \43858 , \43859 , \43860 ,
         \43861 , \43862 , \43863 , \43864 , \43865 , \43866 , \43867 , \43868 , \43869 , \43870 ,
         \43871 , \43872 , \43873 , \43874 , \43875 , \43876 , \43877 , \43878 , \43879 , \43880 ,
         \43881 , \43882 , \43883 , \43884 , \43885 , \43886 , \43887 , \43888 , \43889 , \43890 ,
         \43891 , \43892 , \43893 , \43894 , \43895 , \43896 , \43897 , \43898 , \43899 , \43900 ,
         \43901 , \43902 , \43903 , \43904 , \43905 , \43906 , \43907 , \43908 , \43909 , \43910 ,
         \43911 , \43912 , \43913 , \43914 , \43915 , \43916 , \43917 , \43918 , \43919 , \43920 ,
         \43921 , \43922 , \43923 , \43924 , \43925 , \43926 , \43927 , \43928 , \43929 , \43930 ,
         \43931 , \43932 , \43933 , \43934 , \43935 , \43936 , \43937 , \43938 , \43939 , \43940 ,
         \43941 , \43942 , \43943 , \43944 , \43945 , \43946 , \43947 , \43948 , \43949 , \43950 ,
         \43951 , \43952 , \43953 , \43954 , \43955 , \43956 , \43957 , \43958 , \43959 , \43960 ,
         \43961 , \43962 , \43963 , \43964 , \43965 , \43966 , \43967 , \43968 , \43969 , \43970 ,
         \43971 , \43972 , \43973 , \43974 , \43975 , \43976 , \43977 , \43978 , \43979 , \43980 ,
         \43981 , \43982 , \43983 , \43984 , \43985 , \43986 , \43987 , \43988 , \43989 , \43990 ,
         \43991 , \43992 , \43993 , \43994 , \43995 , \43996 , \43997 , \43998 , \43999 , \44000 ,
         \44001 , \44002 , \44003 , \44004 , \44005 , \44006 , \44007 , \44008 , \44009 , \44010 ,
         \44011 , \44012 , \44013 , \44014 , \44015 , \44016 , \44017 , \44018 , \44019 , \44020 ,
         \44021 , \44022 , \44023 , \44024 , \44025 , \44026 , \44027 , \44028 , \44029 , \44030 ,
         \44031 , \44032 , \44033 , \44034 , \44035 , \44036 , \44037 , \44038 , \44039 , \44040 ,
         \44041 , \44042 , \44043 , \44044 , \44045 , \44046 , \44047 , \44048 , \44049 , \44050 ,
         \44051 , \44052 , \44053 , \44054 , \44055 , \44056 , \44057 , \44058 , \44059 , \44060 ,
         \44061 , \44062 , \44063 , \44064 , \44065 , \44066 , \44067 , \44068 , \44069 , \44070 ,
         \44071 , \44072 , \44073 , \44074 , \44075 , \44076 , \44077 , \44078 , \44079 , \44080 ,
         \44081 , \44082 , \44083 , \44084 , \44085 , \44086 , \44087 , \44088 , \44089 , \44090 ,
         \44091 , \44092 , \44093 , \44094 , \44095 , \44096 , \44097 , \44098 , \44099 , \44100 ,
         \44101 , \44102 , \44103 , \44104 , \44105 , \44106 , \44107 , \44108 , \44109 , \44110 ,
         \44111 , \44112 , \44113 , \44114 , \44115 , \44116 , \44117 , \44118 , \44119 , \44120 ,
         \44121 , \44122 , \44123 , \44124 , \44125 , \44126 , \44127 , \44128 , \44129 , \44130 ,
         \44131 , \44132 , \44133 , \44134 , \44135 , \44136 , \44137 , \44138 , \44139 , \44140 ,
         \44141 , \44142 , \44143 , \44144 , \44145 , \44146 , \44147 , \44148 , \44149 , \44150 ,
         \44151 , \44152 , \44153 , \44154 , \44155 , \44156 , \44157 , \44158 , \44159 , \44160 ,
         \44161 , \44162 , \44163 , \44164 , \44165 , \44166 , \44167 , \44168 , \44169 , \44170 ,
         \44171 , \44172 , \44173 , \44174 , \44175 , \44176 , \44177 , \44178 , \44179 , \44180 ,
         \44181 , \44182 , \44183 , \44184 , \44185 , \44186 , \44187 , \44188 , \44189 , \44190 ,
         \44191 , \44192 , \44193 , \44194 , \44195 , \44196 , \44197 , \44198 , \44199 , \44200 ,
         \44201 , \44202 , \44203 , \44204 , \44205 , \44206 , \44207 , \44208 , \44209 , \44210 ,
         \44211 , \44212 , \44213 , \44214 , \44215 , \44216 , \44217 , \44218 , \44219 , \44220 ,
         \44221 , \44222 , \44223 , \44224 , \44225 , \44226 , \44227 , \44228 , \44229 , \44230 ,
         \44231 , \44232 , \44233 , \44234 , \44235 , \44236 , \44237 , \44238 , \44239 , \44240 ,
         \44241 , \44242 , \44243 , \44244 , \44245 , \44246 , \44247 , \44248 , \44249 , \44250 ,
         \44251 , \44252 , \44253 , \44254 , \44255 , \44256 , \44257 , \44258 , \44259 , \44260 ,
         \44261 , \44262 , \44263 , \44264 , \44265 , \44266 , \44267 , \44268 , \44269 , \44270 ,
         \44271 , \44272 , \44273 , \44274 , \44275 , \44276 , \44277 , \44278 , \44279 , \44280 ,
         \44281 , \44282 , \44283 , \44284 , \44285 , \44286 , \44287 , \44288 , \44289 , \44290 ,
         \44291 , \44292 , \44293 , \44294 , \44295 , \44296 , \44297 , \44298 , \44299 , \44300 ,
         \44301 , \44302 , \44303 , \44304 , \44305 , \44306 , \44307 , \44308 , \44309 , \44310 ,
         \44311 , \44312 , \44313 , \44314 , \44315 , \44316 , \44317 , \44318 , \44319 , \44320 ,
         \44321 , \44322 , \44323 , \44324 , \44325 , \44326 , \44327 , \44328 , \44329 , \44330 ,
         \44331 , \44332 , \44333 , \44334 , \44335 , \44336 , \44337 , \44338 , \44339 , \44340 ,
         \44341 , \44342 , \44343 , \44344 , \44345 , \44346 , \44347 , \44348 , \44349 , \44350 ,
         \44351 , \44352 , \44353 , \44354 , \44355 , \44356 , \44357 , \44358 , \44359 , \44360 ,
         \44361 , \44362 , \44363 , \44364 , \44365 , \44366 , \44367 , \44368 , \44369 , \44370 ,
         \44371 , \44372 , \44373 , \44374 , \44375 , \44376 , \44377 , \44378 , \44379 , \44380 ,
         \44381 , \44382 , \44383 , \44384 , \44385 , \44386 , \44387 , \44388 , \44389 , \44390 ,
         \44391 , \44392 , \44393 , \44394 , \44395 , \44396 , \44397 , \44398 , \44399 , \44400 ,
         \44401 , \44402 , \44403 , \44404 , \44405 , \44406 , \44407 , \44408 , \44409 , \44410 ,
         \44411 , \44412 , \44413 , \44414 , \44415 , \44416 , \44417 , \44418 , \44419 , \44420 ,
         \44421 , \44422 , \44423 , \44424 , \44425 , \44426 , \44427 , \44428 , \44429 , \44430 ,
         \44431 , \44432 , \44433 , \44434 , \44435 , \44436 , \44437 , \44438 , \44439 , \44440 ,
         \44441 , \44442 , \44443 , \44444 , \44445 , \44446 , \44447 , \44448 , \44449 , \44450 ,
         \44451 , \44452 , \44453 , \44454 , \44455 , \44456 , \44457 , \44458 , \44459 , \44460 ,
         \44461 , \44462 , \44463 , \44464 , \44465 , \44466 , \44467 , \44468 , \44469 , \44470 ,
         \44471 , \44472 , \44473 , \44474 , \44475 , \44476 , \44477 , \44478 , \44479 , \44480 ,
         \44481 , \44482 , \44483 , \44484 , \44485 , \44486 , \44487 , \44488 , \44489 , \44490 ,
         \44491 , \44492 , \44493 , \44494 , \44495 , \44496 , \44497 , \44498 , \44499 , \44500 ,
         \44501 , \44502 , \44503 , \44504 , \44505 , \44506 , \44507 , \44508 , \44509 , \44510 ,
         \44511 , \44512 , \44513 , \44514 , \44515 , \44516 , \44517 , \44518 , \44519 , \44520 ,
         \44521 , \44522 , \44523 , \44524 , \44525 , \44526 , \44527 , \44528 , \44529 , \44530 ,
         \44531 , \44532 , \44533 , \44534 , \44535 , \44536 , \44537 , \44538 , \44539 , \44540 ,
         \44541 , \44542 , \44543 , \44544 , \44545 , \44546 , \44547 , \44548 , \44549 , \44550 ,
         \44551 , \44552 , \44553 , \44554 , \44555 , \44556 , \44557 , \44558 , \44559 , \44560 ,
         \44561 , \44562 , \44563 , \44564 , \44565 , \44566 , \44567 , \44568 , \44569 , \44570 ,
         \44571 , \44572 , \44573 , \44574 , \44575 , \44576 , \44577 , \44578 , \44579 , \44580 ,
         \44581 , \44582 , \44583 , \44584 , \44585 , \44586 , \44587 , \44588 , \44589 , \44590 ,
         \44591 , \44592 , \44593 , \44594 , \44595 , \44596 , \44597 , \44598 , \44599 , \44600 ,
         \44601 , \44602 , \44603 , \44604 , \44605 , \44606 , \44607 , \44608 , \44609 , \44610 ,
         \44611 , \44612 , \44613 , \44614 , \44615 , \44616 , \44617 , \44618 , \44619 , \44620 ,
         \44621 , \44622 , \44623 , \44624 , \44625 , \44626 , \44627 , \44628 , \44629 , \44630 ,
         \44631 , \44632 , \44633 , \44634 , \44635 , \44636 , \44637 , \44638 , \44639 , \44640 ,
         \44641 , \44642 , \44643 , \44644 , \44645 , \44646 , \44647 , \44648 , \44649 , \44650 ,
         \44651 , \44652 , \44653 , \44654 , \44655 , \44656 , \44657 , \44658 , \44659 , \44660 ,
         \44661 , \44662 , \44663 , \44664 , \44665 , \44666 , \44667 , \44668 , \44669 , \44670 ,
         \44671 , \44672 , \44673 , \44674 , \44675 , \44676 , \44677 , \44678 , \44679 , \44680 ,
         \44681 , \44682 , \44683 , \44684 , \44685 , \44686 , \44687 , \44688 , \44689 , \44690 ,
         \44691 , \44692 , \44693 , \44694 , \44695 , \44696 , \44697 , \44698 , \44699 , \44700 ,
         \44701 , \44702 , \44703 , \44704 , \44705 , \44706 , \44707 , \44708 , \44709 , \44710 ,
         \44711 , \44712 , \44713 , \44714 , \44715 , \44716 , \44717 , \44718 , \44719 , \44720 ,
         \44721 , \44722 , \44723 , \44724 , \44725 , \44726 , \44727 , \44728 , \44729 , \44730 ,
         \44731 , \44732 , \44733 , \44734 , \44735 , \44736 , \44737 , \44738 , \44739 , \44740 ,
         \44741 , \44742 , \44743 , \44744 , \44745 , \44746 , \44747 , \44748 , \44749 , \44750 ,
         \44751 , \44752 , \44753 , \44754 , \44755 , \44756 , \44757 , \44758 , \44759 , \44760 ,
         \44761 , \44762 , \44763 , \44764 , \44765 , \44766 , \44767 , \44768 , \44769 , \44770 ,
         \44771 , \44772 , \44773 , \44774 , \44775 , \44776 , \44777 , \44778 , \44779 , \44780 ,
         \44781 , \44782 , \44783 , \44784 , \44785 , \44786 , \44787 , \44788 , \44789 , \44790 ,
         \44791 , \44792 , \44793 , \44794 , \44795 , \44796 , \44797 , \44798 , \44799 , \44800 ,
         \44801 , \44802 , \44803 , \44804 , \44805 , \44806 , \44807 , \44808 , \44809 , \44810 ,
         \44811 , \44812 , \44813 , \44814 , \44815 , \44816 , \44817 , \44818 , \44819 , \44820 ,
         \44821 , \44822 , \44823 , \44824 , \44825 , \44826 , \44827 , \44828 , \44829 , \44830 ,
         \44831 , \44832 , \44833 , \44834 , \44835 , \44836 , \44837 , \44838 , \44839 , \44840 ,
         \44841 , \44842 , \44843 , \44844 , \44845 , \44846 , \44847 , \44848 , \44849 , \44850 ,
         \44851 , \44852 , \44853 , \44854 , \44855 , \44856 , \44857 , \44858 , \44859 , \44860 ,
         \44861 , \44862 , \44863 , \44864 , \44865 , \44866 , \44867 , \44868 , \44869 , \44870 ,
         \44871 , \44872 , \44873 , \44874 , \44875 , \44876 , \44877 , \44878 , \44879 , \44880 ,
         \44881 , \44882 , \44883 , \44884 , \44885 , \44886 , \44887 , \44888 , \44889 , \44890 ,
         \44891 , \44892 , \44893 , \44894 , \44895 , \44896 , \44897 , \44898 , \44899 , \44900 ,
         \44901 , \44902 , \44903 , \44904 , \44905 , \44906 , \44907 , \44908 , \44909 , \44910 ,
         \44911 , \44912 , \44913 , \44914 , \44915 , \44916 , \44917 , \44918 , \44919 , \44920 ,
         \44921 , \44922 , \44923 , \44924 , \44925 , \44926 , \44927 , \44928 , \44929 , \44930 ,
         \44931 , \44932 , \44933 , \44934 , \44935 , \44936 , \44937 , \44938 , \44939 , \44940 ,
         \44941 , \44942 , \44943 , \44944 , \44945 , \44946 , \44947 , \44948 , \44949 , \44950 ,
         \44951 , \44952 , \44953 , \44954 , \44955 , \44956 , \44957 , \44958 , \44959 , \44960 ,
         \44961 , \44962 , \44963 , \44964 , \44965 , \44966 , \44967 , \44968 , \44969 , \44970 ,
         \44971 , \44972 , \44973 , \44974 , \44975 , \44976 , \44977 , \44978 , \44979 , \44980 ,
         \44981 , \44982 , \44983 , \44984 , \44985 , \44986 , \44987 , \44988 , \44989 , \44990 ,
         \44991 , \44992 , \44993 , \44994 , \44995 , \44996 , \44997 , \44998 , \44999 , \45000 ,
         \45001 , \45002 , \45003 , \45004 , \45005 , \45006 , \45007 , \45008 , \45009 , \45010 ,
         \45011 , \45012 , \45013 , \45014 , \45015 , \45016 , \45017 , \45018 , \45019 , \45020 ,
         \45021 , \45022 , \45023 , \45024 , \45025 , \45026 , \45027 , \45028 , \45029 , \45030 ,
         \45031 , \45032 , \45033 , \45034 , \45035 , \45036 , \45037 , \45038 , \45039 , \45040 ,
         \45041 , \45042 , \45043 , \45044 , \45045 , \45046 , \45047 , \45048 , \45049 , \45050 ,
         \45051 , \45052 , \45053 , \45054 , \45055 , \45056 , \45057 , \45058 , \45059 , \45060 ,
         \45061 , \45062 , \45063 , \45064 , \45065 , \45066 , \45067 , \45068 , \45069 , \45070 ,
         \45071 , \45072 , \45073 , \45074 , \45075 , \45076 , \45077 , \45078 , \45079 , \45080 ,
         \45081 , \45082 , \45083 , \45084 , \45085 , \45086 , \45087 , \45088 , \45089 , \45090 ,
         \45091 , \45092 , \45093 , \45094 , \45095 , \45096 , \45097 , \45098 , \45099 , \45100 ,
         \45101 , \45102 , \45103 , \45104 , \45105 , \45106 , \45107 , \45108 , \45109 , \45110 ,
         \45111 , \45112 , \45113 , \45114 , \45115 , \45116 , \45117 , \45118 , \45119 , \45120 ,
         \45121 , \45122 , \45123 , \45124 , \45125 , \45126 , \45127 , \45128 , \45129 , \45130 ,
         \45131 , \45132 , \45133 , \45134 , \45135 , \45136 , \45137 , \45138 , \45139 , \45140 ,
         \45141 , \45142 , \45143 , \45144 , \45145 , \45146 , \45147 , \45148 , \45149 , \45150 ,
         \45151 , \45152 , \45153 , \45154 , \45155 , \45156 , \45157 , \45158 , \45159 , \45160 ,
         \45161 , \45162 , \45163 , \45164 , \45165 , \45166 , \45167 , \45168 , \45169 , \45170 ,
         \45171 , \45172 , \45173 , \45174 , \45175 , \45176 , \45177 , \45178 , \45179 , \45180 ,
         \45181 , \45182 , \45183 , \45184 , \45185 , \45186 , \45187 , \45188 , \45189 , \45190 ,
         \45191 , \45192 , \45193 , \45194 , \45195 , \45196 , \45197 , \45198 , \45199 , \45200 ,
         \45201 , \45202 , \45203 , \45204 , \45205 , \45206 , \45207 , \45208 , \45209 , \45210 ,
         \45211 , \45212 , \45213 , \45214 , \45215 , \45216 , \45217 , \45218 , \45219 , \45220 ,
         \45221 , \45222 , \45223 , \45224 , \45225 , \45226 , \45227 , \45228 , \45229 , \45230 ,
         \45231 , \45232 , \45233 , \45234 , \45235 , \45236 , \45237 , \45238 , \45239 , \45240 ,
         \45241 , \45242 , \45243 , \45244 , \45245 , \45246 , \45247 , \45248 , \45249 , \45250 ,
         \45251 , \45252 , \45253 , \45254 , \45255 , \45256 , \45257 , \45258 , \45259 , \45260 ,
         \45261 , \45262 , \45263 , \45264 , \45265 , \45266 , \45267 , \45268 , \45269 , \45270 ,
         \45271 , \45272 , \45273 , \45274 , \45275 , \45276 , \45277 , \45278 , \45279 , \45280 ,
         \45281 , \45282 , \45283 , \45284 , \45285 , \45286 , \45287 , \45288 , \45289 , \45290 ,
         \45291 , \45292 , \45293 , \45294 , \45295 , \45296 , \45297 , \45298 , \45299 , \45300 ,
         \45301 , \45302 , \45303 , \45304 , \45305 , \45306 , \45307 , \45308 , \45309 , \45310 ,
         \45311 , \45312 , \45313 , \45314 , \45315 , \45316 , \45317 , \45318 , \45319 , \45320 ,
         \45321 , \45322 , \45323 , \45324 , \45325 , \45326 , \45327 , \45328 , \45329 , \45330 ,
         \45331 , \45332 , \45333 , \45334 , \45335 , \45336 , \45337 , \45338 , \45339 , \45340 ,
         \45341 , \45342 , \45343 , \45344 , \45345 , \45346 , \45347 , \45348 , \45349 , \45350 ,
         \45351 , \45352 , \45353 , \45354 , \45355 , \45356 , \45357 , \45358 , \45359 , \45360 ,
         \45361 , \45362 , \45363 , \45364 , \45365 , \45366 , \45367 , \45368 , \45369 , \45370 ,
         \45371 , \45372 , \45373 , \45374 , \45375 , \45376 , \45377 , \45378 , \45379 , \45380 ,
         \45381 , \45382 , \45383 , \45384 , \45385 , \45386 , \45387 , \45388 , \45389 , \45390 ,
         \45391 , \45392 , \45393 , \45394 , \45395 , \45396 , \45397 , \45398 , \45399 , \45400 ,
         \45401 , \45402 , \45403 , \45404 , \45405 , \45406 , \45407 , \45408 , \45409 , \45410 ,
         \45411 , \45412 , \45413 , \45414 , \45415 , \45416 , \45417 , \45418 , \45419 , \45420 ,
         \45421 , \45422 , \45423 , \45424 , \45425 , \45426 , \45427 , \45428 , \45429 , \45430 ,
         \45431 , \45432 , \45433 , \45434 , \45435 , \45436 , \45437 , \45438 , \45439 , \45440 ,
         \45441 , \45442 , \45443 , \45444 , \45445 , \45446 , \45447 , \45448 , \45449 , \45450 ,
         \45451 , \45452 , \45453 , \45454 , \45455 , \45456 , \45457 , \45458 , \45459 , \45460 ,
         \45461 , \45462 , \45463 , \45464 , \45465 , \45466 , \45467 , \45468 , \45469 , \45470 ,
         \45471 , \45472 , \45473 , \45474 , \45475 , \45476 , \45477 , \45478 , \45479 , \45480 ,
         \45481 , \45482 , \45483 , \45484 , \45485 , \45486 , \45487 , \45488 , \45489 , \45490 ,
         \45491 , \45492 , \45493 , \45494 , \45495 , \45496 , \45497 , \45498 , \45499 , \45500 ,
         \45501 , \45502 , \45503 , \45504 , \45505 , \45506 , \45507 , \45508 , \45509 , \45510 ,
         \45511 , \45512 , \45513 , \45514 , \45515 , \45516 , \45517 , \45518 , \45519 , \45520 ,
         \45521 , \45522 , \45523 , \45524 , \45525 , \45526 , \45527 , \45528 , \45529 , \45530 ,
         \45531 , \45532 , \45533 , \45534 , \45535 , \45536 , \45537 , \45538 , \45539 , \45540 ,
         \45541 , \45542 , \45543 , \45544 , \45545 , \45546 , \45547 , \45548 , \45549 , \45550 ,
         \45551 , \45552 , \45553 , \45554 , \45555 , \45556 , \45557 , \45558 , \45559 , \45560 ,
         \45561 , \45562 , \45563 , \45564 , \45565 , \45566 , \45567 , \45568 , \45569 , \45570 ,
         \45571 , \45572 , \45573 , \45574 , \45575 , \45576 , \45577 , \45578 , \45579 , \45580 ,
         \45581 , \45582 , \45583 , \45584 , \45585 , \45586 , \45587 , \45588 , \45589 , \45590 ,
         \45591 , \45592 , \45593 , \45594 , \45595 , \45596 , \45597 , \45598 , \45599 , \45600 ,
         \45601 , \45602 , \45603 , \45604 , \45605 , \45606 , \45607 , \45608 , \45609 , \45610 ,
         \45611 , \45612 , \45613 , \45614 , \45615 , \45616 , \45617 , \45618 , \45619 , \45620 ,
         \45621 , \45622 , \45623 , \45624 , \45625 , \45626 , \45627 , \45628 , \45629 , \45630 ,
         \45631 , \45632 , \45633 , \45634 , \45635 , \45636 , \45637 , \45638 , \45639 , \45640 ,
         \45641 , \45642 , \45643 , \45644 , \45645 , \45646 , \45647 , \45648 , \45649 , \45650 ,
         \45651 , \45652 , \45653 , \45654 , \45655 , \45656 , \45657 , \45658 , \45659 , \45660 ,
         \45661 , \45662 , \45663 , \45664 , \45665 , \45666 , \45667 , \45668 , \45669 , \45670 ,
         \45671 , \45672 , \45673 , \45674 , \45675 , \45676 , \45677 , \45678 , \45679 , \45680 ,
         \45681 , \45682 , \45683 , \45684 , \45685 , \45686 , \45687 , \45688 , \45689 , \45690 ,
         \45691 , \45692 , \45693 , \45694 , \45695 , \45696 , \45697 , \45698 , \45699 , \45700 ,
         \45701 , \45702 , \45703 , \45704 , \45705 , \45706 , \45707 , \45708 , \45709 , \45710 ,
         \45711 , \45712 , \45713 , \45714 , \45715 , \45716 , \45717 , \45718 , \45719 , \45720 ,
         \45721 , \45722 , \45723 , \45724 , \45725 , \45726 , \45727 , \45728 , \45729 , \45730 ,
         \45731 , \45732 , \45733 , \45734 , \45735 , \45736 , \45737 , \45738 , \45739 , \45740 ,
         \45741 , \45742 , \45743 , \45744 , \45745 , \45746 , \45747 , \45748 , \45749 , \45750 ,
         \45751 , \45752 , \45753 , \45754 , \45755 , \45756 , \45757 , \45758 , \45759 , \45760 ,
         \45761 , \45762 , \45763 , \45764 , \45765 , \45766 , \45767 , \45768 , \45769 , \45770 ,
         \45771 , \45772 , \45773 , \45774 , \45775 , \45776 , \45777 , \45778 , \45779 , \45780 ,
         \45781 , \45782 , \45783 , \45784 , \45785 , \45786 , \45787 , \45788 , \45789 , \45790 ,
         \45791 , \45792 , \45793 , \45794 , \45795 , \45796 , \45797 , \45798 , \45799 , \45800 ,
         \45801 , \45802 , \45803 , \45804 , \45805 , \45806 , \45807 , \45808 , \45809 , \45810 ,
         \45811 , \45812 , \45813 , \45814 , \45815 , \45816 , \45817 , \45818 , \45819 , \45820 ,
         \45821 , \45822 , \45823 , \45824 , \45825 , \45826 , \45827 , \45828 , \45829 , \45830 ,
         \45831 , \45832 , \45833 , \45834 , \45835 , \45836 , \45837 , \45838 , \45839 , \45840 ,
         \45841 , \45842 , \45843 , \45844 , \45845 , \45846 , \45847 , \45848 , \45849 , \45850 ,
         \45851 , \45852 , \45853 , \45854 , \45855 , \45856 , \45857 , \45858 , \45859 , \45860 ,
         \45861 , \45862 , \45863 , \45864 , \45865 , \45866 , \45867 , \45868 , \45869 , \45870 ,
         \45871 , \45872 , \45873 , \45874 , \45875 , \45876 , \45877 , \45878 , \45879 , \45880 ,
         \45881 , \45882 , \45883 , \45884 , \45885 , \45886 , \45887 , \45888 , \45889 , \45890 ,
         \45891 , \45892 , \45893 , \45894 , \45895 , \45896 , \45897 , \45898 , \45899 , \45900 ,
         \45901 , \45902 , \45903 , \45904 , \45905 , \45906 , \45907 , \45908 , \45909 , \45910 ,
         \45911 , \45912 , \45913 , \45914 , \45915 , \45916 , \45917 , \45918 , \45919 , \45920 ,
         \45921 , \45922 , \45923 , \45924 , \45925 , \45926 , \45927 , \45928 , \45929 , \45930 ,
         \45931 , \45932 , \45933 , \45934 , \45935 , \45936 , \45937 , \45938 , \45939 , \45940 ,
         \45941 , \45942 , \45943 , \45944 , \45945 , \45946 , \45947 , \45948 , \45949 , \45950 ,
         \45951 , \45952 , \45953 , \45954 , \45955 , \45956 , \45957 , \45958 , \45959 , \45960 ,
         \45961 , \45962 , \45963 , \45964 , \45965 , \45966 , \45967 , \45968 , \45969 , \45970 ,
         \45971 , \45972 , \45973 , \45974 , \45975 , \45976 , \45977 , \45978 , \45979 , \45980 ,
         \45981 , \45982 , \45983 , \45984 , \45985 , \45986 , \45987 , \45988 , \45989 , \45990 ,
         \45991 , \45992 , \45993 , \45994 , \45995 , \45996 , \45997 , \45998 , \45999 , \46000 ,
         \46001 , \46002 , \46003 , \46004 , \46005 , \46006 , \46007 , \46008 , \46009 , \46010 ,
         \46011 , \46012 , \46013 , \46014 , \46015 , \46016 , \46017 , \46018 , \46019 , \46020 ,
         \46021 , \46022 , \46023 , \46024 , \46025 , \46026 , \46027 , \46028 , \46029 , \46030 ,
         \46031 , \46032 , \46033 , \46034 , \46035 , \46036 , \46037 , \46038 , \46039 , \46040 ,
         \46041 , \46042 , \46043 , \46044 , \46045 , \46046 , \46047 , \46048 , \46049 , \46050 ,
         \46051 , \46052 , \46053 , \46054 , \46055 , \46056 , \46057 , \46058 , \46059 , \46060 ,
         \46061 , \46062 , \46063 , \46064 , \46065 , \46066 , \46067 , \46068 , \46069 , \46070 ,
         \46071 , \46072 , \46073 , \46074 , \46075 , \46076 , \46077 , \46078 , \46079 , \46080 ,
         \46081 , \46082 , \46083 , \46084 , \46085 , \46086 , \46087 , \46088 , \46089 , \46090 ,
         \46091 , \46092 , \46093 , \46094 , \46095 , \46096 , \46097 , \46098 , \46099 , \46100 ,
         \46101 , \46102 , \46103 , \46104 , \46105 , \46106 , \46107 , \46108 , \46109 , \46110 ,
         \46111 , \46112 , \46113 , \46114 , \46115 , \46116 , \46117 , \46118 , \46119 , \46120 ,
         \46121 , \46122 , \46123 , \46124 , \46125 , \46126 , \46127 , \46128 , \46129 , \46130 ,
         \46131 , \46132 , \46133 , \46134 , \46135 , \46136 , \46137 , \46138 , \46139 , \46140 ,
         \46141 , \46142 , \46143 , \46144 , \46145 , \46146 , \46147 , \46148 , \46149 , \46150 ,
         \46151 , \46152 , \46153 , \46154 , \46155 , \46156 , \46157 , \46158 , \46159 , \46160 ,
         \46161 , \46162 , \46163 , \46164 , \46165 , \46166 , \46167 , \46168 , \46169 , \46170 ,
         \46171 , \46172 , \46173 , \46174 , \46175 , \46176 , \46177 , \46178 , \46179 , \46180 ,
         \46181 , \46182 , \46183 , \46184 , \46185 , \46186 , \46187 , \46188 , \46189 , \46190 ,
         \46191 , \46192 , \46193 , \46194 , \46195 , \46196 , \46197 , \46198 , \46199 , \46200 ,
         \46201 , \46202 , \46203 , \46204 , \46205 , \46206 , \46207 , \46208 , \46209 , \46210 ,
         \46211 , \46212 , \46213 , \46214 , \46215 , \46216 , \46217 , \46218 , \46219 , \46220 ,
         \46221 , \46222 , \46223 , \46224 , \46225 , \46226 , \46227 , \46228 , \46229 , \46230 ,
         \46231 , \46232 , \46233 , \46234 , \46235 , \46236 , \46237 , \46238 , \46239 , \46240 ,
         \46241 , \46242 , \46243 , \46244 , \46245 , \46246 , \46247 , \46248 , \46249 , \46250 ,
         \46251 , \46252 , \46253 , \46254 , \46255 , \46256 , \46257 , \46258 , \46259 , \46260 ,
         \46261 , \46262 , \46263 , \46264 , \46265 , \46266 , \46267 , \46268 , \46269 , \46270 ,
         \46271 , \46272 , \46273 , \46274 , \46275 , \46276 , \46277 , \46278 , \46279 , \46280 ,
         \46281 , \46282 , \46283 , \46284 , \46285 , \46286 , \46287 , \46288 , \46289 , \46290 ,
         \46291 , \46292 , \46293 , \46294 , \46295 , \46296 , \46297 , \46298 , \46299 , \46300 ,
         \46301 , \46302 , \46303 , \46304 , \46305 , \46306 , \46307 , \46308 , \46309 , \46310 ,
         \46311 , \46312 , \46313 , \46314 , \46315 , \46316 , \46317 , \46318 , \46319 , \46320 ,
         \46321 , \46322 , \46323 , \46324 , \46325 , \46326 , \46327 , \46328 , \46329 , \46330 ,
         \46331 , \46332 , \46333 , \46334 , \46335 , \46336 , \46337 , \46338 , \46339 , \46340 ,
         \46341 , \46342 , \46343 , \46344 , \46345 , \46346 , \46347 , \46348 , \46349 , \46350 ,
         \46351 , \46352 , \46353 , \46354 , \46355 , \46356 , \46357 , \46358 , \46359 , \46360 ,
         \46361 , \46362 , \46363 , \46364 , \46365 , \46366 , \46367 , \46368 , \46369 , \46370 ,
         \46371 , \46372 , \46373 , \46374 , \46375 , \46376 , \46377 , \46378 , \46379 , \46380 ,
         \46381 , \46382 , \46383 , \46384 , \46385 , \46386 , \46387 , \46388 , \46389 , \46390 ,
         \46391 , \46392 , \46393 , \46394 , \46395 , \46396 , \46397 , \46398 , \46399 , \46400 ,
         \46401 , \46402 , \46403 , \46404 , \46405 , \46406 , \46407 , \46408 , \46409 , \46410 ,
         \46411 , \46412 , \46413 , \46414 , \46415 , \46416 , \46417 , \46418 , \46419 , \46420 ,
         \46421 , \46422 , \46423 , \46424 , \46425 , \46426 , \46427 , \46428 , \46429 , \46430 ,
         \46431 , \46432 , \46433 , \46434 , \46435 , \46436 , \46437 , \46438 , \46439 , \46440 ,
         \46441 , \46442 , \46443 , \46444 , \46445 , \46446 , \46447 , \46448 , \46449 , \46450 ,
         \46451 , \46452 , \46453 , \46454 , \46455 , \46456 , \46457 , \46458 , \46459 , \46460 ,
         \46461 , \46462 , \46463 , \46464 , \46465 , \46466 , \46467 , \46468 , \46469 , \46470 ,
         \46471 , \46472 , \46473 , \46474 , \46475 , \46476 , \46477 , \46478 , \46479 , \46480 ,
         \46481 , \46482 , \46483 , \46484 , \46485 , \46486 , \46487 , \46488 , \46489 , \46490 ,
         \46491 , \46492 , \46493 , \46494 , \46495 , \46496 , \46497 , \46498 , \46499 , \46500 ,
         \46501 , \46502 , \46503 , \46504 , \46505 , \46506 , \46507 , \46508 , \46509 , \46510 ,
         \46511 , \46512 , \46513 , \46514 , \46515 , \46516 , \46517 , \46518 , \46519 , \46520 ,
         \46521 , \46522 , \46523 , \46524 , \46525 , \46526 , \46527 , \46528 , \46529 , \46530 ,
         \46531 , \46532 , \46533 , \46534 , \46535 , \46536 , \46537 , \46538 , \46539 , \46540 ,
         \46541 , \46542 , \46543 , \46544 , \46545 , \46546 , \46547 , \46548 , \46549 , \46550 ,
         \46551 , \46552 , \46553 , \46554 , \46555 , \46556 , \46557 , \46558 , \46559 , \46560 ,
         \46561 , \46562 , \46563 , \46564 , \46565 , \46566 , \46567 , \46568 , \46569 , \46570 ,
         \46571 , \46572 , \46573 , \46574 , \46575 , \46576 , \46577 , \46578 , \46579 , \46580 ,
         \46581 , \46582 , \46583 , \46584 , \46585 , \46586 , \46587 , \46588 , \46589 , \46590 ,
         \46591 , \46592 , \46593 , \46594 , \46595 , \46596 , \46597 , \46598 , \46599 , \46600 ,
         \46601 , \46602 , \46603 , \46604 , \46605 , \46606 , \46607 , \46608 , \46609 , \46610 ,
         \46611 , \46612 , \46613 , \46614 , \46615 , \46616 , \46617 , \46618 , \46619 , \46620 ,
         \46621 , \46622 , \46623 , \46624 , \46625 , \46626 , \46627 , \46628 , \46629 , \46630 ,
         \46631 , \46632 , \46633 , \46634 , \46635 , \46636 , \46637 , \46638 , \46639 , \46640 ,
         \46641 , \46642 , \46643 , \46644 , \46645 , \46646 , \46647 , \46648 , \46649 , \46650 ,
         \46651 , \46652 , \46653 , \46654 , \46655 , \46656 , \46657 , \46658 , \46659 , \46660 ,
         \46661 , \46662 , \46663 , \46664 , \46665 , \46666 , \46667 , \46668 , \46669 , \46670 ,
         \46671 , \46672 , \46673 , \46674 , \46675 , \46676 , \46677 , \46678 , \46679 , \46680 ,
         \46681 , \46682 , \46683 , \46684 , \46685 , \46686 , \46687 , \46688 , \46689 , \46690 ,
         \46691 , \46692 , \46693 , \46694 , \46695 , \46696 , \46697 , \46698 , \46699 , \46700 ,
         \46701 , \46702 , \46703 , \46704 , \46705 , \46706 , \46707 , \46708 , \46709 , \46710 ,
         \46711 , \46712 , \46713 , \46714 , \46715 , \46716 , \46717 , \46718 , \46719 , \46720 ,
         \46721 , \46722 , \46723 , \46724 , \46725 , \46726 , \46727 , \46728 , \46729 , \46730 ,
         \46731 , \46732 , \46733 , \46734 , \46735 , \46736 , \46737 , \46738 , \46739 , \46740 ,
         \46741 , \46742 , \46743 , \46744 , \46745 , \46746 , \46747 , \46748 , \46749 , \46750 ,
         \46751 , \46752 , \46753 , \46754 , \46755 , \46756 , \46757 , \46758 , \46759 , \46760 ,
         \46761 , \46762 , \46763 , \46764 , \46765 , \46766 , \46767 , \46768 , \46769 , \46770 ,
         \46771 , \46772 , \46773 , \46774 , \46775 , \46776 , \46777 , \46778 , \46779 , \46780 ,
         \46781 , \46782 , \46783 , \46784 , \46785 , \46786 , \46787 , \46788 , \46789 , \46790 ,
         \46791 , \46792 , \46793 , \46794 , \46795 , \46796 , \46797 , \46798 , \46799 , \46800 ,
         \46801 , \46802 , \46803 , \46804 , \46805 , \46806 , \46807 , \46808 , \46809 , \46810 ,
         \46811 , \46812 , \46813 , \46814 , \46815 , \46816 , \46817 , \46818 , \46819 , \46820 ,
         \46821 , \46822 , \46823 , \46824 , \46825 , \46826 , \46827 , \46828 , \46829 , \46830 ,
         \46831 , \46832 , \46833 , \46834 , \46835 , \46836 , \46837 , \46838 , \46839 , \46840 ,
         \46841 , \46842 , \46843 , \46844 , \46845 , \46846 , \46847 , \46848 , \46849 , \46850 ,
         \46851 , \46852 , \46853 , \46854 , \46855 , \46856 , \46857 , \46858 , \46859 , \46860 ,
         \46861 , \46862 , \46863 , \46864 , \46865 , \46866 , \46867 , \46868 , \46869 , \46870 ,
         \46871 , \46872 , \46873 , \46874 , \46875 , \46876 , \46877 , \46878 , \46879 , \46880 ,
         \46881 , \46882 , \46883 , \46884 , \46885 , \46886 , \46887 , \46888 , \46889 , \46890 ,
         \46891 , \46892 , \46893 , \46894 , \46895 , \46896 , \46897 , \46898 , \46899 , \46900 ,
         \46901 , \46902 , \46903 , \46904 , \46905 , \46906 , \46907 , \46908 , \46909 , \46910 ,
         \46911 , \46912 , \46913 , \46914 , \46915 , \46916 , \46917 , \46918 , \46919 , \46920 ,
         \46921 , \46922 , \46923 , \46924 , \46925 , \46926 , \46927 , \46928 , \46929 , \46930 ,
         \46931 , \46932 , \46933 , \46934 , \46935 , \46936 , \46937 , \46938 , \46939 , \46940 ,
         \46941 , \46942 , \46943 , \46944 , \46945 , \46946 , \46947 , \46948 , \46949 , \46950 ,
         \46951 , \46952 , \46953 , \46954 , \46955 , \46956 , \46957 , \46958 , \46959 , \46960 ,
         \46961 , \46962 , \46963 , \46964 , \46965 , \46966 , \46967 , \46968 , \46969 , \46970 ,
         \46971 , \46972 , \46973 , \46974 , \46975 , \46976 , \46977 , \46978 , \46979 , \46980 ,
         \46981 , \46982 , \46983 , \46984 , \46985 , \46986 , \46987 , \46988 , \46989 , \46990 ,
         \46991 , \46992 , \46993 , \46994 , \46995 , \46996 , \46997 , \46998 , \46999 , \47000 ,
         \47001 , \47002 , \47003 , \47004 , \47005 , \47006 , \47007 , \47008 , \47009 , \47010 ,
         \47011 , \47012 , \47013 , \47014 , \47015 , \47016 , \47017 , \47018 , \47019 , \47020 ,
         \47021 , \47022 , \47023 , \47024 , \47025 , \47026 , \47027 , \47028 , \47029 , \47030 ,
         \47031 , \47032 , \47033 , \47034 , \47035 , \47036 , \47037 , \47038 , \47039 , \47040 ,
         \47041 , \47042 , \47043 , \47044 , \47045 , \47046 , \47047 , \47048 , \47049 , \47050 ,
         \47051 , \47052 , \47053 , \47054 , \47055 , \47056 , \47057 , \47058 , \47059 , \47060 ,
         \47061 , \47062 , \47063 , \47064 , \47065 , \47066 , \47067 , \47068 , \47069 , \47070 ,
         \47071 , \47072 , \47073 , \47074 , \47075 , \47076 , \47077 , \47078 , \47079 , \47080 ,
         \47081 , \47082 , \47083 , \47084 , \47085 , \47086 , \47087 , \47088 , \47089 , \47090 ,
         \47091 , \47092 , \47093 , \47094 , \47095 , \47096 , \47097 , \47098 , \47099 , \47100 ,
         \47101 , \47102 , \47103 , \47104 , \47105 , \47106 , \47107 , \47108 , \47109 , \47110 ,
         \47111 , \47112 , \47113 , \47114 , \47115 , \47116 , \47117 , \47118 , \47119 , \47120 ,
         \47121 , \47122 , \47123 , \47124 , \47125 , \47126 , \47127 , \47128 , \47129 , \47130 ,
         \47131 , \47132 , \47133 , \47134 , \47135 , \47136 , \47137 , \47138 , \47139 , \47140 ,
         \47141 , \47142 , \47143 , \47144 , \47145 , \47146 , \47147 , \47148 , \47149 , \47150 ,
         \47151 , \47152 , \47153 , \47154 , \47155 , \47156 , \47157 , \47158 , \47159 , \47160 ,
         \47161 , \47162 , \47163 , \47164 , \47165 , \47166 , \47167 , \47168 , \47169 , \47170 ,
         \47171 , \47172 , \47173 , \47174 , \47175 , \47176 , \47177 , \47178 , \47179 , \47180 ,
         \47181 , \47182 , \47183 , \47184 , \47185 , \47186 , \47187 , \47188 , \47189 , \47190 ,
         \47191 , \47192 , \47193 , \47194 , \47195 , \47196 , \47197 , \47198 , \47199 , \47200 ,
         \47201 , \47202 , \47203 , \47204 , \47205 , \47206 , \47207 , \47208 , \47209 , \47210 ,
         \47211 , \47212 , \47213 , \47214 , \47215 , \47216 , \47217 , \47218 , \47219 , \47220 ,
         \47221 , \47222 , \47223 , \47224 , \47225 , \47226 , \47227 , \47228 , \47229 , \47230 ,
         \47231 , \47232 , \47233 , \47234 , \47235 , \47236 , \47237 , \47238 , \47239 , \47240 ,
         \47241 , \47242 , \47243 , \47244 , \47245 , \47246 , \47247 , \47248 , \47249 , \47250 ,
         \47251 , \47252 , \47253 , \47254 , \47255 , \47256 , \47257 , \47258 , \47259 , \47260 ,
         \47261 , \47262 , \47263 , \47264 , \47265 , \47266 , \47267 , \47268 , \47269 , \47270 ,
         \47271 , \47272 , \47273 , \47274 , \47275 , \47276 , \47277 , \47278 , \47279 , \47280 ,
         \47281 , \47282 , \47283 , \47284 , \47285 , \47286 , \47287 , \47288 , \47289 , \47290 ,
         \47291 , \47292 , \47293 , \47294 , \47295 , \47296 , \47297 , \47298 , \47299 , \47300 ,
         \47301 , \47302 , \47303 , \47304 , \47305 , \47306 , \47307 , \47308 , \47309 , \47310 ,
         \47311 , \47312 , \47313 , \47314 , \47315 , \47316 , \47317 , \47318 , \47319 , \47320 ,
         \47321 , \47322 , \47323 , \47324 , \47325 , \47326 , \47327 , \47328 , \47329 , \47330 ,
         \47331 , \47332 , \47333 , \47334 , \47335 , \47336 , \47337 , \47338 , \47339 , \47340 ,
         \47341 , \47342 , \47343 , \47344 , \47345 , \47346 , \47347 , \47348 , \47349 , \47350 ,
         \47351 , \47352 , \47353 , \47354 , \47355 , \47356 , \47357 , \47358 , \47359 , \47360 ,
         \47361 , \47362 , \47363 , \47364 , \47365 , \47366 , \47367 , \47368 , \47369 , \47370 ,
         \47371 , \47372 , \47373 , \47374 , \47375 , \47376 , \47377 , \47378 , \47379 , \47380 ,
         \47381 , \47382 , \47383 , \47384 , \47385 , \47386 , \47387 , \47388 , \47389 , \47390 ,
         \47391 , \47392 , \47393 , \47394 , \47395 , \47396 , \47397 , \47398 , \47399 , \47400 ,
         \47401 , \47402 , \47403 , \47404 , \47405 , \47406 , \47407 , \47408 , \47409 , \47410 ,
         \47411 , \47412 , \47413 , \47414 , \47415 , \47416 , \47417 , \47418 , \47419 , \47420 ,
         \47421 , \47422 , \47423 , \47424 , \47425 , \47426 , \47427 , \47428 , \47429 , \47430 ,
         \47431 , \47432 , \47433 , \47434 , \47435 , \47436 , \47437 , \47438 , \47439 , \47440 ,
         \47441 , \47442 , \47443 , \47444 , \47445 , \47446 , \47447 , \47448 , \47449 , \47450 ,
         \47451 , \47452 , \47453 , \47454 , \47455 , \47456 , \47457 , \47458 , \47459 , \47460 ,
         \47461 , \47462 , \47463 , \47464 , \47465 , \47466 , \47467 , \47468 , \47469 , \47470 ,
         \47471 , \47472 , \47473 , \47474 , \47475 , \47476 , \47477 , \47478 , \47479 , \47480 ,
         \47481 , \47482 , \47483 , \47484 , \47485 , \47486 , \47487 , \47488 , \47489 , \47490 ,
         \47491 , \47492 , \47493 , \47494 , \47495 , \47496 , \47497 , \47498 , \47499 , \47500 ,
         \47501 , \47502 , \47503 , \47504 , \47505 , \47506 , \47507 , \47508 , \47509 , \47510 ,
         \47511 , \47512 , \47513 , \47514 , \47515 , \47516 , \47517 , \47518 , \47519 , \47520 ,
         \47521 , \47522 , \47523 , \47524 , \47525 , \47526 , \47527 , \47528 , \47529 , \47530 ,
         \47531 , \47532 , \47533 , \47534 , \47535 , \47536 , \47537 , \47538 , \47539 , \47540 ,
         \47541 , \47542 , \47543 , \47544 , \47545 , \47546 , \47547 , \47548 , \47549 , \47550 ,
         \47551 , \47552 , \47553 , \47554 , \47555 , \47556 , \47557 , \47558 , \47559 , \47560 ,
         \47561 , \47562 , \47563 , \47564 , \47565 , \47566 , \47567 , \47568 , \47569 , \47570 ,
         \47571 , \47572 , \47573 , \47574 , \47575 , \47576 , \47577 , \47578 , \47579 , \47580 ,
         \47581 , \47582 , \47583 , \47584 , \47585 , \47586 , \47587 , \47588 , \47589 , \47590 ,
         \47591 , \47592 , \47593 , \47594 , \47595 , \47596 , \47597 , \47598 , \47599 , \47600 ,
         \47601 , \47602 , \47603 , \47604 , \47605 , \47606 , \47607 , \47608 , \47609 , \47610 ,
         \47611 , \47612 , \47613 , \47614 , \47615 , \47616 , \47617 , \47618 , \47619 , \47620 ,
         \47621 , \47622 , \47623 , \47624 , \47625 , \47626 , \47627 , \47628 , \47629 , \47630 ,
         \47631 , \47632 , \47633 , \47634 , \47635 , \47636 , \47637 , \47638 , \47639 , \47640 ,
         \47641 , \47642 , \47643 , \47644 , \47645 , \47646 , \47647 , \47648 , \47649 , \47650 ,
         \47651 , \47652 , \47653 , \47654 , \47655 , \47656 , \47657 , \47658 , \47659 , \47660 ,
         \47661 , \47662 , \47663 , \47664 , \47665 , \47666 , \47667 , \47668 , \47669 , \47670 ,
         \47671 , \47672 , \47673 , \47674 , \47675 , \47676 , \47677 , \47678 , \47679 , \47680 ,
         \47681 , \47682 , \47683 , \47684 , \47685 , \47686 , \47687 , \47688 , \47689 , \47690 ,
         \47691 , \47692 , \47693 , \47694 , \47695 , \47696 , \47697 , \47698 , \47699 , \47700 ,
         \47701 , \47702 , \47703 , \47704 , \47705 , \47706 , \47707 , \47708 , \47709 , \47710 ,
         \47711 , \47712 , \47713 , \47714 , \47715 , \47716 , \47717 , \47718 , \47719 , \47720 ,
         \47721 , \47722 , \47723 , \47724 , \47725 , \47726 , \47727 , \47728 , \47729 , \47730 ,
         \47731 , \47732 , \47733 , \47734 , \47735 , \47736 , \47737 , \47738 , \47739 , \47740 ,
         \47741 , \47742 , \47743 , \47744 , \47745 , \47746 , \47747 , \47748 , \47749 , \47750 ,
         \47751 , \47752 , \47753 , \47754 , \47755 , \47756 , \47757 , \47758 , \47759 , \47760 ,
         \47761 , \47762 , \47763 , \47764 , \47765 , \47766 , \47767 , \47768 , \47769 , \47770 ,
         \47771 , \47772 , \47773 , \47774 , \47775 , \47776 , \47777 , \47778 , \47779 , \47780 ,
         \47781 , \47782 , \47783 , \47784 , \47785 , \47786 , \47787 , \47788 , \47789 , \47790 ,
         \47791 , \47792 , \47793 , \47794 , \47795 , \47796 , \47797 , \47798 , \47799 , \47800 ,
         \47801 , \47802 , \47803 , \47804 , \47805 , \47806 , \47807 , \47808 , \47809 , \47810 ,
         \47811 , \47812 , \47813 , \47814 , \47815 , \47816 , \47817 , \47818 , \47819 , \47820 ,
         \47821 , \47822 , \47823 , \47824 , \47825 , \47826 , \47827 , \47828 , \47829 , \47830 ,
         \47831 , \47832 , \47833 , \47834 , \47835 , \47836 , \47837 , \47838 , \47839 , \47840 ,
         \47841 , \47842 , \47843 , \47844 , \47845 , \47846 , \47847 , \47848 , \47849 , \47850 ,
         \47851 , \47852 , \47853 , \47854 , \47855 , \47856 , \47857 , \47858 , \47859 , \47860 ,
         \47861 , \47862 , \47863 , \47864 , \47865 , \47866 , \47867 , \47868 , \47869 , \47870 ,
         \47871 , \47872 , \47873 , \47874 , \47875 , \47876 , \47877 , \47878 , \47879 , \47880 ,
         \47881 , \47882 , \47883 , \47884 , \47885 , \47886 , \47887 , \47888 , \47889 , \47890 ,
         \47891 , \47892 , \47893 , \47894 , \47895 , \47896 , \47897 , \47898 , \47899 , \47900 ,
         \47901 , \47902 , \47903 , \47904 , \47905 , \47906 , \47907 , \47908 , \47909 , \47910 ,
         \47911 , \47912 , \47913 , \47914 , \47915 , \47916 , \47917 , \47918 , \47919 , \47920 ,
         \47921 , \47922 , \47923 , \47924 , \47925 , \47926 , \47927 , \47928 , \47929 , \47930 ,
         \47931 , \47932 , \47933 , \47934 , \47935 , \47936 , \47937 , \47938 , \47939 , \47940 ,
         \47941 , \47942 , \47943 , \47944 , \47945 , \47946 , \47947 , \47948 , \47949 , \47950 ,
         \47951 , \47952 , \47953 , \47954 , \47955 , \47956 , \47957 , \47958 , \47959 , \47960 ,
         \47961 , \47962 , \47963 , \47964 , \47965 , \47966 , \47967 , \47968 , \47969 , \47970 ,
         \47971 , \47972 , \47973 , \47974 , \47975 , \47976 , \47977 , \47978 , \47979 , \47980 ,
         \47981 , \47982 , \47983 , \47984 , \47985 , \47986 , \47987 , \47988 , \47989 , \47990 ,
         \47991 , \47992 , \47993 , \47994 , \47995 , \47996 , \47997 , \47998 , \47999 , \48000 ,
         \48001 , \48002 , \48003 , \48004 , \48005 , \48006 , \48007 , \48008 , \48009 , \48010 ,
         \48011 , \48012 , \48013 , \48014 , \48015 , \48016 , \48017 , \48018 , \48019 , \48020 ,
         \48021 , \48022 , \48023 , \48024 , \48025 , \48026 , \48027 , \48028 , \48029 , \48030 ,
         \48031 , \48032 , \48033 , \48034 , \48035 , \48036 , \48037 , \48038 , \48039 , \48040 ,
         \48041 , \48042 , \48043 , \48044 , \48045 , \48046 , \48047 , \48048 , \48049 , \48050 ,
         \48051 , \48052 , \48053 , \48054 , \48055 , \48056 , \48057 , \48058 , \48059 , \48060 ,
         \48061 , \48062 , \48063 , \48064 , \48065 , \48066 , \48067 , \48068 , \48069 , \48070 ,
         \48071 , \48072 , \48073 , \48074 , \48075 , \48076 , \48077 , \48078 , \48079 , \48080 ,
         \48081 , \48082 , \48083 , \48084 , \48085 , \48086 , \48087 , \48088 , \48089 , \48090 ,
         \48091 , \48092 , \48093 , \48094 , \48095 , \48096 , \48097 , \48098 , \48099 , \48100 ,
         \48101 , \48102 , \48103 , \48104 , \48105 , \48106 , \48107 , \48108 , \48109 , \48110 ,
         \48111 , \48112 , \48113 , \48114 , \48115 , \48116 , \48117 , \48118 , \48119 , \48120 ,
         \48121 , \48122 , \48123 , \48124 , \48125 , \48126 , \48127 , \48128 , \48129 , \48130 ,
         \48131 , \48132 , \48133 , \48134 , \48135 , \48136 , \48137 , \48138 , \48139 , \48140 ,
         \48141 , \48142 , \48143 , \48144 , \48145 , \48146 , \48147 , \48148 , \48149 , \48150 ,
         \48151 , \48152 , \48153 , \48154 , \48155 , \48156 , \48157 , \48158 , \48159 , \48160 ,
         \48161 , \48162 , \48163 , \48164 , \48165 , \48166 , \48167 , \48168 , \48169 , \48170 ,
         \48171 , \48172 , \48173 , \48174 , \48175 , \48176 , \48177 , \48178 , \48179 , \48180 ,
         \48181 , \48182 , \48183 , \48184 , \48185 , \48186 , \48187 , \48188 , \48189 , \48190 ,
         \48191 , \48192 , \48193 , \48194 , \48195 , \48196 , \48197 , \48198 , \48199 , \48200 ,
         \48201 , \48202 , \48203 , \48204 , \48205 , \48206 , \48207 , \48208 , \48209 , \48210 ,
         \48211 , \48212 , \48213 , \48214 , \48215 , \48216 , \48217 , \48218 , \48219 , \48220 ,
         \48221 , \48222 , \48223 , \48224 , \48225 , \48226 , \48227 , \48228 , \48229 , \48230 ,
         \48231 , \48232 , \48233 , \48234 , \48235 , \48236 , \48237 , \48238 , \48239 , \48240 ,
         \48241 , \48242 , \48243 , \48244 , \48245 , \48246 , \48247 , \48248 , \48249 , \48250 ,
         \48251 , \48252 , \48253 , \48254 , \48255 , \48256 , \48257 , \48258 , \48259 , \48260 ,
         \48261 , \48262 , \48263 , \48264 , \48265 , \48266 , \48267 , \48268 , \48269 , \48270 ,
         \48271 , \48272 , \48273 , \48274 , \48275 , \48276 , \48277 , \48278 , \48279 , \48280 ,
         \48281 , \48282 , \48283 , \48284 , \48285 , \48286 , \48287 , \48288 , \48289 , \48290 ,
         \48291 , \48292 , \48293 , \48294 , \48295 , \48296 , \48297 , \48298 , \48299 , \48300 ,
         \48301 , \48302 , \48303 , \48304 , \48305 , \48306 , \48307 , \48308 , \48309 , \48310 ,
         \48311 , \48312 , \48313 , \48314 , \48315 , \48316 , \48317 , \48318 , \48319 , \48320 ,
         \48321 , \48322 , \48323 , \48324 , \48325 , \48326 , \48327 , \48328 , \48329 , \48330 ,
         \48331 , \48332 , \48333 , \48334 , \48335 , \48336 , \48337 , \48338 , \48339 , \48340 ,
         \48341 , \48342 , \48343 , \48344 , \48345 , \48346 , \48347 , \48348 , \48349 , \48350 ,
         \48351 , \48352 , \48353 , \48354 , \48355 , \48356 , \48357 , \48358 , \48359 , \48360 ,
         \48361 , \48362 , \48363 , \48364 , \48365 , \48366 , \48367 , \48368 , \48369 , \48370 ,
         \48371 , \48372 , \48373 , \48374 , \48375 , \48376 , \48377 , \48378 , \48379 , \48380 ,
         \48381 , \48382 , \48383 , \48384 , \48385 , \48386 , \48387 , \48388 , \48389 , \48390 ,
         \48391 , \48392 , \48393 , \48394 , \48395 , \48396 , \48397 , \48398 , \48399 , \48400 ,
         \48401 , \48402 , \48403 , \48404 , \48405 , \48406 , \48407 , \48408 , \48409 , \48410 ,
         \48411 , \48412 , \48413 , \48414 , \48415 , \48416 , \48417 , \48418 , \48419 , \48420 ,
         \48421 , \48422 , \48423 , \48424 , \48425 , \48426 , \48427 , \48428 , \48429 , \48430 ,
         \48431 , \48432 , \48433 , \48434 , \48435 , \48436 , \48437 , \48438 , \48439 , \48440 ,
         \48441 , \48442 , \48443 , \48444 , \48445 , \48446 , \48447 , \48448 , \48449 , \48450 ,
         \48451 , \48452 , \48453 , \48454 , \48455 , \48456 , \48457 , \48458 , \48459 , \48460 ,
         \48461 , \48462 , \48463 , \48464 , \48465 , \48466 , \48467 , \48468 , \48469 , \48470 ,
         \48471 , \48472 , \48473 , \48474 , \48475 , \48476 , \48477 , \48478 , \48479 , \48480 ,
         \48481 , \48482 , \48483 , \48484 , \48485 , \48486 , \48487 , \48488 , \48489 , \48490 ,
         \48491 , \48492 , \48493 , \48494 , \48495 , \48496 , \48497 , \48498 , \48499 , \48500 ,
         \48501 , \48502 , \48503 , \48504 , \48505 , \48506 , \48507 , \48508 , \48509 , \48510 ,
         \48511 , \48512 , \48513 , \48514 , \48515 , \48516 , \48517 , \48518 , \48519 , \48520 ,
         \48521 , \48522 , \48523 , \48524 , \48525 , \48526 , \48527 , \48528 , \48529 , \48530 ,
         \48531 , \48532 , \48533 , \48534 , \48535 , \48536 , \48537 , \48538 , \48539 , \48540 ,
         \48541 , \48542 , \48543 , \48544 , \48545 , \48546 , \48547 , \48548 , \48549 , \48550 ,
         \48551 , \48552 , \48553 , \48554 , \48555 , \48556 , \48557 , \48558 , \48559 , \48560 ,
         \48561 , \48562 , \48563 , \48564 , \48565 , \48566 , \48567 , \48568 , \48569 , \48570 ,
         \48571 , \48572 , \48573 , \48574 , \48575 , \48576 , \48577 , \48578 , \48579 , \48580 ,
         \48581 , \48582 , \48583 , \48584 , \48585 , \48586 , \48587 , \48588 , \48589 , \48590 ,
         \48591 , \48592 , \48593 , \48594 , \48595 , \48596 , \48597 , \48598 , \48599 , \48600 ,
         \48601 , \48602 , \48603 , \48604 , \48605 , \48606 , \48607 , \48608 , \48609 , \48610 ,
         \48611 , \48612 , \48613 , \48614 , \48615 , \48616 , \48617 , \48618 , \48619 , \48620 ,
         \48621 , \48622 , \48623 , \48624 , \48625 , \48626 , \48627 , \48628 , \48629 , \48630 ,
         \48631 , \48632 , \48633 , \48634 , \48635 , \48636 , \48637 , \48638 , \48639 , \48640 ,
         \48641 , \48642 , \48643 , \48644 , \48645 , \48646 , \48647 , \48648 , \48649 , \48650 ,
         \48651 , \48652 , \48653 , \48654 , \48655 , \48656 , \48657 , \48658 , \48659 , \48660 ,
         \48661 , \48662 , \48663 , \48664 , \48665 , \48666 , \48667 , \48668 , \48669 , \48670 ,
         \48671 , \48672 , \48673 , \48674 , \48675 , \48676 , \48677 , \48678 , \48679 , \48680 ,
         \48681 , \48682 , \48683 , \48684 , \48685 , \48686 , \48687 , \48688 , \48689 , \48690 ,
         \48691 , \48692 , \48693 , \48694 , \48695 , \48696 , \48697 , \48698 , \48699 , \48700 ,
         \48701 , \48702 , \48703 , \48704 , \48705 , \48706 , \48707 , \48708 , \48709 , \48710 ,
         \48711 , \48712 , \48713 , \48714 , \48715 , \48716 , \48717 , \48718 , \48719 , \48720 ,
         \48721 , \48722 , \48723 , \48724 , \48725 , \48726 , \48727 , \48728 , \48729 , \48730 ,
         \48731 , \48732 , \48733 , \48734 , \48735 , \48736 , \48737 , \48738 , \48739 , \48740 ,
         \48741 , \48742 , \48743 , \48744 , \48745 , \48746 , \48747 , \48748 , \48749 , \48750 ,
         \48751 , \48752 , \48753 , \48754 , \48755 , \48756 , \48757 , \48758 , \48759 , \48760 ,
         \48761 , \48762 , \48763 , \48764 , \48765 , \48766 , \48767 , \48768 , \48769 , \48770 ,
         \48771 , \48772 , \48773 , \48774 , \48775 , \48776 , \48777 , \48778 , \48779 , \48780 ,
         \48781 , \48782 , \48783 , \48784 , \48785 , \48786 , \48787 , \48788 , \48789 , \48790 ,
         \48791 , \48792 , \48793 , \48794 , \48795 , \48796 , \48797 , \48798 , \48799 , \48800 ,
         \48801 , \48802 , \48803 , \48804 , \48805 , \48806 , \48807 , \48808 , \48809 , \48810 ,
         \48811 , \48812 , \48813 , \48814 , \48815 , \48816 , \48817 , \48818 , \48819 , \48820 ,
         \48821 , \48822 , \48823 , \48824 , \48825 , \48826 , \48827 , \48828 , \48829 , \48830 ,
         \48831 , \48832 , \48833 , \48834 , \48835 , \48836 , \48837 , \48838 , \48839 , \48840 ,
         \48841 , \48842 , \48843 , \48844 , \48845 , \48846 , \48847 , \48848 , \48849 , \48850 ,
         \48851 , \48852 , \48853 , \48854 , \48855 , \48856 , \48857 , \48858 , \48859 , \48860 ,
         \48861 , \48862 , \48863 , \48864 , \48865 , \48866 , \48867 , \48868 , \48869 , \48870 ,
         \48871 , \48872 , \48873 , \48874 , \48875 , \48876 , \48877 , \48878 , \48879 , \48880 ,
         \48881 , \48882 , \48883 , \48884 , \48885 , \48886 , \48887 , \48888 , \48889 , \48890 ,
         \48891 , \48892 , \48893 , \48894 , \48895 , \48896 , \48897 , \48898 , \48899 , \48900 ,
         \48901 , \48902 , \48903 , \48904 , \48905 , \48906 , \48907 , \48908 , \48909 , \48910 ,
         \48911 , \48912 , \48913 , \48914 , \48915 , \48916 , \48917 , \48918 , \48919 , \48920 ,
         \48921 , \48922 , \48923 , \48924 , \48925 , \48926 , \48927 , \48928 , \48929 , \48930 ,
         \48931 , \48932 , \48933 , \48934 , \48935 , \48936 , \48937 , \48938 , \48939 , \48940 ,
         \48941 , \48942 , \48943 , \48944 , \48945 , \48946 , \48947 , \48948 , \48949 , \48950 ,
         \48951 , \48952 , \48953 , \48954 , \48955 , \48956 , \48957 , \48958 , \48959 , \48960 ,
         \48961 , \48962 , \48963 , \48964 , \48965 , \48966 , \48967 , \48968 , \48969 , \48970 ,
         \48971 , \48972 , \48973 , \48974 , \48975 , \48976 , \48977 , \48978 , \48979 , \48980 ,
         \48981 , \48982 , \48983 , \48984 , \48985 , \48986 , \48987 , \48988 , \48989 , \48990 ,
         \48991 , \48992 , \48993 , \48994 , \48995 , \48996 , \48997 , \48998 , \48999 , \49000 ,
         \49001 , \49002 , \49003 , \49004 , \49005 , \49006 , \49007 , \49008 , \49009 , \49010 ,
         \49011 , \49012 , \49013 , \49014 , \49015 , \49016 , \49017 , \49018 , \49019 , \49020 ,
         \49021 , \49022 , \49023 , \49024 , \49025 , \49026 , \49027 , \49028 , \49029 , \49030 ,
         \49031 , \49032 , \49033 , \49034 , \49035 , \49036 , \49037 , \49038 , \49039 , \49040 ,
         \49041 , \49042 , \49043 , \49044 , \49045 , \49046 , \49047 , \49048 , \49049 , \49050 ,
         \49051 , \49052 , \49053 , \49054 , \49055 , \49056 , \49057 , \49058 , \49059 , \49060 ,
         \49061 , \49062 , \49063 , \49064 , \49065 , \49066 , \49067 , \49068 , \49069 , \49070 ,
         \49071 , \49072 , \49073 , \49074 , \49075 , \49076 , \49077 , \49078 , \49079 , \49080 ,
         \49081 , \49082 , \49083 , \49084 , \49085 , \49086 , \49087 , \49088 , \49089 , \49090 ,
         \49091 , \49092 , \49093 , \49094 , \49095 , \49096 , \49097 , \49098 , \49099 , \49100 ,
         \49101 , \49102 , \49103 , \49104 , \49105 , \49106 , \49107 , \49108 , \49109 , \49110 ,
         \49111 , \49112 , \49113 , \49114 , \49115 , \49116 , \49117 , \49118 , \49119 , \49120 ,
         \49121 , \49122 , \49123 , \49124 , \49125 , \49126 , \49127 , \49128 , \49129 , \49130 ,
         \49131 , \49132 , \49133 , \49134 , \49135 , \49136 , \49137 , \49138 , \49139 , \49140 ,
         \49141 , \49142 , \49143 , \49144 , \49145 , \49146 , \49147 , \49148 , \49149 , \49150 ,
         \49151 , \49152 , \49153 , \49154 , \49155 , \49156 , \49157 , \49158 , \49159 , \49160 ,
         \49161 , \49162 , \49163 , \49164 , \49165 , \49166 , \49167 , \49168 , \49169 , \49170 ,
         \49171 , \49172 , \49173 , \49174 , \49175 , \49176 , \49177 , \49178 , \49179 , \49180 ,
         \49181 , \49182 , \49183 , \49184 , \49185 , \49186 , \49187 , \49188 , \49189 , \49190 ,
         \49191 , \49192 , \49193 , \49194 , \49195 , \49196 , \49197 , \49198 , \49199 , \49200 ,
         \49201 , \49202 , \49203 , \49204 , \49205 , \49206 , \49207 , \49208 , \49209 , \49210 ,
         \49211 , \49212 , \49213 , \49214 , \49215 , \49216 , \49217 , \49218 , \49219 , \49220 ,
         \49221 , \49222 , \49223 , \49224 , \49225 , \49226 , \49227 , \49228 , \49229 , \49230 ,
         \49231 , \49232 , \49233 , \49234 , \49235 , \49236 , \49237 , \49238 , \49239 , \49240 ,
         \49241 , \49242 , \49243 , \49244 , \49245 , \49246 , \49247 , \49248 , \49249 , \49250 ,
         \49251 , \49252 , \49253 , \49254 , \49255 , \49256 , \49257 , \49258 , \49259 , \49260 ,
         \49261 , \49262 , \49263 , \49264 , \49265 , \49266 , \49267 , \49268 , \49269 , \49270 ,
         \49271 , \49272 , \49273 , \49274 , \49275 , \49276 , \49277 , \49278 , \49279 , \49280 ,
         \49281 , \49282 , \49283 , \49284 , \49285 , \49286 , \49287 , \49288 , \49289 , \49290 ,
         \49291 , \49292 , \49293 , \49294 , \49295 , \49296 , \49297 , \49298 , \49299 , \49300 ,
         \49301 , \49302 , \49303 , \49304 , \49305 , \49306 , \49307 , \49308 , \49309 , \49310 ,
         \49311 , \49312 , \49313 , \49314 , \49315 , \49316 , \49317 , \49318 , \49319 , \49320 ,
         \49321 , \49322 , \49323 , \49324 , \49325 , \49326 , \49327 , \49328 , \49329 , \49330 ,
         \49331 , \49332 , \49333 , \49334 , \49335 , \49336 , \49337 , \49338 , \49339 , \49340 ,
         \49341 , \49342 , \49343 , \49344 , \49345 , \49346 , \49347 , \49348 , \49349 , \49350 ,
         \49351 , \49352 , \49353 , \49354 , \49355 , \49356 , \49357 , \49358 , \49359 , \49360 ,
         \49361 , \49362 , \49363 , \49364 , \49365 , \49366 , \49367 , \49368 , \49369 , \49370 ,
         \49371 , \49372 , \49373 , \49374 , \49375 , \49376 , \49377 , \49378 , \49379 , \49380 ,
         \49381 , \49382 , \49383 , \49384 , \49385 , \49386 , \49387 , \49388 , \49389 , \49390 ,
         \49391 , \49392 , \49393 , \49394 , \49395 , \49396 , \49397 , \49398 , \49399 , \49400 ,
         \49401 , \49402 , \49403 , \49404 , \49405 , \49406 , \49407 , \49408 , \49409 , \49410 ,
         \49411 , \49412 , \49413 , \49414 , \49415 , \49416 , \49417 , \49418 , \49419 , \49420 ,
         \49421 , \49422 , \49423 , \49424 , \49425 , \49426 , \49427 , \49428 , \49429 , \49430 ,
         \49431 , \49432 , \49433 , \49434 , \49435 , \49436 , \49437 , \49438 , \49439 , \49440 ,
         \49441 , \49442 , \49443 , \49444 , \49445 , \49446 , \49447 , \49448 , \49449 , \49450 ,
         \49451 , \49452 , \49453 , \49454 , \49455 , \49456 , \49457 , \49458 , \49459 , \49460 ,
         \49461 , \49462 , \49463 , \49464 , \49465 , \49466 , \49467 , \49468 , \49469 , \49470 ,
         \49471 , \49472 , \49473 , \49474 , \49475 , \49476 , \49477 , \49478 , \49479 , \49480 ,
         \49481 , \49482 , \49483 , \49484 , \49485 , \49486 , \49487 , \49488 , \49489 , \49490 ,
         \49491 , \49492 , \49493 , \49494 , \49495 , \49496 , \49497 , \49498 , \49499 , \49500 ,
         \49501 , \49502 , \49503 , \49504 , \49505 , \49506 , \49507 , \49508 , \49509 , \49510 ,
         \49511 , \49512 , \49513 , \49514 , \49515 , \49516 , \49517 , \49518 , \49519 , \49520 ,
         \49521 , \49522 , \49523 , \49524 , \49525 , \49526 , \49527 , \49528 , \49529 , \49530 ,
         \49531 , \49532 , \49533 , \49534 , \49535 , \49536 , \49537 , \49538 , \49539 , \49540 ,
         \49541 , \49542 , \49543 , \49544 , \49545 , \49546 , \49547 , \49548 , \49549 , \49550 ,
         \49551 , \49552 , \49553 , \49554 , \49555 , \49556 , \49557 , \49558 , \49559 , \49560 ,
         \49561 , \49562 , \49563 , \49564 , \49565 , \49566 , \49567 , \49568 , \49569 , \49570 ,
         \49571 , \49572 , \49573 , \49574 , \49575 , \49576 , \49577 , \49578 , \49579 , \49580 ,
         \49581 , \49582 , \49583 , \49584 , \49585 , \49586 , \49587 , \49588 , \49589 , \49590 ,
         \49591 , \49592 , \49593 , \49594 , \49595 , \49596 , \49597 , \49598 , \49599 , \49600 ,
         \49601 , \49602 , \49603 , \49604 , \49605 , \49606 , \49607 , \49608 , \49609 , \49610 ,
         \49611 , \49612 , \49613 , \49614 , \49615 , \49616 , \49617 , \49618 , \49619 , \49620 ,
         \49621 , \49622 , \49623 , \49624 , \49625 , \49626 , \49627 , \49628 , \49629 , \49630 ,
         \49631 , \49632 , \49633 , \49634 , \49635 , \49636 , \49637 , \49638 , \49639 , \49640 ,
         \49641 , \49642 , \49643 , \49644 , \49645 , \49646 , \49647 , \49648 , \49649 , \49650 ,
         \49651 , \49652 , \49653 , \49654 , \49655 , \49656 , \49657 , \49658 , \49659 , \49660 ,
         \49661 , \49662 , \49663 , \49664 , \49665 , \49666 , \49667 , \49668 , \49669 , \49670 ,
         \49671 , \49672 , \49673 , \49674 , \49675 , \49676 , \49677 , \49678 , \49679 , \49680 ,
         \49681 , \49682 , \49683 , \49684 , \49685 , \49686 , \49687 , \49688 , \49689 , \49690 ,
         \49691 , \49692 , \49693 , \49694 , \49695 , \49696 , \49697 , \49698 , \49699 , \49700 ,
         \49701 , \49702 , \49703 , \49704 , \49705 , \49706 , \49707 , \49708 , \49709 , \49710 ,
         \49711 , \49712 , \49713 , \49714 , \49715 , \49716 , \49717 , \49718 , \49719 , \49720 ,
         \49721 , \49722 , \49723 , \49724 , \49725 , \49726 , \49727 , \49728 , \49729 , \49730 ,
         \49731 , \49732 , \49733 , \49734 , \49735 , \49736 , \49737 , \49738 , \49739 , \49740 ,
         \49741 , \49742 , \49743 , \49744 , \49745 , \49746 , \49747 , \49748 , \49749 , \49750 ,
         \49751 , \49752 , \49753 , \49754 , \49755 , \49756 , \49757 , \49758 , \49759 , \49760 ,
         \49761 , \49762 , \49763 , \49764 , \49765 , \49766 , \49767 , \49768 , \49769 , \49770 ,
         \49771 , \49772 , \49773 , \49774 , \49775 , \49776 , \49777 , \49778 , \49779 , \49780 ,
         \49781 , \49782 , \49783 , \49784 , \49785 , \49786 , \49787 , \49788 , \49789 , \49790 ,
         \49791 , \49792 , \49793 , \49794 , \49795 , \49796 , \49797 , \49798 , \49799 , \49800 ,
         \49801 , \49802 , \49803 , \49804 , \49805 , \49806 , \49807 , \49808 , \49809 , \49810 ,
         \49811 , \49812 , \49813 , \49814 , \49815 , \49816 , \49817 , \49818 , \49819 , \49820 ,
         \49821 , \49822 , \49823 , \49824 , \49825 , \49826 , \49827 , \49828 , \49829 , \49830 ,
         \49831 , \49832 , \49833 , \49834 , \49835 , \49836 , \49837 , \49838 , \49839 , \49840 ,
         \49841 , \49842 , \49843 , \49844 , \49845 , \49846 , \49847 , \49848 , \49849 , \49850 ,
         \49851 , \49852 , \49853 , \49854 , \49855 , \49856 , \49857 , \49858 , \49859 , \49860 ,
         \49861 , \49862 , \49863 , \49864 , \49865 , \49866 , \49867 , \49868 , \49869 , \49870 ,
         \49871 , \49872 , \49873 , \49874 , \49875 , \49876 , \49877 , \49878 , \49879 , \49880 ,
         \49881 , \49882 , \49883 , \49884 , \49885 , \49886 , \49887 , \49888 , \49889 , \49890 ,
         \49891 , \49892 , \49893 , \49894 , \49895 , \49896 , \49897 , \49898 , \49899 , \49900 ,
         \49901 , \49902 , \49903 , \49904 , \49905 , \49906 , \49907 , \49908 , \49909 , \49910 ,
         \49911 , \49912 , \49913 , \49914 , \49915 , \49916 , \49917 , \49918 , \49919 , \49920 ,
         \49921 , \49922 , \49923 , \49924 , \49925 , \49926 , \49927 , \49928 , \49929 , \49930 ,
         \49931 , \49932 , \49933 , \49934 , \49935 , \49936 , \49937 , \49938 , \49939 , \49940 ,
         \49941 , \49942 , \49943 , \49944 , \49945 , \49946 , \49947 , \49948 , \49949 , \49950 ,
         \49951 , \49952 , \49953 , \49954 , \49955 , \49956 , \49957 , \49958 , \49959 , \49960 ,
         \49961 , \49962 , \49963 , \49964 , \49965 , \49966 , \49967 , \49968 , \49969 , \49970 ,
         \49971 , \49972 , \49973 , \49974 , \49975 , \49976 , \49977 , \49978 , \49979 , \49980 ,
         \49981 , \49982 , \49983 , \49984 , \49985 , \49986 , \49987 , \49988 , \49989 , \49990 ,
         \49991 , \49992 , \49993 , \49994 , \49995 , \49996 , \49997 , \49998 , \49999 , \50000 ,
         \50001 , \50002 , \50003 , \50004 , \50005 , \50006 , \50007 , \50008 , \50009 , \50010 ,
         \50011 , \50012 , \50013 , \50014 , \50015 , \50016 , \50017 , \50018 , \50019 , \50020 ,
         \50021 , \50022 , \50023 , \50024 , \50025 , \50026 , \50027 , \50028 , \50029 , \50030 ,
         \50031 , \50032 , \50033 , \50034 , \50035 , \50036 , \50037 , \50038 , \50039 , \50040 ,
         \50041 , \50042 , \50043 , \50044 , \50045 , \50046 , \50047 , \50048 , \50049 , \50050 ,
         \50051 , \50052 , \50053 , \50054 , \50055 , \50056 , \50057 , \50058 , \50059 , \50060 ,
         \50061 , \50062 , \50063 , \50064 , \50065 , \50066 , \50067 , \50068 , \50069 , \50070 ,
         \50071 , \50072 , \50073 , \50074 , \50075 , \50076 , \50077 , \50078 , \50079 , \50080 ,
         \50081 , \50082 , \50083 , \50084 , \50085 , \50086 , \50087 , \50088 , \50089 , \50090 ,
         \50091 , \50092 , \50093 , \50094 , \50095 , \50096 , \50097 , \50098 , \50099 , \50100 ,
         \50101 , \50102 , \50103 , \50104 , \50105 , \50106 , \50107 , \50108 , \50109 , \50110 ,
         \50111 , \50112 , \50113 , \50114 , \50115 , \50116 , \50117 , \50118 , \50119 , \50120 ,
         \50121 , \50122 , \50123 , \50124 , \50125 , \50126 , \50127 , \50128 , \50129 , \50130 ,
         \50131 , \50132 , \50133 , \50134 , \50135 , \50136 , \50137 , \50138 , \50139 , \50140 ,
         \50141 , \50142 , \50143 , \50144 , \50145 , \50146 , \50147 , \50148 , \50149 , \50150 ,
         \50151 , \50152 , \50153 , \50154 , \50155 , \50156 , \50157 , \50158 , \50159 , \50160 ,
         \50161 , \50162 , \50163 , \50164 , \50165 , \50166 , \50167 , \50168 , \50169 , \50170 ,
         \50171 , \50172 , \50173 , \50174 , \50175 , \50176 , \50177 , \50178 , \50179 , \50180 ,
         \50181 , \50182 , \50183 , \50184 , \50185 , \50186 , \50187 , \50188 , \50189 , \50190 ,
         \50191 , \50192 , \50193 , \50194 , \50195 , \50196 , \50197 , \50198 , \50199 , \50200 ,
         \50201 , \50202 , \50203 , \50204 , \50205 , \50206 , \50207 , \50208 , \50209 , \50210 ,
         \50211 , \50212 , \50213 , \50214 , \50215 , \50216 , \50217 , \50218 , \50219 , \50220 ,
         \50221 , \50222 , \50223 , \50224 , \50225 , \50226 , \50227 , \50228 , \50229 , \50230 ,
         \50231 , \50232 , \50233 , \50234 , \50235 , \50236 , \50237 , \50238 , \50239 , \50240 ,
         \50241 , \50242 , \50243 , \50244 , \50245 , \50246 , \50247 , \50248 , \50249 , \50250 ,
         \50251 , \50252 , \50253 , \50254 , \50255 , \50256 , \50257 , \50258 , \50259 , \50260 ,
         \50261 , \50262 , \50263 , \50264 , \50265 , \50266 , \50267 , \50268 , \50269 , \50270 ,
         \50271 , \50272 , \50273 , \50274 , \50275 , \50276 , \50277 , \50278 , \50279 , \50280 ,
         \50281 , \50282 , \50283 , \50284 , \50285 , \50286 , \50287 , \50288 , \50289 , \50290 ,
         \50291 , \50292 , \50293 , \50294 , \50295 , \50296 , \50297 , \50298 , \50299 , \50300 ,
         \50301 , \50302 , \50303 , \50304 , \50305 , \50306 , \50307 , \50308 , \50309 , \50310 ,
         \50311 , \50312 , \50313 , \50314 , \50315 , \50316 , \50317 , \50318 , \50319 , \50320 ,
         \50321 , \50322 , \50323 , \50324 , \50325 , \50326 , \50327 , \50328 , \50329 , \50330 ,
         \50331 , \50332 , \50333 , \50334 , \50335 , \50336 , \50337 , \50338 , \50339 , \50340 ,
         \50341 , \50342 , \50343 , \50344 , \50345 , \50346 , \50347 , \50348 , \50349 , \50350 ,
         \50351 , \50352 , \50353 , \50354 , \50355 , \50356 , \50357 , \50358 , \50359 , \50360 ,
         \50361 , \50362 , \50363 , \50364 , \50365 , \50366 , \50367 , \50368 , \50369 , \50370 ,
         \50371 , \50372 , \50373 , \50374 , \50375 , \50376 , \50377 , \50378 , \50379 , \50380 ,
         \50381 , \50382 , \50383 , \50384 , \50385 , \50386 , \50387 , \50388 , \50389 , \50390 ,
         \50391 , \50392 , \50393 , \50394 , \50395 , \50396 , \50397 , \50398 , \50399 , \50400 ,
         \50401 , \50402 , \50403 , \50404 , \50405 , \50406 , \50407 , \50408 , \50409 , \50410 ,
         \50411 , \50412 , \50413 , \50414 , \50415 , \50416 , \50417 , \50418 , \50419 , \50420 ,
         \50421 , \50422 , \50423 , \50424 , \50425 , \50426 , \50427 , \50428 , \50429 , \50430 ,
         \50431 , \50432 , \50433 , \50434 , \50435 , \50436 , \50437 , \50438 , \50439 , \50440 ,
         \50441 , \50442 , \50443 , \50444 , \50445 , \50446 , \50447 , \50448 , \50449 , \50450 ,
         \50451 , \50452 , \50453 , \50454 , \50455 , \50456 , \50457 , \50458 , \50459 , \50460 ,
         \50461 , \50462 , \50463 , \50464 , \50465 , \50466 , \50467 , \50468 , \50469 , \50470 ,
         \50471 , \50472 , \50473 , \50474 , \50475 , \50476 , \50477 , \50478 , \50479 , \50480 ,
         \50481 , \50482 , \50483 , \50484 , \50485 , \50486 , \50487 , \50488 , \50489 , \50490 ,
         \50491 , \50492 , \50493 , \50494 , \50495 , \50496 , \50497 , \50498 , \50499 , \50500 ,
         \50501 , \50502 , \50503 , \50504 , \50505 , \50506 , \50507 , \50508 , \50509 , \50510 ,
         \50511 , \50512 , \50513 , \50514 , \50515 , \50516 , \50517 , \50518 , \50519 , \50520 ,
         \50521 , \50522 , \50523 , \50524 , \50525 , \50526 , \50527 , \50528 , \50529 , \50530 ,
         \50531 , \50532 , \50533 , \50534 , \50535 , \50536 , \50537 , \50538 , \50539 , \50540 ,
         \50541 , \50542 , \50543 , \50544 , \50545 , \50546 , \50547 , \50548 , \50549 , \50550 ,
         \50551 , \50552 , \50553 , \50554 , \50555 , \50556 , \50557 , \50558 , \50559 , \50560 ,
         \50561 , \50562 , \50563 , \50564 , \50565 , \50566 , \50567 , \50568 , \50569 , \50570 ,
         \50571 , \50572 , \50573 , \50574 , \50575 , \50576 , \50577 , \50578 , \50579 , \50580 ,
         \50581 , \50582 , \50583 , \50584 , \50585 , \50586 , \50587 , \50588 , \50589 , \50590 ,
         \50591 , \50592 , \50593 , \50594 , \50595 , \50596 , \50597 , \50598 , \50599 , \50600 ,
         \50601 , \50602 , \50603 , \50604 , \50605 , \50606 , \50607 , \50608 , \50609 , \50610 ,
         \50611 , \50612 , \50613 , \50614 , \50615 , \50616 , \50617 , \50618 , \50619 , \50620 ,
         \50621 , \50622 , \50623 , \50624 , \50625 , \50626 , \50627 , \50628 , \50629 , \50630 ,
         \50631 , \50632 , \50633 , \50634 , \50635 , \50636 , \50637 , \50638 , \50639 , \50640 ,
         \50641 , \50642 , \50643 , \50644 , \50645 , \50646 , \50647 , \50648 , \50649 , \50650 ,
         \50651 , \50652 , \50653 , \50654 , \50655 , \50656 , \50657 , \50658 , \50659 , \50660 ,
         \50661 , \50662 , \50663 , \50664 , \50665 , \50666 , \50667 , \50668 , \50669 , \50670 ,
         \50671 , \50672 , \50673 , \50674 , \50675 , \50676 , \50677 , \50678 , \50679 , \50680 ,
         \50681 , \50682 , \50683 , \50684 , \50685 , \50686 , \50687 , \50688 , \50689 , \50690 ,
         \50691 , \50692 , \50693 , \50694 , \50695 , \50696 , \50697 , \50698 , \50699 , \50700 ,
         \50701 , \50702 , \50703 , \50704 , \50705 , \50706 , \50707 , \50708 , \50709 , \50710 ,
         \50711 , \50712 , \50713 , \50714 , \50715 , \50716 , \50717 , \50718 , \50719 , \50720 ,
         \50721 , \50722 , \50723 , \50724 , \50725 , \50726 , \50727 , \50728 , \50729 , \50730 ,
         \50731 , \50732 , \50733 , \50734 , \50735 , \50736 , \50737 , \50738 , \50739 , \50740 ,
         \50741 , \50742 , \50743 , \50744 , \50745 , \50746 , \50747 , \50748 , \50749 , \50750 ,
         \50751 , \50752 , \50753 , \50754 , \50755 , \50756 , \50757 , \50758 , \50759 , \50760 ,
         \50761 , \50762 , \50763 , \50764 , \50765 , \50766 , \50767 , \50768 , \50769 , \50770 ,
         \50771 , \50772 , \50773 , \50774 , \50775 , \50776 , \50777 , \50778 , \50779 , \50780 ,
         \50781 , \50782 , \50783 , \50784 , \50785 , \50786 , \50787 , \50788 , \50789 , \50790 ,
         \50791 , \50792 , \50793 , \50794 , \50795 , \50796 , \50797 , \50798 , \50799 , \50800 ,
         \50801 , \50802 , \50803 , \50804 , \50805 , \50806 , \50807 , \50808 , \50809 , \50810 ,
         \50811 , \50812 , \50813 , \50814 , \50815 , \50816 , \50817 , \50818 , \50819 , \50820 ,
         \50821 , \50822 , \50823 , \50824 , \50825 , \50826 , \50827 , \50828 , \50829 , \50830 ,
         \50831 , \50832 , \50833 , \50834 , \50835 , \50836 , \50837 , \50838 , \50839 , \50840 ,
         \50841 , \50842 , \50843 , \50844 , \50845 , \50846 , \50847 , \50848 , \50849 , \50850 ,
         \50851 , \50852 , \50853 , \50854 , \50855 , \50856 , \50857 , \50858 , \50859 , \50860 ,
         \50861 , \50862 , \50863 , \50864 , \50865 , \50866 , \50867 , \50868 , \50869 , \50870 ,
         \50871 , \50872 , \50873 , \50874 , \50875 , \50876 , \50877 , \50878 , \50879 , \50880 ,
         \50881 , \50882 , \50883 , \50884 , \50885 , \50886 , \50887 , \50888 , \50889 , \50890 ,
         \50891 , \50892 , \50893 , \50894 , \50895 , \50896 , \50897 , \50898 , \50899 , \50900 ,
         \50901 , \50902 , \50903 , \50904 , \50905 , \50906 , \50907 , \50908 , \50909 , \50910 ,
         \50911 , \50912 , \50913 , \50914 , \50915 , \50916 , \50917 , \50918 , \50919 , \50920 ,
         \50921 , \50922 , \50923 , \50924 , \50925 , \50926 , \50927 , \50928 , \50929 , \50930 ,
         \50931 , \50932 , \50933 , \50934 , \50935 , \50936 , \50937 , \50938 , \50939 , \50940 ,
         \50941 , \50942 , \50943 , \50944 , \50945 , \50946 , \50947 , \50948 , \50949 , \50950 ,
         \50951 , \50952 , \50953 , \50954 , \50955 , \50956 , \50957 , \50958 , \50959 , \50960 ,
         \50961 , \50962 , \50963 , \50964 , \50965 , \50966 , \50967 , \50968 , \50969 , \50970 ,
         \50971 , \50972 , \50973 , \50974 , \50975 , \50976 , \50977 , \50978 , \50979 , \50980 ,
         \50981 , \50982 , \50983 , \50984 , \50985 , \50986 , \50987 , \50988 , \50989 , \50990 ,
         \50991 , \50992 , \50993 , \50994 , \50995 , \50996 , \50997 , \50998 , \50999 , \51000 ,
         \51001 , \51002 , \51003 , \51004 , \51005 , \51006 , \51007 , \51008 , \51009 , \51010 ,
         \51011 , \51012 , \51013 , \51014 , \51015 , \51016 , \51017 , \51018 , \51019 , \51020 ,
         \51021 , \51022 , \51023 , \51024 , \51025 , \51026 , \51027 , \51028 , \51029 , \51030 ,
         \51031 , \51032 , \51033 , \51034 , \51035 , \51036 , \51037 , \51038 , \51039 , \51040 ,
         \51041 , \51042 , \51043 , \51044 , \51045 , \51046 , \51047 , \51048 , \51049 , \51050 ,
         \51051 , \51052 , \51053 , \51054 , \51055 , \51056 , \51057 , \51058 , \51059 , \51060 ,
         \51061 , \51062 , \51063 , \51064 , \51065 , \51066 , \51067 , \51068 , \51069 , \51070 ,
         \51071 , \51072 , \51073 , \51074 , \51075 , \51076 , \51077 , \51078 , \51079 , \51080 ,
         \51081 , \51082 , \51083 , \51084 , \51085 , \51086 , \51087 , \51088 , \51089 , \51090 ,
         \51091 , \51092 , \51093 , \51094 , \51095 , \51096 , \51097 , \51098 , \51099 , \51100 ,
         \51101 , \51102 , \51103 , \51104 , \51105 , \51106 , \51107 , \51108 , \51109 , \51110 ,
         \51111 , \51112 , \51113 , \51114 , \51115 , \51116 , \51117 , \51118 , \51119 , \51120 ,
         \51121 , \51122 , \51123 , \51124 , \51125 , \51126 , \51127 , \51128 , \51129 , \51130 ,
         \51131 , \51132 , \51133 , \51134 , \51135 , \51136 , \51137 , \51138 , \51139 , \51140 ,
         \51141 , \51142 , \51143 , \51144 , \51145 , \51146 , \51147 , \51148 , \51149 , \51150 ,
         \51151 , \51152 , \51153 , \51154 , \51155 , \51156 , \51157 , \51158 , \51159 , \51160 ,
         \51161 , \51162 , \51163 , \51164 , \51165 , \51166 , \51167 , \51168 , \51169 , \51170 ,
         \51171 , \51172 , \51173 , \51174 , \51175 , \51176 , \51177 , \51178 , \51179 , \51180 ,
         \51181 , \51182 , \51183 , \51184 , \51185 , \51186 , \51187 , \51188 , \51189 , \51190 ,
         \51191 , \51192 , \51193 , \51194 , \51195 , \51196 , \51197 , \51198 , \51199 , \51200 ,
         \51201 , \51202 , \51203 , \51204 , \51205 , \51206 , \51207 , \51208 , \51209 , \51210 ,
         \51211 , \51212 , \51213 , \51214 , \51215 , \51216 , \51217 , \51218 , \51219 , \51220 ,
         \51221 , \51222 , \51223 , \51224 , \51225 , \51226 , \51227 , \51228 , \51229 , \51230 ,
         \51231 , \51232 , \51233 , \51234 , \51235 , \51236 , \51237 , \51238 , \51239 , \51240 ,
         \51241 , \51242 , \51243 , \51244 , \51245 , \51246 , \51247 , \51248 , \51249 , \51250 ,
         \51251 , \51252 , \51253 , \51254 , \51255 , \51256 , \51257 , \51258 , \51259 , \51260 ,
         \51261 , \51262 , \51263 , \51264 , \51265 , \51266 , \51267 , \51268 , \51269 , \51270 ,
         \51271 , \51272 , \51273 , \51274 , \51275 , \51276 , \51277 , \51278 , \51279 , \51280 ,
         \51281 , \51282 , \51283 , \51284 , \51285 , \51286 , \51287 , \51288 , \51289 , \51290 ,
         \51291 , \51292 , \51293 , \51294 , \51295 , \51296 , \51297 , \51298 , \51299 , \51300 ,
         \51301 , \51302 , \51303 , \51304 , \51305 , \51306 , \51307 , \51308 , \51309 , \51310 ,
         \51311 , \51312 , \51313 , \51314 , \51315 , \51316 , \51317 , \51318 , \51319 , \51320 ,
         \51321 , \51322 , \51323 , \51324 , \51325 , \51326 , \51327 , \51328 , \51329 , \51330 ,
         \51331 , \51332 , \51333 , \51334 , \51335 , \51336 , \51337 , \51338 , \51339 , \51340 ,
         \51341 , \51342 , \51343 , \51344 , \51345 , \51346 , \51347 , \51348 , \51349 , \51350 ,
         \51351 , \51352 , \51353 , \51354 , \51355 , \51356 , \51357 , \51358 , \51359 , \51360 ,
         \51361 , \51362 , \51363 , \51364 , \51365 , \51366 , \51367 , \51368 , \51369 , \51370 ,
         \51371 , \51372 , \51373 , \51374 , \51375 , \51376 , \51377 , \51378 , \51379 , \51380 ,
         \51381 , \51382 , \51383 , \51384 , \51385 , \51386 , \51387 , \51388 , \51389 , \51390 ,
         \51391 , \51392 , \51393 , \51394 , \51395 , \51396 , \51397 , \51398 , \51399 , \51400 ,
         \51401 , \51402 , \51403 , \51404 , \51405 , \51406 , \51407 , \51408 , \51409 , \51410 ,
         \51411 , \51412 , \51413 , \51414 , \51415 , \51416 , \51417 , \51418 , \51419 , \51420 ,
         \51421 , \51422 , \51423 , \51424 , \51425 , \51426 , \51427 , \51428 , \51429 , \51430 ,
         \51431 , \51432 , \51433 , \51434 , \51435 , \51436 , \51437 , \51438 , \51439 , \51440 ,
         \51441 , \51442 , \51443 , \51444 , \51445 , \51446 , \51447 , \51448 , \51449 , \51450 ,
         \51451 , \51452 , \51453 , \51454 , \51455 , \51456 , \51457 , \51458 , \51459 , \51460 ,
         \51461 , \51462 , \51463 , \51464 , \51465 , \51466 , \51467 , \51468 , \51469 , \51470 ,
         \51471 , \51472 , \51473 , \51474 , \51475 , \51476 , \51477 , \51478 , \51479 , \51480 ,
         \51481 , \51482 , \51483 , \51484 , \51485 , \51486 , \51487 , \51488 , \51489 , \51490 ,
         \51491 , \51492 , \51493 , \51494 , \51495 , \51496 , \51497 , \51498 , \51499 , \51500 ,
         \51501 , \51502 , \51503 , \51504 , \51505 , \51506 , \51507 , \51508 , \51509 , \51510 ,
         \51511 , \51512 , \51513 , \51514 , \51515 , \51516 , \51517 , \51518 , \51519 , \51520 ,
         \51521 , \51522 , \51523 , \51524 , \51525 , \51526 , \51527 , \51528 , \51529 , \51530 ,
         \51531 , \51532 , \51533 , \51534 , \51535 , \51536 , \51537 , \51538 , \51539 , \51540 ,
         \51541 , \51542 , \51543 , \51544 , \51545 , \51546 , \51547 , \51548 , \51549 , \51550 ,
         \51551 , \51552 , \51553 , \51554 , \51555 , \51556 , \51557 , \51558 , \51559 , \51560 ,
         \51561 , \51562 , \51563 , \51564 , \51565 , \51566 , \51567 , \51568 , \51569 , \51570 ,
         \51571 , \51572 , \51573 , \51574 , \51575 , \51576 , \51577 , \51578 , \51579 , \51580 ,
         \51581 , \51582 , \51583 , \51584 , \51585 , \51586 , \51587 , \51588 , \51589 , \51590 ,
         \51591 , \51592 , \51593 , \51594 , \51595 , \51596 , \51597 , \51598 , \51599 , \51600 ,
         \51601 , \51602 , \51603 , \51604 , \51605 , \51606 , \51607 , \51608 , \51609 , \51610 ,
         \51611 , \51612 , \51613 , \51614 , \51615 , \51616 , \51617 , \51618 , \51619 , \51620 ,
         \51621 , \51622 , \51623 , \51624 , \51625 , \51626 , \51627 , \51628 , \51629 , \51630 ,
         \51631 , \51632 , \51633 , \51634 , \51635 , \51636 , \51637 , \51638 , \51639 , \51640 ,
         \51641 , \51642 , \51643 , \51644 , \51645 , \51646 , \51647 , \51648 , \51649 , \51650 ,
         \51651 , \51652 , \51653 , \51654 , \51655 , \51656 , \51657 , \51658 , \51659 , \51660 ,
         \51661 , \51662 , \51663 , \51664 , \51665 , \51666 , \51667 , \51668 , \51669 , \51670 ,
         \51671 , \51672 , \51673 , \51674 , \51675 , \51676 , \51677 , \51678 , \51679 , \51680 ,
         \51681 , \51682 , \51683 , \51684 , \51685 , \51686 , \51687 , \51688 , \51689 , \51690 ,
         \51691 , \51692 , \51693 , \51694 , \51695 , \51696 , \51697 , \51698 , \51699 , \51700 ,
         \51701 , \51702 , \51703 , \51704 , \51705 , \51706 , \51707 , \51708 , \51709 , \51710 ,
         \51711 , \51712 , \51713 , \51714 , \51715 , \51716 , \51717 , \51718 , \51719 , \51720 ,
         \51721 , \51722 , \51723 , \51724 , \51725 , \51726 , \51727 , \51728 , \51729 , \51730 ,
         \51731 , \51732 , \51733 , \51734 , \51735 , \51736 , \51737 , \51738 , \51739 , \51740 ,
         \51741 , \51742 , \51743 , \51744 , \51745 , \51746 , \51747 , \51748 , \51749 , \51750 ,
         \51751 , \51752 , \51753 , \51754 , \51755 , \51756 , \51757 , \51758 , \51759 , \51760 ,
         \51761 , \51762 , \51763 , \51764 , \51765 , \51766 , \51767 , \51768 , \51769 , \51770 ,
         \51771 , \51772 , \51773 , \51774 , \51775 , \51776 , \51777 , \51778 , \51779 , \51780 ,
         \51781 , \51782 , \51783 , \51784 , \51785 , \51786 , \51787 , \51788 , \51789 , \51790 ,
         \51791 , \51792 , \51793 , \51794 , \51795 , \51796 , \51797 , \51798 , \51799 , \51800 ,
         \51801 , \51802 , \51803 , \51804 , \51805 , \51806 , \51807 , \51808 , \51809 , \51810 ,
         \51811 , \51812 , \51813 , \51814 , \51815 , \51816 , \51817 , \51818 , \51819 , \51820 ,
         \51821 , \51822 , \51823 , \51824 , \51825 , \51826 , \51827 , \51828 , \51829 , \51830 ,
         \51831 , \51832 , \51833 , \51834 , \51835 , \51836 , \51837 , \51838 , \51839 , \51840 ,
         \51841 , \51842 , \51843 , \51844 , \51845 , \51846 , \51847 , \51848 , \51849 , \51850 ,
         \51851 , \51852 , \51853 , \51854 , \51855 , \51856 , \51857 , \51858 , \51859 , \51860 ,
         \51861 , \51862 , \51863 , \51864 , \51865 , \51866 , \51867 , \51868 , \51869 , \51870 ,
         \51871 , \51872 , \51873 , \51874 , \51875 , \51876 , \51877 , \51878 , \51879 , \51880 ,
         \51881 , \51882 , \51883 , \51884 , \51885 , \51886 , \51887 , \51888 , \51889 , \51890 ,
         \51891 , \51892 , \51893 , \51894 , \51895 , \51896 , \51897 , \51898 , \51899 , \51900 ,
         \51901 , \51902 , \51903 , \51904 , \51905 , \51906 , \51907 , \51908 , \51909 , \51910 ,
         \51911 , \51912 , \51913 , \51914 , \51915 , \51916 , \51917 , \51918 , \51919 , \51920 ,
         \51921 , \51922 , \51923 , \51924 , \51925 , \51926 , \51927 , \51928 , \51929 , \51930 ,
         \51931 , \51932 , \51933 , \51934 , \51935 , \51936 , \51937 , \51938 , \51939 , \51940 ,
         \51941 , \51942 , \51943 , \51944 , \51945 , \51946 , \51947 , \51948 , \51949 , \51950 ,
         \51951 , \51952 , \51953 , \51954 , \51955 , \51956 , \51957 , \51958 , \51959 , \51960 ,
         \51961 , \51962 , \51963 , \51964 , \51965 , \51966 , \51967 , \51968 , \51969 , \51970 ,
         \51971 , \51972 , \51973 , \51974 , \51975 , \51976 , \51977 , \51978 , \51979 , \51980 ,
         \51981 , \51982 , \51983 , \51984 , \51985 , \51986 , \51987 , \51988 , \51989 , \51990 ,
         \51991 , \51992 , \51993 , \51994 , \51995 , \51996 , \51997 , \51998 , \51999 , \52000 ,
         \52001 , \52002 , \52003 , \52004 , \52005 , \52006 , \52007 , \52008 , \52009 , \52010 ,
         \52011 , \52012 , \52013 , \52014 , \52015 , \52016 , \52017 , \52018 , \52019 , \52020 ,
         \52021 , \52022 , \52023 , \52024 , \52025 , \52026 , \52027 , \52028 , \52029 , \52030 ,
         \52031 , \52032 , \52033 , \52034 , \52035 , \52036 , \52037 , \52038 , \52039 , \52040 ,
         \52041 , \52042 , \52043 , \52044 , \52045 , \52046 , \52047 , \52048 , \52049 , \52050 ,
         \52051 , \52052 , \52053 , \52054 , \52055 , \52056 , \52057 , \52058 , \52059 , \52060 ,
         \52061 , \52062 , \52063 , \52064 , \52065 , \52066 , \52067 , \52068 , \52069 , \52070 ,
         \52071 , \52072 , \52073 , \52074 , \52075 , \52076 , \52077 , \52078 , \52079 , \52080 ,
         \52081 , \52082 , \52083 , \52084 , \52085 , \52086 , \52087 , \52088 , \52089 , \52090 ,
         \52091 , \52092 , \52093 , \52094 , \52095 , \52096 , \52097 , \52098 , \52099 , \52100 ,
         \52101 , \52102 , \52103 , \52104 , \52105 , \52106 , \52107 , \52108 , \52109 , \52110 ,
         \52111 , \52112 , \52113 , \52114 , \52115 , \52116 , \52117 , \52118 , \52119 , \52120 ,
         \52121 , \52122 , \52123 , \52124 , \52125 , \52126 , \52127 , \52128 , \52129 , \52130 ,
         \52131 , \52132 , \52133 , \52134 , \52135 , \52136 , \52137 , \52138 , \52139 , \52140 ,
         \52141 , \52142 , \52143 , \52144 , \52145 , \52146 , \52147 , \52148 , \52149 , \52150 ,
         \52151 , \52152 , \52153 , \52154 , \52155 , \52156 , \52157 , \52158 , \52159 , \52160 ,
         \52161 , \52162 , \52163 , \52164 , \52165 , \52166 , \52167 , \52168 , \52169 , \52170 ,
         \52171 , \52172 , \52173 , \52174 , \52175 , \52176 , \52177 , \52178 , \52179 , \52180 ,
         \52181 , \52182 , \52183 , \52184 , \52185 , \52186 , \52187 , \52188 , \52189 , \52190 ,
         \52191 , \52192 , \52193 , \52194 , \52195 , \52196 , \52197 , \52198 , \52199 , \52200 ,
         \52201 , \52202 , \52203 , \52204 , \52205 , \52206 , \52207 , \52208 , \52209 , \52210 ,
         \52211 , \52212 , \52213 , \52214 , \52215 , \52216 , \52217 , \52218 , \52219 , \52220 ,
         \52221 , \52222 , \52223 , \52224 , \52225 , \52226 , \52227 , \52228 , \52229 , \52230 ,
         \52231 , \52232 , \52233 , \52234 , \52235 , \52236 , \52237 , \52238 , \52239 , \52240 ,
         \52241 , \52242 , \52243 , \52244 , \52245 , \52246 , \52247 , \52248 , \52249 , \52250 ,
         \52251 , \52252 , \52253 , \52254 , \52255 , \52256 , \52257 , \52258 , \52259 , \52260 ,
         \52261 , \52262 , \52263 , \52264 , \52265 , \52266 , \52267 , \52268 , \52269 , \52270 ,
         \52271 , \52272 , \52273 , \52274 , \52275 , \52276 , \52277 , \52278 , \52279 , \52280 ,
         \52281 , \52282 , \52283 , \52284 , \52285 , \52286 , \52287 , \52288 , \52289 , \52290 ,
         \52291 , \52292 , \52293 , \52294 , \52295 , \52296 , \52297 , \52298 , \52299 , \52300 ,
         \52301 , \52302 , \52303 , \52304 , \52305 , \52306 , \52307 , \52308 , \52309 , \52310 ,
         \52311 , \52312 , \52313 , \52314 , \52315 , \52316 , \52317 , \52318 , \52319 , \52320 ,
         \52321 , \52322 , \52323 , \52324 , \52325 , \52326 , \52327 , \52328 , \52329 , \52330 ,
         \52331 , \52332 , \52333 , \52334 , \52335 , \52336 , \52337 , \52338 , \52339 , \52340 ,
         \52341 , \52342 , \52343 , \52344 , \52345 , \52346 , \52347 , \52348 , \52349 , \52350 ,
         \52351 , \52352 , \52353 , \52354 , \52355 , \52356 , \52357 , \52358 , \52359 , \52360 ,
         \52361 , \52362 , \52363 , \52364 , \52365 , \52366 , \52367 , \52368 , \52369 , \52370 ,
         \52371 , \52372 , \52373 , \52374 , \52375 , \52376 , \52377 , \52378 , \52379 , \52380 ,
         \52381 , \52382 , \52383 , \52384 , \52385 , \52386 , \52387 , \52388 , \52389 , \52390 ,
         \52391 , \52392 , \52393 , \52394 , \52395 , \52396 , \52397 , \52398 , \52399 , \52400 ,
         \52401 , \52402 , \52403 , \52404 , \52405 , \52406 , \52407 , \52408 , \52409 , \52410 ,
         \52411 , \52412 , \52413 , \52414 , \52415 , \52416 , \52417 , \52418 , \52419 , \52420 ,
         \52421 , \52422 , \52423 , \52424 , \52425 , \52426 , \52427 , \52428 , \52429 , \52430 ,
         \52431 , \52432 , \52433 , \52434 , \52435 , \52436 , \52437 , \52438 , \52439 , \52440 ,
         \52441 , \52442 , \52443 , \52444 , \52445 , \52446 , \52447 , \52448 , \52449 , \52450 ,
         \52451 , \52452 , \52453 , \52454 , \52455 , \52456 , \52457 , \52458 , \52459 , \52460 ,
         \52461 , \52462 , \52463 , \52464 , \52465 , \52466 , \52467 , \52468 , \52469 , \52470 ,
         \52471 , \52472 , \52473 , \52474 , \52475 , \52476 , \52477 , \52478 , \52479 , \52480 ,
         \52481 , \52482 , \52483 , \52484 , \52485 , \52486 , \52487 , \52488 , \52489 , \52490 ,
         \52491 , \52492 , \52493 , \52494 , \52495 , \52496 , \52497 , \52498 , \52499 , \52500 ,
         \52501 , \52502 , \52503 , \52504 , \52505 , \52506 , \52507 , \52508 , \52509 , \52510 ,
         \52511 , \52512 , \52513 , \52514 , \52515 , \52516 , \52517 , \52518 , \52519 , \52520 ,
         \52521 , \52522 , \52523 , \52524 , \52525 , \52526 , \52527 , \52528 , \52529 , \52530 ,
         \52531 , \52532 , \52533 , \52534 , \52535 , \52536 , \52537 , \52538 , \52539 , \52540 ,
         \52541 , \52542 , \52543 , \52544 , \52545 , \52546 , \52547 , \52548 , \52549 , \52550 ,
         \52551 , \52552 , \52553 , \52554 , \52555 , \52556 , \52557 , \52558 , \52559 , \52560 ,
         \52561 , \52562 , \52563 , \52564 , \52565 , \52566 , \52567 , \52568 , \52569 , \52570 ,
         \52571 , \52572 , \52573 , \52574 , \52575 , \52576 , \52577 , \52578 , \52579 , \52580 ,
         \52581 , \52582 , \52583 , \52584 , \52585 , \52586 , \52587 , \52588 , \52589 , \52590 ,
         \52591 , \52592 , \52593 , \52594 , \52595 , \52596 , \52597 , \52598 , \52599 , \52600 ,
         \52601 , \52602 , \52603 , \52604 , \52605 , \52606 , \52607 , \52608 , \52609 , \52610 ,
         \52611 , \52612 , \52613 , \52614 , \52615 , \52616 , \52617 , \52618 , \52619 , \52620 ,
         \52621 , \52622 , \52623 , \52624 , \52625 , \52626 , \52627 , \52628 , \52629 , \52630 ,
         \52631 , \52632 , \52633 , \52634 , \52635 , \52636 , \52637 , \52638 , \52639 , \52640 ,
         \52641 , \52642 , \52643 , \52644 , \52645 , \52646 , \52647 , \52648 , \52649 , \52650 ,
         \52651 , \52652 , \52653 , \52654 , \52655 , \52656 , \52657 , \52658 , \52659 , \52660 ,
         \52661 , \52662 , \52663 , \52664 , \52665 , \52666 , \52667 , \52668 , \52669 , \52670 ,
         \52671 , \52672 , \52673 , \52674 , \52675 , \52676 , \52677 , \52678 , \52679 , \52680 ,
         \52681 , \52682 , \52683 , \52684 , \52685 , \52686 , \52687 , \52688 , \52689 , \52690 ,
         \52691 , \52692 , \52693 , \52694 , \52695 , \52696 , \52697 , \52698 , \52699 , \52700 ,
         \52701 , \52702 , \52703 , \52704 , \52705 , \52706 , \52707 , \52708 , \52709 , \52710 ,
         \52711 , \52712 , \52713 , \52714 , \52715 , \52716 , \52717 , \52718 , \52719 , \52720 ,
         \52721 , \52722 , \52723 , \52724 , \52725 , \52726 , \52727 , \52728 , \52729 , \52730 ,
         \52731 , \52732 , \52733 , \52734 , \52735 , \52736 , \52737 , \52738 , \52739 , \52740 ,
         \52741 , \52742 , \52743 , \52744 , \52745 , \52746 , \52747 , \52748 , \52749 , \52750 ,
         \52751 , \52752 , \52753 , \52754 , \52755 , \52756 , \52757 , \52758 , \52759 , \52760 ,
         \52761 , \52762 , \52763 , \52764 , \52765 , \52766 , \52767 , \52768 , \52769 , \52770 ,
         \52771 , \52772 , \52773 , \52774 , \52775 , \52776 , \52777 , \52778 , \52779 , \52780 ,
         \52781 , \52782 , \52783 , \52784 , \52785 , \52786 , \52787 , \52788 , \52789 , \52790 ,
         \52791 , \52792 , \52793 , \52794 , \52795 , \52796 , \52797 , \52798 , \52799 , \52800 ,
         \52801 , \52802 , \52803 , \52804 , \52805 , \52806 , \52807 , \52808 , \52809 , \52810 ,
         \52811 , \52812 , \52813 , \52814 , \52815 , \52816 , \52817 , \52818 , \52819 , \52820 ,
         \52821 , \52822 , \52823 , \52824 , \52825 , \52826 , \52827 , \52828 , \52829 , \52830 ,
         \52831 , \52832 , \52833 , \52834 , \52835 , \52836 , \52837 , \52838 , \52839 , \52840 ,
         \52841 , \52842 , \52843 , \52844 , \52845 , \52846 , \52847 , \52848 , \52849 , \52850 ,
         \52851 , \52852 , \52853 , \52854 , \52855 , \52856 , \52857 , \52858 , \52859 , \52860 ,
         \52861 , \52862 , \52863 , \52864 , \52865 , \52866 , \52867 , \52868 , \52869 , \52870 ,
         \52871 , \52872 , \52873 , \52874 , \52875 , \52876 , \52877 , \52878 , \52879 , \52880 ,
         \52881 , \52882 , \52883 , \52884 , \52885 , \52886 , \52887 , \52888 , \52889 , \52890 ,
         \52891 , \52892 , \52893 , \52894 , \52895 , \52896 , \52897 , \52898 , \52899 , \52900 ,
         \52901 , \52902 , \52903 , \52904 , \52905 , \52906 , \52907 , \52908 , \52909 , \52910 ,
         \52911 , \52912 , \52913 , \52914 , \52915 , \52916 , \52917 , \52918 , \52919 , \52920 ,
         \52921 , \52922 , \52923 , \52924 , \52925 , \52926 , \52927 , \52928 , \52929 , \52930 ,
         \52931 , \52932 , \52933 , \52934 , \52935 , \52936 , \52937 , \52938 , \52939 , \52940 ,
         \52941 , \52942 , \52943 , \52944 , \52945 , \52946 , \52947 , \52948 , \52949 , \52950 ,
         \52951 , \52952 , \52953 , \52954 , \52955 , \52956 , \52957 , \52958 , \52959 , \52960 ,
         \52961 , \52962 , \52963 , \52964 , \52965 , \52966 , \52967 , \52968 , \52969 , \52970 ,
         \52971 , \52972 , \52973 , \52974 , \52975 , \52976 , \52977 , \52978 , \52979 , \52980 ,
         \52981 , \52982 , \52983 , \52984 , \52985 , \52986 , \52987 , \52988 , \52989 , \52990 ,
         \52991 , \52992 , \52993 , \52994 , \52995 , \52996 , \52997 , \52998 , \52999 , \53000 ,
         \53001 , \53002 , \53003 , \53004 , \53005 , \53006 , \53007 , \53008 , \53009 , \53010 ,
         \53011 , \53012 , \53013 , \53014 , \53015 , \53016 , \53017 , \53018 , \53019 , \53020 ,
         \53021 , \53022 , \53023 , \53024 , \53025 , \53026 , \53027 , \53028 , \53029 , \53030 ,
         \53031 , \53032 , \53033 , \53034 , \53035 , \53036 , \53037 , \53038 , \53039 , \53040 ,
         \53041 , \53042 , \53043 , \53044 , \53045 , \53046 , \53047 , \53048 , \53049 , \53050 ,
         \53051 , \53052 , \53053 , \53054 , \53055 , \53056 , \53057 , \53058 , \53059 , \53060 ,
         \53061 , \53062 , \53063 , \53064 , \53065 , \53066 , \53067 , \53068 , \53069 , \53070 ,
         \53071 , \53072 , \53073 , \53074 , \53075 , \53076 , \53077 , \53078 , \53079 , \53080 ,
         \53081 , \53082 , \53083 , \53084 , \53085 , \53086 , \53087 , \53088 , \53089 , \53090 ,
         \53091 , \53092 , \53093 , \53094 , \53095 , \53096 , \53097 , \53098 , \53099 , \53100 ,
         \53101 , \53102 , \53103 , \53104 , \53105 , \53106 , \53107 , \53108 , \53109 , \53110 ,
         \53111 , \53112 , \53113 , \53114 , \53115 , \53116 , \53117 , \53118 , \53119 , \53120 ,
         \53121 , \53122 , \53123 , \53124 , \53125 , \53126 , \53127 , \53128 , \53129 , \53130 ,
         \53131 , \53132 , \53133 , \53134 , \53135 , \53136 , \53137 , \53138 , \53139 , \53140 ,
         \53141 , \53142 , \53143 , \53144 , \53145 , \53146 , \53147 , \53148 , \53149 , \53150 ,
         \53151 , \53152 , \53153 , \53154 , \53155 , \53156 , \53157 , \53158 , \53159 , \53160 ,
         \53161 , \53162 , \53163 , \53164 , \53165 , \53166 , \53167 , \53168 , \53169 , \53170 ,
         \53171 , \53172 , \53173 , \53174 , \53175 , \53176 , \53177 , \53178 , \53179 , \53180 ,
         \53181 , \53182 , \53183 , \53184 , \53185 , \53186 , \53187 , \53188 , \53189 , \53190 ,
         \53191 , \53192 , \53193 , \53194 , \53195 , \53196 , \53197 , \53198 , \53199 , \53200 ,
         \53201 , \53202 , \53203 , \53204 , \53205 , \53206 , \53207 , \53208 , \53209 , \53210 ,
         \53211 , \53212 , \53213 , \53214 , \53215 , \53216 , \53217 , \53218 , \53219 , \53220 ,
         \53221 , \53222 , \53223 , \53224 , \53225 , \53226 , \53227 , \53228 , \53229 , \53230 ,
         \53231 , \53232 , \53233 , \53234 , \53235 , \53236 , \53237 , \53238 , \53239 , \53240 ,
         \53241 , \53242 , \53243 , \53244 , \53245 , \53246 , \53247 , \53248 , \53249 , \53250 ,
         \53251 , \53252 , \53253 , \53254 , \53255 , \53256 , \53257 , \53258 , \53259 , \53260 ,
         \53261 , \53262 , \53263 , \53264 , \53265 , \53266 , \53267 , \53268 , \53269 , \53270 ,
         \53271 , \53272 , \53273 , \53274 , \53275 , \53276 , \53277 , \53278 , \53279 , \53280 ,
         \53281 , \53282 , \53283 , \53284 , \53285 , \53286 , \53287 , \53288 , \53289 , \53290 ,
         \53291 , \53292 , \53293 , \53294 , \53295 , \53296 , \53297 , \53298 , \53299 , \53300 ,
         \53301 , \53302 , \53303 , \53304 , \53305 , \53306 , \53307 , \53308 , \53309 , \53310 ,
         \53311 , \53312 , \53313 , \53314 , \53315 , \53316 , \53317 , \53318 , \53319 , \53320 ,
         \53321 , \53322 , \53323 , \53324 , \53325 , \53326 , \53327 , \53328 , \53329 , \53330 ,
         \53331 , \53332 , \53333 , \53334 , \53335 , \53336 , \53337 , \53338 , \53339 , \53340 ,
         \53341 , \53342 , \53343 , \53344 , \53345 , \53346 , \53347 , \53348 , \53349 , \53350 ,
         \53351 , \53352 , \53353 , \53354 , \53355 , \53356 , \53357 , \53358 , \53359 , \53360 ,
         \53361 , \53362 , \53363 , \53364 , \53365 , \53366 , \53367 , \53368 , \53369 , \53370 ,
         \53371 , \53372 , \53373 , \53374 , \53375 , \53376 , \53377 , \53378 , \53379 , \53380 ,
         \53381 , \53382 , \53383 , \53384 , \53385 , \53386 , \53387 , \53388 , \53389 , \53390 ,
         \53391 , \53392 , \53393 , \53394 , \53395 , \53396 , \53397 , \53398 , \53399 , \53400 ,
         \53401 , \53402 , \53403 , \53404 , \53405 , \53406 , \53407 , \53408 , \53409 , \53410 ,
         \53411 , \53412 , \53413 , \53414 , \53415 , \53416 , \53417 , \53418 , \53419 , \53420 ,
         \53421 , \53422 , \53423 , \53424 , \53425 , \53426 , \53427 , \53428 , \53429 , \53430 ,
         \53431 , \53432 , \53433 , \53434 , \53435 , \53436 , \53437 , \53438 , \53439 , \53440 ,
         \53441 , \53442 , \53443 , \53444 , \53445 , \53446 , \53447 , \53448 , \53449 , \53450 ,
         \53451 , \53452 , \53453 , \53454 , \53455 , \53456 , \53457 , \53458 , \53459 , \53460 ,
         \53461 , \53462 , \53463 , \53464 , \53465 , \53466 , \53467 , \53468 , \53469 , \53470 ,
         \53471 , \53472 , \53473 , \53474 , \53475 , \53476 , \53477 , \53478 , \53479 , \53480 ,
         \53481 , \53482 , \53483 , \53484 , \53485 , \53486 , \53487 , \53488 , \53489 , \53490 ,
         \53491 , \53492 , \53493 , \53494 , \53495 , \53496 , \53497 , \53498 , \53499 , \53500 ,
         \53501 , \53502 , \53503 , \53504 , \53505 , \53506 , \53507 , \53508 , \53509 , \53510 ,
         \53511 , \53512 , \53513 , \53514 , \53515 , \53516 , \53517 , \53518 , \53519 , \53520 ,
         \53521 , \53522 , \53523 , \53524 , \53525 , \53526 , \53527 , \53528 , \53529 , \53530 ,
         \53531 , \53532 , \53533 , \53534 , \53535 , \53536 , \53537 , \53538 , \53539 , \53540 ,
         \53541 , \53542 , \53543 , \53544 , \53545 , \53546 , \53547 , \53548 , \53549 , \53550 ,
         \53551 , \53552 , \53553 , \53554 , \53555 , \53556 , \53557 , \53558 , \53559 , \53560 ,
         \53561 , \53562 , \53563 , \53564 , \53565 , \53566 , \53567 , \53568 , \53569 , \53570 ,
         \53571 , \53572 , \53573 , \53574 , \53575 , \53576 , \53577 , \53578 , \53579 , \53580 ,
         \53581 , \53582 , \53583 , \53584 , \53585 , \53586 , \53587 , \53588 , \53589 , \53590 ,
         \53591 , \53592 , \53593 , \53594 , \53595 , \53596 , \53597 , \53598 , \53599 , \53600 ,
         \53601 , \53602 , \53603 , \53604 , \53605 , \53606 , \53607 , \53608 , \53609 , \53610 ,
         \53611 , \53612 , \53613 , \53614 , \53615 , \53616 , \53617 , \53618 , \53619 , \53620 ,
         \53621 , \53622 , \53623 , \53624 , \53625 , \53626 , \53627 , \53628 , \53629 , \53630 ,
         \53631 , \53632 , \53633 , \53634 , \53635 , \53636 , \53637 , \53638 , \53639 , \53640 ,
         \53641 , \53642 , \53643 , \53644 , \53645 , \53646 , \53647 , \53648 , \53649 , \53650 ,
         \53651 , \53652 , \53653 , \53654 , \53655 , \53656 , \53657 , \53658 , \53659 , \53660 ,
         \53661 , \53662 , \53663 , \53664 , \53665 , \53666 , \53667 , \53668 , \53669 , \53670 ,
         \53671 , \53672 , \53673 , \53674 , \53675 , \53676 , \53677 , \53678 , \53679 , \53680 ,
         \53681 , \53682 , \53683 , \53684 , \53685 , \53686 , \53687 , \53688 , \53689 , \53690 ,
         \53691 , \53692 , \53693 , \53694 , \53695 , \53696 , \53697 , \53698 , \53699 , \53700 ,
         \53701 , \53702 , \53703 , \53704 , \53705 , \53706 , \53707 , \53708 , \53709 , \53710 ,
         \53711 , \53712 , \53713 , \53714 , \53715 , \53716 , \53717 , \53718 , \53719 , \53720 ,
         \53721 , \53722 , \53723 , \53724 , \53725 , \53726 , \53727 , \53728 , \53729 , \53730 ,
         \53731 , \53732 , \53733 , \53734 , \53735 , \53736 , \53737 , \53738 , \53739 , \53740 ,
         \53741 , \53742 , \53743 , \53744 , \53745 , \53746 , \53747 , \53748 , \53749 , \53750 ,
         \53751 , \53752 , \53753 , \53754 , \53755 , \53756 , \53757 , \53758 , \53759 , \53760 ,
         \53761 , \53762 , \53763 , \53764 , \53765 , \53766 , \53767 , \53768 , \53769 , \53770 ,
         \53771 , \53772 , \53773 , \53774 , \53775 , \53776 , \53777 , \53778 , \53779 , \53780 ,
         \53781 , \53782 , \53783 , \53784 , \53785 , \53786 , \53787 , \53788 , \53789 , \53790 ,
         \53791 , \53792 , \53793 , \53794 , \53795 , \53796 , \53797 , \53798 , \53799 , \53800 ,
         \53801 , \53802 , \53803 , \53804 , \53805 , \53806 , \53807 , \53808 , \53809 , \53810 ,
         \53811 , \53812 , \53813 , \53814 , \53815 , \53816 , \53817 , \53818 , \53819 , \53820 ,
         \53821 , \53822 , \53823 , \53824 , \53825 , \53826 , \53827 , \53828 , \53829 , \53830 ,
         \53831 , \53832 , \53833 , \53834 , \53835 , \53836 , \53837 , \53838 , \53839 , \53840 ,
         \53841 , \53842 , \53843 , \53844 , \53845 , \53846 , \53847 , \53848 , \53849 , \53850 ,
         \53851 , \53852 , \53853 , \53854 , \53855 , \53856 , \53857 , \53858 , \53859 , \53860 ,
         \53861 , \53862 , \53863 , \53864 , \53865 , \53866 , \53867 , \53868 , \53869 , \53870 ,
         \53871 , \53872 , \53873 , \53874 , \53875 , \53876 , \53877 , \53878 , \53879 , \53880 ,
         \53881 , \53882 , \53883 , \53884 , \53885 , \53886 , \53887 , \53888 , \53889 , \53890 ,
         \53891 , \53892 , \53893 , \53894 , \53895 , \53896 , \53897 , \53898 , \53899 , \53900 ,
         \53901 , \53902 , \53903 , \53904 , \53905 , \53906 , \53907 , \53908 , \53909 , \53910 ,
         \53911 , \53912 , \53913 , \53914 , \53915 , \53916 , \53917 , \53918 , \53919 , \53920 ,
         \53921 , \53922 , \53923 , \53924 , \53925 , \53926 , \53927 , \53928 , \53929 , \53930 ,
         \53931 , \53932 , \53933 , \53934 , \53935 , \53936 , \53937 , \53938 , \53939 , \53940 ,
         \53941 , \53942 , \53943 , \53944 , \53945 , \53946 , \53947 , \53948 , \53949 , \53950 ,
         \53951 , \53952 , \53953 , \53954 , \53955 , \53956 , \53957 , \53958 , \53959 , \53960 ,
         \53961 , \53962 , \53963 , \53964 , \53965 , \53966 , \53967 , \53968 , \53969 , \53970 ,
         \53971 , \53972 , \53973 , \53974 , \53975 , \53976 , \53977 , \53978 , \53979 , \53980 ,
         \53981 , \53982 , \53983 , \53984 , \53985 , \53986 , \53987 , \53988 , \53989 , \53990 ,
         \53991 , \53992 , \53993 , \53994 , \53995 , \53996 , \53997 , \53998 , \53999 , \54000 ,
         \54001 , \54002 , \54003 , \54004 , \54005 , \54006 , \54007 , \54008 , \54009 , \54010 ,
         \54011 , \54012 , \54013 , \54014 , \54015 , \54016 , \54017 , \54018 , \54019 , \54020 ,
         \54021 , \54022 , \54023 , \54024 , \54025 , \54026 , \54027 , \54028 , \54029 , \54030 ,
         \54031 , \54032 , \54033 , \54034 , \54035 , \54036 , \54037 , \54038 , \54039 , \54040 ,
         \54041 , \54042 , \54043 , \54044 , \54045 , \54046 , \54047 , \54048 , \54049 , \54050 ,
         \54051 , \54052 , \54053 , \54054 , \54055 , \54056 , \54057 , \54058 , \54059 , \54060 ,
         \54061 , \54062 , \54063 , \54064 , \54065 , \54066 , \54067 , \54068 , \54069 , \54070 ,
         \54071 , \54072 , \54073 , \54074 , \54075 , \54076 , \54077 , \54078 , \54079 , \54080 ,
         \54081 , \54082 , \54083 , \54084 , \54085 , \54086 , \54087 , \54088 , \54089 , \54090 ,
         \54091 , \54092 , \54093 , \54094 , \54095 , \54096 , \54097 , \54098 , \54099 , \54100 ,
         \54101 , \54102 , \54103 , \54104 , \54105 , \54106 , \54107 , \54108 , \54109 , \54110 ,
         \54111 , \54112 , \54113 , \54114 , \54115 , \54116 , \54117 , \54118 , \54119 , \54120 ,
         \54121 , \54122 , \54123 , \54124 , \54125 , \54126 , \54127 , \54128 , \54129 , \54130 ,
         \54131 , \54132 , \54133 , \54134 , \54135 , \54136 , \54137 , \54138 , \54139 , \54140 ,
         \54141 , \54142 , \54143 , \54144 , \54145 , \54146 , \54147 , \54148 , \54149 , \54150 ,
         \54151 , \54152 , \54153 , \54154 , \54155 , \54156 , \54157 , \54158 , \54159 , \54160 ,
         \54161 , \54162 , \54163 , \54164 , \54165 , \54166 , \54167 , \54168 , \54169 , \54170 ,
         \54171 , \54172 , \54173 , \54174 , \54175 , \54176 , \54177 , \54178 , \54179 , \54180 ,
         \54181 , \54182 , \54183 , \54184 , \54185 , \54186 , \54187 , \54188 , \54189 , \54190 ,
         \54191 , \54192 , \54193 , \54194 , \54195 , \54196 , \54197 , \54198 , \54199 , \54200 ,
         \54201 , \54202 , \54203 , \54204 , \54205 , \54206 , \54207 , \54208 , \54209 , \54210 ,
         \54211 , \54212 , \54213 , \54214 , \54215 , \54216 , \54217 , \54218 , \54219 , \54220 ,
         \54221 , \54222 , \54223 , \54224 , \54225 , \54226 , \54227 , \54228 , \54229 , \54230 ,
         \54231 , \54232 , \54233 , \54234 , \54235 , \54236 , \54237 , \54238 , \54239 , \54240 ,
         \54241 , \54242 , \54243 , \54244 , \54245 , \54246 , \54247 , \54248 , \54249 , \54250 ,
         \54251 , \54252 , \54253 , \54254 , \54255 , \54256 , \54257 , \54258 , \54259 , \54260 ,
         \54261 , \54262 , \54263 , \54264 , \54265 , \54266 , \54267 , \54268 , \54269 , \54270 ,
         \54271 , \54272 , \54273 , \54274 , \54275 , \54276 , \54277 , \54278 , \54279 , \54280 ,
         \54281 , \54282 , \54283 , \54284 , \54285 , \54286 , \54287 , \54288 , \54289 , \54290 ,
         \54291 , \54292 , \54293 , \54294 , \54295 , \54296 , \54297 , \54298 , \54299 , \54300 ,
         \54301 , \54302 , \54303 , \54304 , \54305 , \54306 , \54307 , \54308 , \54309 , \54310 ,
         \54311 , \54312 , \54313 , \54314 , \54315 , \54316 , \54317 , \54318 , \54319 , \54320 ,
         \54321 , \54322 , \54323 , \54324 , \54325 , \54326 , \54327 , \54328 , \54329 , \54330 ,
         \54331 , \54332 , \54333 , \54334 , \54335 , \54336 , \54337 , \54338 , \54339 , \54340 ,
         \54341 , \54342 , \54343 , \54344 , \54345 , \54346 , \54347 , \54348 , \54349 , \54350 ,
         \54351 , \54352 , \54353 , \54354 , \54355 , \54356 , \54357 , \54358 , \54359 , \54360 ,
         \54361 , \54362 , \54363 , \54364 , \54365 , \54366 , \54367 , \54368 , \54369 , \54370 ,
         \54371 , \54372 , \54373 , \54374 , \54375 , \54376 , \54377 , \54378 , \54379 , \54380 ,
         \54381 , \54382 , \54383 , \54384 , \54385 , \54386 , \54387 , \54388 , \54389 , \54390 ,
         \54391 , \54392 , \54393 , \54394 , \54395 , \54396 , \54397 , \54398 , \54399 , \54400 ,
         \54401 , \54402 , \54403 , \54404 , \54405 , \54406 , \54407 , \54408 , \54409 , \54410 ,
         \54411 , \54412 , \54413 , \54414 , \54415 , \54416 , \54417 , \54418 , \54419 , \54420 ,
         \54421 , \54422 , \54423 , \54424 , \54425 , \54426 , \54427 , \54428 , \54429 , \54430 ,
         \54431 , \54432 , \54433 , \54434 , \54435 , \54436 , \54437 , \54438 , \54439 , \54440 ,
         \54441 , \54442 , \54443 , \54444 , \54445 , \54446 , \54447 , \54448 , \54449 , \54450 ,
         \54451 , \54452 , \54453 , \54454 , \54455 , \54456 , \54457 , \54458 , \54459 , \54460 ,
         \54461 , \54462 , \54463 , \54464 , \54465 , \54466 , \54467 , \54468 , \54469 , \54470 ,
         \54471 , \54472 , \54473 , \54474 , \54475 , \54476 , \54477 , \54478 , \54479 , \54480 ,
         \54481 , \54482 , \54483 , \54484 , \54485 , \54486 , \54487 , \54488 , \54489 , \54490 ,
         \54491 , \54492 , \54493 , \54494 , \54495 , \54496 , \54497 , \54498 , \54499 , \54500 ,
         \54501 , \54502 , \54503 , \54504 , \54505 , \54506 , \54507 , \54508 , \54509 , \54510 ,
         \54511 , \54512 , \54513 , \54514 , \54515 , \54516 , \54517 , \54518 , \54519 , \54520 ,
         \54521 , \54522 , \54523 , \54524 , \54525 , \54526 , \54527 , \54528 , \54529 , \54530 ,
         \54531 , \54532 , \54533 , \54534 , \54535 , \54536 , \54537 , \54538 , \54539 , \54540 ,
         \54541 , \54542 , \54543 , \54544 , \54545 , \54546 , \54547 , \54548 , \54549 , \54550 ,
         \54551 , \54552 , \54553 , \54554 , \54555 , \54556 , \54557 , \54558 , \54559 , \54560 ,
         \54561 , \54562 , \54563 , \54564 , \54565 , \54566 , \54567 , \54568 , \54569 , \54570 ,
         \54571 , \54572 , \54573 , \54574 , \54575 , \54576 , \54577 , \54578 , \54579 , \54580 ,
         \54581 , \54582 , \54583 , \54584 , \54585 , \54586 , \54587 , \54588 , \54589 , \54590 ,
         \54591 , \54592 , \54593 , \54594 , \54595 , \54596 , \54597 , \54598 , \54599 , \54600 ,
         \54601 , \54602 , \54603 , \54604 , \54605 , \54606 , \54607 , \54608 , \54609 , \54610 ,
         \54611 , \54612 , \54613 , \54614 , \54615 , \54616 , \54617 , \54618 , \54619 , \54620 ,
         \54621 , \54622 , \54623 , \54624 , \54625 , \54626 , \54627 , \54628 , \54629 , \54630 ,
         \54631 , \54632 , \54633 , \54634 , \54635 , \54636 , \54637 , \54638 , \54639 , \54640 ,
         \54641 , \54642 , \54643 , \54644 , \54645 , \54646 , \54647 , \54648 , \54649 , \54650 ,
         \54651 , \54652 , \54653 , \54654 , \54655 , \54656 , \54657 , \54658 , \54659 , \54660 ,
         \54661 , \54662 , \54663 , \54664 , \54665 , \54666 , \54667 , \54668 , \54669 , \54670 ,
         \54671 , \54672 , \54673 , \54674 , \54675 , \54676 , \54677 , \54678 , \54679 , \54680 ,
         \54681 , \54682 , \54683 , \54684 , \54685 , \54686 , \54687 , \54688 , \54689 , \54690 ,
         \54691 , \54692 , \54693 , \54694 , \54695 , \54696 , \54697 , \54698 , \54699 , \54700 ,
         \54701 , \54702 , \54703 , \54704 , \54705 , \54706 , \54707 , \54708 , \54709 , \54710 ,
         \54711 , \54712 , \54713 , \54714 , \54715 , \54716 , \54717 , \54718 , \54719 , \54720 ,
         \54721 , \54722 , \54723 , \54724 , \54725 , \54726 , \54727 , \54728 , \54729 , \54730 ,
         \54731 , \54732 , \54733 , \54734 , \54735 , \54736 , \54737 , \54738 , \54739 , \54740 ,
         \54741 , \54742 , \54743 , \54744 , \54745 , \54746 , \54747 , \54748 , \54749 , \54750 ,
         \54751 , \54752 , \54753 , \54754 , \54755 , \54756 , \54757 , \54758 , \54759 , \54760 ,
         \54761 , \54762 , \54763 , \54764 , \54765 , \54766 , \54767 , \54768 , \54769 , \54770 ,
         \54771 , \54772 , \54773 , \54774 , \54775 , \54776 , \54777 , \54778 , \54779 , \54780 ,
         \54781 , \54782 , \54783 , \54784 , \54785 , \54786 , \54787 , \54788 , \54789 , \54790 ,
         \54791 , \54792 , \54793 , \54794 , \54795 , \54796 , \54797 , \54798 , \54799 , \54800 ,
         \54801 , \54802 , \54803 , \54804 , \54805 , \54806 , \54807 , \54808 , \54809 , \54810 ,
         \54811 , \54812 , \54813 , \54814 , \54815 , \54816 , \54817 , \54818 , \54819 , \54820 ,
         \54821 , \54822 , \54823 , \54824 , \54825 , \54826 , \54827 , \54828 , \54829 , \54830 ,
         \54831 , \54832 , \54833 , \54834 , \54835 , \54836 , \54837 , \54838 , \54839 , \54840 ,
         \54841 , \54842 , \54843 , \54844 , \54845 , \54846 , \54847 , \54848 , \54849 , \54850 ,
         \54851 , \54852 , \54853 , \54854 , \54855 , \54856 , \54857 , \54858 , \54859 , \54860 ,
         \54861 , \54862 , \54863 , \54864 , \54865 , \54866 , \54867 , \54868 , \54869 , \54870 ,
         \54871 , \54872 , \54873 , \54874 , \54875 , \54876 , \54877 , \54878 , \54879 , \54880 ,
         \54881 , \54882 , \54883 , \54884 , \54885 , \54886 , \54887 , \54888 , \54889 , \54890 ,
         \54891 , \54892 , \54893 , \54894 , \54895 , \54896 , \54897 , \54898 , \54899 , \54900 ,
         \54901 , \54902 , \54903 , \54904 , \54905 , \54906 , \54907 , \54908 , \54909 , \54910 ,
         \54911 , \54912 , \54913 , \54914 , \54915 , \54916 , \54917 , \54918 , \54919 , \54920 ,
         \54921 , \54922 , \54923 , \54924 , \54925 , \54926 , \54927 , \54928 , \54929 , \54930 ,
         \54931 , \54932 , \54933 , \54934 , \54935 , \54936 , \54937 , \54938 , \54939 , \54940 ,
         \54941 , \54942 , \54943 , \54944 , \54945 , \54946 , \54947 , \54948 , \54949 , \54950 ,
         \54951 , \54952 , \54953 , \54954 , \54955 , \54956 , \54957 , \54958 , \54959 , \54960 ,
         \54961 , \54962 , \54963 , \54964 , \54965 , \54966 , \54967 , \54968 , \54969 , \54970 ,
         \54971 , \54972 , \54973 , \54974 , \54975 , \54976 , \54977 , \54978 , \54979 , \54980 ,
         \54981 , \54982 , \54983 , \54984 , \54985 , \54986 , \54987 , \54988 , \54989 , \54990 ,
         \54991 , \54992 , \54993 , \54994 , \54995 , \54996 , \54997 , \54998 , \54999 , \55000 ,
         \55001 , \55002 , \55003 , \55004 , \55005 , \55006 , \55007 , \55008 , \55009 , \55010 ,
         \55011 , \55012 , \55013 , \55014 , \55015 , \55016 , \55017 , \55018 , \55019 , \55020 ,
         \55021 , \55022 , \55023 , \55024 , \55025 , \55026 , \55027 , \55028 , \55029 , \55030 ,
         \55031 , \55032 , \55033 , \55034 , \55035 , \55036 , \55037 , \55038 , \55039 , \55040 ,
         \55041 , \55042 , \55043 , \55044 , \55045 , \55046 , \55047 , \55048 , \55049 , \55050 ,
         \55051 , \55052 , \55053 , \55054 , \55055 , \55056 , \55057 , \55058 , \55059 , \55060 ,
         \55061 , \55062 , \55063 , \55064 , \55065 , \55066 , \55067 , \55068 , \55069 , \55070 ,
         \55071 , \55072 , \55073 , \55074 , \55075 , \55076 , \55077 , \55078 , \55079 , \55080 ,
         \55081 , \55082 , \55083 , \55084 , \55085 , \55086 , \55087 , \55088 , \55089 , \55090 ,
         \55091 , \55092 , \55093 , \55094 , \55095 , \55096 , \55097 , \55098 , \55099 , \55100 ,
         \55101 , \55102 , \55103 , \55104 , \55105 , \55106 , \55107 , \55108 , \55109 , \55110 ,
         \55111 , \55112 , \55113 , \55114 , \55115 , \55116 , \55117 , \55118 , \55119 , \55120 ,
         \55121 , \55122 , \55123 , \55124 , \55125 , \55126 , \55127 , \55128 , \55129 , \55130 ,
         \55131 , \55132 , \55133 , \55134 , \55135 , \55136 , \55137 , \55138 , \55139 , \55140 ,
         \55141 , \55142 , \55143 , \55144 , \55145 , \55146 , \55147 , \55148 , \55149 , \55150 ,
         \55151 , \55152 , \55153 , \55154 , \55155 , \55156 , \55157 , \55158 , \55159 , \55160 ,
         \55161 , \55162 , \55163 , \55164 , \55165 , \55166 , \55167 , \55168 , \55169 , \55170 ,
         \55171 , \55172 , \55173 , \55174 , \55175 , \55176 , \55177 , \55178 , \55179 , \55180 ,
         \55181 , \55182 , \55183 , \55184 , \55185 , \55186 , \55187 , \55188 , \55189 , \55190 ,
         \55191 , \55192 , \55193 , \55194 , \55195 , \55196 , \55197 , \55198 , \55199 , \55200 ,
         \55201 , \55202 , \55203 , \55204 , \55205 , \55206 , \55207 , \55208 , \55209 , \55210 ,
         \55211 , \55212 , \55213 , \55214 , \55215 , \55216 , \55217 , \55218 , \55219 , \55220 ,
         \55221 , \55222 , \55223 , \55224 , \55225 , \55226 , \55227 , \55228 , \55229 , \55230 ,
         \55231 , \55232 , \55233 , \55234 , \55235 , \55236 , \55237 , \55238 , \55239 , \55240 ,
         \55241 , \55242 , \55243 , \55244 , \55245 , \55246 , \55247 , \55248 , \55249 , \55250 ,
         \55251 , \55252 , \55253 , \55254 , \55255 , \55256 , \55257 , \55258 , \55259 , \55260 ,
         \55261 , \55262 , \55263 , \55264 , \55265 , \55266 , \55267 , \55268 , \55269 , \55270 ,
         \55271 , \55272 , \55273 , \55274 , \55275 , \55276 , \55277 , \55278 , \55279 , \55280 ,
         \55281 , \55282 , \55283 , \55284 , \55285 , \55286 , \55287 , \55288 , \55289 , \55290 ,
         \55291 , \55292 , \55293 , \55294 , \55295 , \55296 , \55297 , \55298 , \55299 , \55300 ,
         \55301 , \55302 , \55303 , \55304 , \55305 , \55306 , \55307 , \55308 , \55309 , \55310 ,
         \55311 , \55312 , \55313 , \55314 , \55315 , \55316 , \55317 , \55318 , \55319 , \55320 ,
         \55321 , \55322 , \55323 , \55324 , \55325 , \55326 , \55327 , \55328 , \55329 , \55330 ,
         \55331 , \55332 , \55333 , \55334 , \55335 , \55336 , \55337 , \55338 , \55339 , \55340 ,
         \55341 , \55342 , \55343 , \55344 , \55345 , \55346 , \55347 , \55348 , \55349 , \55350 ,
         \55351 , \55352 , \55353 , \55354 , \55355 , \55356 , \55357 , \55358 , \55359 , \55360 ,
         \55361 , \55362 , \55363 , \55364 , \55365 , \55366 , \55367 , \55368 , \55369 , \55370 ,
         \55371 , \55372 , \55373 , \55374 , \55375 , \55376 , \55377 , \55378 , \55379 , \55380 ,
         \55381 , \55382 , \55383 , \55384 , \55385 , \55386 , \55387 , \55388 , \55389 , \55390 ,
         \55391 , \55392 , \55393 , \55394 , \55395 , \55396 , \55397 , \55398 , \55399 , \55400 ,
         \55401 , \55402 , \55403 , \55404 , \55405 , \55406 , \55407 , \55408 , \55409 , \55410 ,
         \55411 , \55412 , \55413 , \55414 , \55415 , \55416 , \55417 , \55418 , \55419 , \55420 ,
         \55421 , \55422 , \55423 , \55424 , \55425 , \55426 , \55427 , \55428 , \55429 , \55430 ,
         \55431 , \55432 , \55433 , \55434 , \55435 , \55436 , \55437 , \55438 , \55439 , \55440 ,
         \55441 , \55442 , \55443 , \55444 , \55445 , \55446 , \55447 , \55448 , \55449 , \55450 ,
         \55451 , \55452 , \55453 , \55454 , \55455 , \55456 , \55457 , \55458 , \55459 , \55460 ,
         \55461 , \55462 , \55463 , \55464 , \55465 , \55466 , \55467 , \55468 , \55469 , \55470 ,
         \55471 , \55472 , \55473 , \55474 , \55475 , \55476 , \55477 , \55478 , \55479 , \55480 ,
         \55481 , \55482 , \55483 , \55484 , \55485 , \55486 , \55487 , \55488 , \55489 , \55490 ,
         \55491 , \55492 , \55493 , \55494 , \55495 , \55496 , \55497 , \55498 , \55499 , \55500 ,
         \55501 , \55502 , \55503 , \55504 , \55505 , \55506 , \55507 , \55508 , \55509 , \55510 ,
         \55511 , \55512 , \55513 , \55514 , \55515 , \55516 , \55517 , \55518 , \55519 , \55520 ,
         \55521 , \55522 , \55523 , \55524 , \55525 , \55526 , \55527 , \55528 , \55529 , \55530 ,
         \55531 , \55532 , \55533 , \55534 , \55535 , \55536 , \55537 , \55538 , \55539 , \55540 ,
         \55541 , \55542 , \55543 , \55544 , \55545 , \55546 , \55547 , \55548 , \55549 , \55550 ,
         \55551 , \55552 , \55553 , \55554 , \55555 , \55556 , \55557 , \55558 , \55559 , \55560 ,
         \55561 , \55562 , \55563 , \55564 , \55565 , \55566 , \55567 , \55568 , \55569 , \55570 ,
         \55571 , \55572 , \55573 , \55574 , \55575 , \55576 , \55577 , \55578 , \55579 , \55580 ,
         \55581 , \55582 , \55583 , \55584 , \55585 , \55586 , \55587 , \55588 , \55589 , \55590 ,
         \55591 , \55592 , \55593 , \55594 , \55595 , \55596 , \55597 , \55598 , \55599 , \55600 ,
         \55601 , \55602 , \55603 , \55604 , \55605 , \55606 , \55607 , \55608 , \55609 , \55610 ,
         \55611 , \55612 , \55613 , \55614 , \55615 , \55616 , \55617 , \55618 , \55619 , \55620 ,
         \55621 , \55622 , \55623 , \55624 , \55625 , \55626 , \55627 , \55628 , \55629 , \55630 ,
         \55631 , \55632 , \55633 , \55634 , \55635 , \55636 , \55637 , \55638 , \55639 , \55640 ,
         \55641 , \55642 , \55643 , \55644 , \55645 , \55646 , \55647 , \55648 , \55649 , \55650 ,
         \55651 , \55652 , \55653 , \55654 , \55655 , \55656 , \55657 , \55658 , \55659 , \55660 ,
         \55661 , \55662 , \55663 , \55664 , \55665 , \55666 , \55667 , \55668 , \55669 , \55670 ,
         \55671 , \55672 , \55673 , \55674 , \55675 , \55676 , \55677 , \55678 , \55679 , \55680 ,
         \55681 , \55682 , \55683 , \55684 , \55685 , \55686 , \55687 , \55688 , \55689 , \55690 ,
         \55691 , \55692 , \55693 , \55694 , \55695 , \55696 , \55697 , \55698 , \55699 , \55700 ,
         \55701 , \55702 , \55703 , \55704 , \55705 , \55706 , \55707 , \55708 , \55709 , \55710 ,
         \55711 , \55712 , \55713 , \55714 , \55715 , \55716 , \55717 , \55718 , \55719 , \55720 ,
         \55721 , \55722 , \55723 , \55724 , \55725 , \55726 , \55727 , \55728 , \55729 , \55730 ,
         \55731 , \55732 , \55733 , \55734 , \55735 , \55736 , \55737 , \55738 , \55739 , \55740 ,
         \55741 , \55742 , \55743 , \55744 , \55745 , \55746 , \55747 , \55748 , \55749 , \55750 ,
         \55751 , \55752 , \55753 , \55754 , \55755 , \55756 , \55757 , \55758 , \55759 , \55760 ,
         \55761 , \55762 , \55763 , \55764 , \55765 , \55766 , \55767 , \55768 , \55769 , \55770 ,
         \55771 , \55772 , \55773 , \55774 , \55775 , \55776 , \55777 , \55778 , \55779 , \55780 ,
         \55781 , \55782 , \55783 , \55784 , \55785 , \55786 , \55787 , \55788 , \55789 , \55790 ,
         \55791 , \55792 , \55793 , \55794 , \55795 , \55796 , \55797 , \55798 , \55799 , \55800 ,
         \55801 , \55802 , \55803 , \55804 , \55805 , \55806 , \55807 , \55808 , \55809 , \55810 ,
         \55811 , \55812 , \55813 , \55814 , \55815 , \55816 , \55817 , \55818 , \55819 , \55820 ,
         \55821 , \55822 , \55823 , \55824 , \55825 , \55826 , \55827 , \55828 , \55829 , \55830 ,
         \55831 , \55832 , \55833 , \55834 , \55835 , \55836 , \55837 , \55838 , \55839 , \55840 ,
         \55841 , \55842 , \55843 , \55844 , \55845 , \55846 , \55847 , \55848 , \55849 , \55850 ,
         \55851 , \55852 , \55853 , \55854 , \55855 , \55856 , \55857 , \55858 , \55859 , \55860 ,
         \55861 , \55862 , \55863 , \55864 , \55865 , \55866 , \55867 , \55868 , \55869 , \55870 ,
         \55871 , \55872 , \55873 , \55874 , \55875 , \55876 , \55877 , \55878 , \55879 , \55880 ,
         \55881 , \55882 , \55883 , \55884 , \55885 , \55886 , \55887 , \55888 , \55889 , \55890 ,
         \55891 , \55892 , \55893 , \55894 , \55895 , \55896 , \55897 , \55898 , \55899 , \55900 ,
         \55901 , \55902 , \55903 , \55904 , \55905 , \55906 , \55907 , \55908 , \55909 , \55910 ,
         \55911 , \55912 , \55913 , \55914 , \55915 , \55916 , \55917 , \55918 , \55919 , \55920 ,
         \55921 , \55922 , \55923 , \55924 , \55925 , \55926 , \55927 , \55928 , \55929 , \55930 ,
         \55931 , \55932 , \55933 , \55934 , \55935 , \55936 , \55937 , \55938 , \55939 , \55940 ,
         \55941 , \55942 , \55943 , \55944 , \55945 , \55946 , \55947 , \55948 , \55949 , \55950 ,
         \55951 , \55952 , \55953 , \55954 , \55955 , \55956 , \55957 , \55958 , \55959 , \55960 ,
         \55961 , \55962 , \55963 , \55964 , \55965 , \55966 , \55967 , \55968 , \55969 , \55970 ,
         \55971 , \55972 , \55973 , \55974 , \55975 , \55976 , \55977 , \55978 , \55979 , \55980 ,
         \55981 , \55982 , \55983 , \55984 , \55985 , \55986 , \55987 , \55988 , \55989 , \55990 ,
         \55991 , \55992 , \55993 , \55994 , \55995 , \55996 , \55997 , \55998 , \55999 , \56000 ,
         \56001 , \56002 , \56003 , \56004 , \56005 , \56006 , \56007 , \56008 , \56009 , \56010 ,
         \56011 , \56012 , \56013 , \56014 , \56015 , \56016 , \56017 , \56018 , \56019 , \56020 ,
         \56021 , \56022 , \56023 , \56024 , \56025 , \56026 , \56027 , \56028 , \56029 , \56030 ,
         \56031 , \56032 , \56033 , \56034 , \56035 , \56036 , \56037 , \56038 , \56039 , \56040 ,
         \56041 , \56042 , \56043 , \56044 , \56045 , \56046 , \56047 , \56048 , \56049 , \56050 ,
         \56051 , \56052 , \56053 , \56054 , \56055 , \56056 , \56057 , \56058 , \56059 , \56060 ,
         \56061 , \56062 , \56063 , \56064 , \56065 , \56066 , \56067 , \56068 , \56069 , \56070 ,
         \56071 , \56072 , \56073 , \56074 , \56075 , \56076 , \56077 , \56078 , \56079 , \56080 ,
         \56081 , \56082 , \56083 , \56084 , \56085 , \56086 , \56087 , \56088 , \56089 , \56090 ,
         \56091 , \56092 , \56093 , \56094 , \56095 , \56096 , \56097 , \56098 , \56099 , \56100 ,
         \56101 , \56102 , \56103 , \56104 , \56105 , \56106 , \56107 , \56108 , \56109 , \56110 ,
         \56111 , \56112 , \56113 , \56114 , \56115 , \56116 , \56117 , \56118 , \56119 , \56120 ,
         \56121 , \56122 , \56123 , \56124 , \56125 , \56126 , \56127 , \56128 , \56129 , \56130 ,
         \56131 , \56132 , \56133 , \56134 , \56135 , \56136 , \56137 , \56138 , \56139 , \56140 ,
         \56141 , \56142 , \56143 , \56144 , \56145 , \56146 , \56147 , \56148 , \56149 , \56150 ,
         \56151 , \56152 , \56153 , \56154 , \56155 , \56156 , \56157 , \56158 , \56159 , \56160 ,
         \56161 , \56162 , \56163 , \56164 , \56165 , \56166 , \56167 , \56168 , \56169 , \56170 ,
         \56171 , \56172 , \56173 , \56174 , \56175 , \56176 , \56177 , \56178 , \56179 , \56180 ,
         \56181 , \56182 , \56183 , \56184 , \56185 , \56186 , \56187 , \56188 , \56189 , \56190 ,
         \56191 , \56192 , \56193 , \56194 , \56195 , \56196 , \56197 , \56198 , \56199 , \56200 ,
         \56201 , \56202 , \56203 , \56204 , \56205 , \56206 , \56207 , \56208 , \56209 , \56210 ,
         \56211 , \56212 , \56213 , \56214 , \56215 , \56216 , \56217 , \56218 , \56219 , \56220 ,
         \56221 , \56222 , \56223 , \56224 , \56225 , \56226 , \56227 , \56228 , \56229 , \56230 ,
         \56231 , \56232 , \56233 , \56234 , \56235 , \56236 , \56237 , \56238 , \56239 , \56240 ,
         \56241 , \56242 , \56243 , \56244 , \56245 , \56246 , \56247 , \56248 , \56249 , \56250 ,
         \56251 , \56252 , \56253 , \56254 , \56255 , \56256 , \56257 , \56258 , \56259 , \56260 ,
         \56261 , \56262 , \56263 , \56264 , \56265 , \56266 , \56267 , \56268 , \56269 , \56270 ,
         \56271 , \56272 , \56273 , \56274 , \56275 , \56276 , \56277 , \56278 , \56279 , \56280 ,
         \56281 , \56282 , \56283 , \56284 , \56285 , \56286 , \56287 , \56288 , \56289 , \56290 ,
         \56291 , \56292 , \56293 , \56294 , \56295 , \56296 , \56297 , \56298 , \56299 , \56300 ,
         \56301 , \56302 , \56303 , \56304 , \56305 , \56306 , \56307 , \56308 , \56309 , \56310 ,
         \56311 , \56312 , \56313 , \56314 , \56315 , \56316 , \56317 , \56318 , \56319 , \56320 ,
         \56321 , \56322 , \56323 , \56324 , \56325 , \56326 , \56327 , \56328 , \56329 , \56330 ,
         \56331 , \56332 , \56333 , \56334 , \56335 , \56336 , \56337 , \56338 , \56339 , \56340 ,
         \56341 , \56342 , \56343 , \56344 , \56345 , \56346 , \56347 , \56348 , \56349 , \56350 ,
         \56351 , \56352 , \56353 , \56354 , \56355 , \56356 , \56357 , \56358 , \56359 , \56360 ,
         \56361 , \56362 , \56363 , \56364 , \56365 , \56366 , \56367 , \56368 , \56369 , \56370 ,
         \56371 , \56372 , \56373 , \56374 , \56375 , \56376 , \56377 , \56378 , \56379 , \56380 ,
         \56381 , \56382 , \56383 , \56384 , \56385 , \56386 , \56387 , \56388 , \56389 , \56390 ,
         \56391 , \56392 , \56393 , \56394 , \56395 , \56396 , \56397 , \56398 , \56399 , \56400 ,
         \56401 , \56402 , \56403 , \56404 , \56405 , \56406 , \56407 , \56408 , \56409 , \56410 ,
         \56411 , \56412 , \56413 , \56414 , \56415 , \56416 , \56417 , \56418 , \56419 , \56420 ,
         \56421 , \56422 , \56423 , \56424 , \56425 , \56426 , \56427 , \56428 , \56429 , \56430 ,
         \56431 , \56432 , \56433 , \56434 , \56435 , \56436 , \56437 , \56438 , \56439 , \56440 ,
         \56441 , \56442 , \56443 , \56444 , \56445 , \56446 , \56447 , \56448 , \56449 , \56450 ,
         \56451 , \56452 , \56453 , \56454 , \56455 , \56456 , \56457 , \56458 , \56459 , \56460 ,
         \56461 , \56462 , \56463 , \56464 , \56465 , \56466 , \56467 , \56468 , \56469 , \56470 ,
         \56471 , \56472 , \56473 , \56474 , \56475 , \56476 , \56477 , \56478 , \56479 , \56480 ,
         \56481 , \56482 , \56483 , \56484 , \56485 , \56486 , \56487 , \56488 , \56489 , \56490 ,
         \56491 , \56492 , \56493 , \56494 , \56495 , \56496 , \56497 , \56498 , \56499 , \56500 ,
         \56501 , \56502 , \56503 , \56504 , \56505 , \56506 , \56507 , \56508 , \56509 , \56510 ,
         \56511 , \56512 , \56513 , \56514 , \56515 , \56516 , \56517 , \56518 , \56519 , \56520 ,
         \56521 , \56522 , \56523 , \56524 , \56525 , \56526 , \56527 , \56528 , \56529 , \56530 ,
         \56531 , \56532 , \56533 , \56534 , \56535 , \56536 , \56537 , \56538 , \56539 , \56540 ,
         \56541 , \56542 , \56543 , \56544 , \56545 , \56546 , \56547 , \56548 , \56549 , \56550 ,
         \56551 , \56552 , \56553 , \56554 , \56555 , \56556 , \56557 , \56558 , \56559 , \56560 ,
         \56561 , \56562 , \56563 , \56564 , \56565 , \56566 , \56567 , \56568 , \56569 , \56570 ,
         \56571 , \56572 , \56573 , \56574 , \56575 , \56576 , \56577 , \56578 , \56579 , \56580 ,
         \56581 , \56582 , \56583 , \56584 , \56585 , \56586 , \56587 , \56588 , \56589 , \56590 ,
         \56591 , \56592 , \56593 , \56594 , \56595 , \56596 , \56597 , \56598 , \56599 , \56600 ,
         \56601 , \56602 , \56603 , \56604 , \56605 , \56606 , \56607 , \56608 , \56609 , \56610 ,
         \56611 , \56612 , \56613 , \56614 , \56615 , \56616 , \56617 , \56618 , \56619 , \56620 ,
         \56621 , \56622 , \56623 , \56624 , \56625 , \56626 , \56627 , \56628 , \56629 , \56630 ,
         \56631 , \56632 , \56633 , \56634 , \56635 , \56636 , \56637 , \56638 , \56639 , \56640 ,
         \56641 , \56642 , \56643 , \56644 , \56645 , \56646 , \56647 , \56648 , \56649 , \56650 ,
         \56651 , \56652 , \56653 , \56654 , \56655 , \56656 , \56657 , \56658 , \56659 , \56660 ,
         \56661 , \56662 , \56663 , \56664 , \56665 , \56666 , \56667 , \56668 , \56669 , \56670 ,
         \56671 , \56672 , \56673 , \56674 , \56675 , \56676 , \56677 , \56678 , \56679 , \56680 ,
         \56681 , \56682 , \56683 , \56684 , \56685 , \56686 , \56687 , \56688 , \56689 , \56690 ,
         \56691 , \56692 , \56693 , \56694 , \56695 , \56696 , \56697 , \56698 , \56699 , \56700 ,
         \56701 , \56702 , \56703 , \56704 , \56705 , \56706 , \56707 , \56708 , \56709 , \56710 ,
         \56711 , \56712 , \56713 , \56714 , \56715 , \56716 , \56717 , \56718 , \56719 , \56720 ,
         \56721 , \56722 , \56723 , \56724 , \56725 , \56726 , \56727 , \56728 , \56729 , \56730 ,
         \56731 , \56732 , \56733 , \56734 , \56735 , \56736 , \56737 , \56738 , \56739 , \56740 ,
         \56741 , \56742 , \56743 , \56744 , \56745 , \56746 , \56747 , \56748 , \56749 , \56750 ,
         \56751 , \56752 , \56753 , \56754 , \56755 , \56756 , \56757 , \56758 , \56759 , \56760 ,
         \56761 , \56762 , \56763 , \56764 , \56765 , \56766 , \56767 , \56768 , \56769 , \56770 ,
         \56771 , \56772 , \56773 , \56774 , \56775 , \56776 , \56777 , \56778 , \56779 , \56780 ,
         \56781 , \56782 , \56783 , \56784 , \56785 , \56786 , \56787 , \56788 , \56789 , \56790 ,
         \56791 , \56792 , \56793 , \56794 , \56795 , \56796 , \56797 , \56798 , \56799 , \56800 ,
         \56801 , \56802 , \56803 , \56804 , \56805 , \56806 , \56807 , \56808 , \56809 , \56810 ,
         \56811 , \56812 , \56813 , \56814 , \56815 , \56816 , \56817 , \56818 , \56819 , \56820 ,
         \56821 , \56822 , \56823 , \56824 , \56825 , \56826 , \56827 , \56828 , \56829 , \56830 ,
         \56831 , \56832 , \56833 , \56834 , \56835 , \56836 , \56837 , \56838 , \56839 , \56840 ,
         \56841 , \56842 , \56843 , \56844 , \56845 , \56846 , \56847 , \56848 , \56849 , \56850 ,
         \56851 , \56852 , \56853 , \56854 , \56855 , \56856 , \56857 , \56858 , \56859 , \56860 ,
         \56861 , \56862 , \56863 , \56864 , \56865 , \56866 , \56867 , \56868 , \56869 , \56870 ,
         \56871 , \56872 , \56873 , \56874 , \56875 , \56876 , \56877 , \56878 , \56879 , \56880 ,
         \56881 , \56882 , \56883 , \56884 , \56885 , \56886 , \56887 , \56888 , \56889 , \56890 ,
         \56891 , \56892 , \56893 , \56894 , \56895 , \56896 , \56897 , \56898 , \56899 , \56900 ,
         \56901 , \56902 , \56903 , \56904 , \56905 , \56906 , \56907 , \56908 , \56909 , \56910 ,
         \56911 , \56912 , \56913 , \56914 , \56915 , \56916 , \56917 , \56918 , \56919 , \56920 ,
         \56921 , \56922 , \56923 , \56924 , \56925 , \56926 , \56927 , \56928 , \56929 , \56930 ,
         \56931 , \56932 , \56933 , \56934 , \56935 , \56936 , \56937 , \56938 , \56939 , \56940 ,
         \56941 , \56942 , \56943 , \56944 , \56945 , \56946 , \56947 , \56948 , \56949 , \56950 ,
         \56951 , \56952 , \56953 , \56954 , \56955 , \56956 , \56957 , \56958 , \56959 , \56960 ,
         \56961 , \56962 , \56963 , \56964 , \56965 , \56966 , \56967 , \56968 , \56969 , \56970 ,
         \56971 , \56972 , \56973 , \56974 , \56975 , \56976 , \56977 , \56978 , \56979 , \56980 ,
         \56981 , \56982 , \56983 , \56984 , \56985 , \56986 , \56987 , \56988 , \56989 , \56990 ,
         \56991 , \56992 , \56993 , \56994 , \56995 , \56996 , \56997 , \56998 , \56999 , \57000 ,
         \57001 , \57002 , \57003 , \57004 , \57005 , \57006 , \57007 , \57008 , \57009 , \57010 ,
         \57011 , \57012 , \57013 , \57014 , \57015 , \57016 , \57017 , \57018 , \57019 , \57020 ,
         \57021 , \57022 , \57023 , \57024 , \57025 , \57026 , \57027 , \57028 , \57029 , \57030 ,
         \57031 , \57032 , \57033 , \57034 , \57035 , \57036 , \57037 , \57038 , \57039 , \57040 ,
         \57041 , \57042 , \57043 , \57044 , \57045 , \57046 , \57047 , \57048 , \57049 , \57050 ,
         \57051 , \57052 , \57053 , \57054 , \57055 , \57056 , \57057 , \57058 , \57059 , \57060 ,
         \57061 , \57062 , \57063 , \57064 , \57065 , \57066 , \57067 , \57068 , \57069 , \57070 ,
         \57071 , \57072 , \57073 , \57074 , \57075 , \57076 , \57077 , \57078 , \57079 , \57080 ,
         \57081 , \57082 , \57083 , \57084 , \57085 , \57086 , \57087 , \57088 , \57089 , \57090 ,
         \57091 , \57092 , \57093 , \57094 , \57095 , \57096 , \57097 , \57098 , \57099 , \57100 ,
         \57101 , \57102 , \57103 , \57104 , \57105 , \57106 , \57107 , \57108 , \57109 , \57110 ,
         \57111 , \57112 , \57113 , \57114 , \57115 , \57116 , \57117 , \57118 , \57119 , \57120 ,
         \57121 , \57122 , \57123 , \57124 , \57125 , \57126 , \57127 , \57128 , \57129 , \57130 ,
         \57131 , \57132 , \57133 , \57134 , \57135 , \57136 , \57137 , \57138 , \57139 , \57140 ,
         \57141 , \57142 , \57143 , \57144 , \57145 , \57146 , \57147 , \57148 , \57149 , \57150 ,
         \57151 , \57152 , \57153 , \57154 , \57155 , \57156 , \57157 , \57158 , \57159 , \57160 ,
         \57161 , \57162 , \57163 , \57164 , \57165 , \57166 , \57167 , \57168 , \57169 , \57170 ,
         \57171 , \57172 , \57173 , \57174 , \57175 , \57176 , \57177 , \57178 , \57179 , \57180 ,
         \57181 , \57182 , \57183 , \57184 , \57185 , \57186 , \57187 , \57188 , \57189 , \57190 ,
         \57191 , \57192 , \57193 , \57194 , \57195 , \57196 , \57197 , \57198 , \57199 , \57200 ,
         \57201 , \57202 , \57203 , \57204 , \57205 , \57206 , \57207 , \57208 , \57209 , \57210 ,
         \57211 , \57212 , \57213 , \57214 , \57215 , \57216 , \57217 , \57218 , \57219 , \57220 ,
         \57221 , \57222 , \57223 , \57224 , \57225 , \57226 , \57227 , \57228 , \57229 , \57230 ,
         \57231 , \57232 , \57233 , \57234 , \57235 , \57236 , \57237 , \57238 , \57239 , \57240 ,
         \57241 , \57242 , \57243 , \57244 , \57245 , \57246 , \57247 , \57248 , \57249 , \57250 ,
         \57251 , \57252 , \57253 , \57254 , \57255 , \57256 , \57257 , \57258 , \57259 , \57260 ,
         \57261 , \57262 , \57263 , \57264 , \57265 , \57266 , \57267 , \57268 , \57269 , \57270 ,
         \57271 , \57272 , \57273 , \57274 , \57275 , \57276 , \57277 , \57278 , \57279 , \57280 ,
         \57281 , \57282 , \57283 , \57284 , \57285 , \57286 , \57287 , \57288 , \57289 , \57290 ,
         \57291 , \57292 , \57293 , \57294 , \57295 , \57296 , \57297 , \57298 , \57299 , \57300 ,
         \57301 , \57302 , \57303 , \57304 , \57305 , \57306 , \57307 , \57308 , \57309 , \57310 ,
         \57311 , \57312 , \57313 , \57314 , \57315 , \57316 , \57317 , \57318 , \57319 , \57320 ,
         \57321 , \57322 , \57323 , \57324 , \57325 , \57326 , \57327 , \57328 , \57329 , \57330 ,
         \57331 , \57332 , \57333 , \57334 , \57335 , \57336 , \57337 , \57338 , \57339 , \57340 ,
         \57341 , \57342 , \57343 , \57344 , \57345 , \57346 , \57347 , \57348 , \57349 , \57350 ,
         \57351 , \57352 , \57353 , \57354 , \57355 , \57356 , \57357 , \57358 , \57359 , \57360 ,
         \57361 , \57362 , \57363 , \57364 , \57365 , \57366 , \57367 , \57368 , \57369 , \57370 ,
         \57371 , \57372 , \57373 , \57374 , \57375 , \57376 , \57377 , \57378 , \57379 , \57380 ,
         \57381 , \57382 , \57383 , \57384 , \57385 , \57386 , \57387 , \57388 , \57389 , \57390 ,
         \57391 , \57392 , \57393 , \57394 , \57395 , \57396 , \57397 , \57398 , \57399 , \57400 ,
         \57401 , \57402 , \57403 , \57404 , \57405 , \57406 , \57407 , \57408 , \57409 , \57410 ,
         \57411 , \57412 , \57413 , \57414 , \57415 , \57416 , \57417 , \57418 , \57419 , \57420 ,
         \57421 , \57422 , \57423 , \57424 , \57425 , \57426 , \57427 , \57428 , \57429 , \57430 ,
         \57431 , \57432 , \57433 , \57434 , \57435 , \57436 , \57437 , \57438 , \57439 , \57440 ,
         \57441 , \57442 , \57443 , \57444 , \57445 , \57446 , \57447 , \57448 , \57449 , \57450 ,
         \57451 , \57452 , \57453 , \57454 , \57455 , \57456 , \57457 , \57458 , \57459 , \57460 ,
         \57461 , \57462 , \57463 , \57464 , \57465 , \57466 , \57467 , \57468 , \57469 , \57470 ,
         \57471 , \57472 , \57473 , \57474 , \57475 , \57476 , \57477 , \57478 , \57479 , \57480 ,
         \57481 , \57482 , \57483 , \57484 , \57485 , \57486 , \57487 , \57488 , \57489 , \57490 ,
         \57491 , \57492 , \57493 , \57494 , \57495 , \57496 , \57497 , \57498 , \57499 , \57500 ,
         \57501 , \57502 , \57503 , \57504 , \57505 , \57506 , \57507 , \57508 , \57509 , \57510 ,
         \57511 , \57512 , \57513 , \57514 , \57515 , \57516 , \57517 , \57518 , \57519 , \57520 ,
         \57521 , \57522 , \57523 , \57524 , \57525 , \57526 , \57527 , \57528 , \57529 , \57530 ,
         \57531 , \57532 , \57533 , \57534 , \57535 , \57536 , \57537 , \57538 , \57539 , \57540 ,
         \57541 , \57542 , \57543 , \57544 , \57545 , \57546 , \57547 , \57548 , \57549 , \57550 ,
         \57551 , \57552 , \57553 , \57554 , \57555 , \57556 , \57557 , \57558 , \57559 , \57560 ,
         \57561 , \57562 , \57563 , \57564 , \57565 , \57566 , \57567 , \57568 , \57569 , \57570 ,
         \57571 , \57572 , \57573 , \57574 , \57575 , \57576 , \57577 , \57578 , \57579 , \57580 ,
         \57581 , \57582 , \57583 , \57584 , \57585 , \57586 , \57587 , \57588 , \57589 , \57590 ,
         \57591 , \57592 , \57593 , \57594 , \57595 , \57596 , \57597 , \57598 , \57599 , \57600 ,
         \57601 , \57602 , \57603 , \57604 , \57605 , \57606 , \57607 , \57608 , \57609 , \57610 ,
         \57611 , \57612 , \57613 , \57614 , \57615 , \57616 , \57617 , \57618 , \57619 , \57620 ,
         \57621 , \57622 , \57623 , \57624 , \57625 , \57626 , \57627 , \57628 , \57629 , \57630 ,
         \57631 , \57632 , \57633 , \57634 , \57635 , \57636 , \57637 , \57638 , \57639 , \57640 ,
         \57641 , \57642 , \57643 , \57644 , \57645 , \57646 , \57647 , \57648 , \57649 , \57650 ,
         \57651 , \57652 , \57653 , \57654 , \57655 , \57656 , \57657 , \57658 , \57659 , \57660 ,
         \57661 , \57662 , \57663 , \57664 , \57665 , \57666 , \57667 , \57668 , \57669 , \57670 ,
         \57671 , \57672 , \57673 , \57674 , \57675 , \57676 , \57677 , \57678 , \57679 , \57680 ,
         \57681 , \57682 , \57683 , \57684 , \57685 , \57686 , \57687 , \57688 , \57689 , \57690 ,
         \57691 , \57692 , \57693 , \57694 , \57695 , \57696 , \57697 , \57698 , \57699 , \57700 ,
         \57701 , \57702 , \57703 , \57704 , \57705 , \57706 , \57707 , \57708 , \57709 , \57710 ,
         \57711 , \57712 , \57713 , \57714 , \57715 , \57716 , \57717 , \57718 , \57719 , \57720 ,
         \57721 , \57722 , \57723 , \57724 , \57725 , \57726 , \57727 , \57728 , \57729 , \57730 ,
         \57731 , \57732 , \57733 , \57734 , \57735 , \57736 , \57737 , \57738 , \57739 , \57740 ,
         \57741 , \57742 , \57743 , \57744 , \57745 , \57746 , \57747 , \57748 , \57749 , \57750 ,
         \57751 , \57752 , \57753 , \57754 , \57755 , \57756 , \57757 , \57758 , \57759 , \57760 ,
         \57761 , \57762 , \57763 , \57764 , \57765 , \57766 , \57767 , \57768 , \57769 , \57770 ,
         \57771 , \57772 , \57773 , \57774 , \57775 , \57776 , \57777 , \57778 , \57779 , \57780 ,
         \57781 , \57782 , \57783 , \57784 , \57785 , \57786 , \57787 , \57788 , \57789 , \57790 ,
         \57791 , \57792 , \57793 , \57794 , \57795 , \57796 , \57797 , \57798 , \57799 , \57800 ,
         \57801 , \57802 , \57803 , \57804 , \57805 , \57806 , \57807 , \57808 , \57809 , \57810 ,
         \57811 , \57812 , \57813 , \57814 , \57815 , \57816 , \57817 , \57818 , \57819 , \57820 ,
         \57821 , \57822 , \57823 , \57824 , \57825 , \57826 , \57827 , \57828 , \57829 , \57830 ,
         \57831 , \57832 , \57833 , \57834 , \57835 , \57836 , \57837 , \57838 , \57839 , \57840 ,
         \57841 , \57842 , \57843 , \57844 , \57845 , \57846 , \57847 , \57848 , \57849 , \57850 ,
         \57851 , \57852 , \57853 , \57854 , \57855 , \57856 , \57857 , \57858 , \57859 , \57860 ,
         \57861 , \57862 , \57863 , \57864 , \57865 , \57866 , \57867 , \57868 , \57869 , \57870 ,
         \57871 , \57872 , \57873 , \57874 , \57875 , \57876 , \57877 , \57878 , \57879 , \57880 ,
         \57881 , \57882 , \57883 , \57884 , \57885 , \57886 , \57887 , \57888 , \57889 , \57890 ,
         \57891 , \57892 , \57893 , \57894 , \57895 , \57896 , \57897 , \57898 , \57899 , \57900 ,
         \57901 , \57902 , \57903 , \57904 , \57905 , \57906 , \57907 , \57908 , \57909 , \57910 ,
         \57911 , \57912 , \57913 , \57914 , \57915 , \57916 , \57917 , \57918 , \57919 , \57920 ,
         \57921 , \57922 , \57923 , \57924 , \57925 , \57926 , \57927 , \57928 , \57929 , \57930 ,
         \57931 , \57932 , \57933 , \57934 , \57935 , \57936 , \57937 , \57938 , \57939 , \57940 ,
         \57941 , \57942 , \57943 , \57944 , \57945 , \57946 , \57947 , \57948 , \57949 , \57950 ,
         \57951 , \57952 , \57953 , \57954 , \57955 , \57956 , \57957 , \57958 , \57959 , \57960 ,
         \57961 , \57962 , \57963 , \57964 , \57965 , \57966 , \57967 , \57968 , \57969 , \57970 ,
         \57971 , \57972 , \57973 , \57974 , \57975 , \57976 , \57977 , \57978 , \57979 , \57980 ,
         \57981 , \57982 , \57983 , \57984 , \57985 , \57986 , \57987 , \57988 , \57989 , \57990 ,
         \57991 , \57992 , \57993 , \57994 , \57995 , \57996 , \57997 , \57998 , \57999 , \58000 ,
         \58001 , \58002 , \58003 , \58004 , \58005 , \58006 , \58007 , \58008 , \58009 , \58010 ,
         \58011 , \58012 , \58013 , \58014 , \58015 , \58016 , \58017 , \58018 , \58019 , \58020 ,
         \58021 , \58022 , \58023 , \58024 , \58025 , \58026 , \58027 , \58028 , \58029 , \58030 ,
         \58031 , \58032 , \58033 , \58034 , \58035 , \58036 , \58037 , \58038 , \58039 , \58040 ,
         \58041 , \58042 , \58043 , \58044 , \58045 , \58046 , \58047 , \58048 , \58049 , \58050 ,
         \58051 , \58052 , \58053 , \58054 , \58055 , \58056 , \58057 , \58058 , \58059 , \58060 ,
         \58061 , \58062 , \58063 , \58064 , \58065 , \58066 , \58067 , \58068 , \58069 , \58070 ,
         \58071 , \58072 , \58073 , \58074 , \58075 , \58076 , \58077 , \58078 , \58079 , \58080 ,
         \58081 , \58082 , \58083 , \58084 , \58085 , \58086 , \58087 , \58088 , \58089 , \58090 ,
         \58091 , \58092 , \58093 , \58094 , \58095 , \58096 , \58097 , \58098 , \58099 , \58100 ,
         \58101 , \58102 , \58103 , \58104 , \58105 , \58106 , \58107 , \58108 , \58109 , \58110 ,
         \58111 , \58112 , \58113 , \58114 , \58115 , \58116 , \58117 , \58118 , \58119 , \58120 ,
         \58121 , \58122 , \58123 , \58124 , \58125 , \58126 , \58127 , \58128 , \58129 , \58130 ,
         \58131 , \58132 , \58133 , \58134 , \58135 , \58136 , \58137 , \58138 , \58139 , \58140 ,
         \58141 , \58142 , \58143 , \58144 , \58145 , \58146 , \58147 , \58148 , \58149 , \58150 ,
         \58151 , \58152 , \58153 , \58154 , \58155 , \58156 , \58157 , \58158 , \58159 , \58160 ,
         \58161 , \58162 , \58163 , \58164 , \58165 , \58166 , \58167 , \58168 , \58169 , \58170 ,
         \58171 , \58172 , \58173 , \58174 , \58175 , \58176 , \58177 , \58178 , \58179 , \58180 ,
         \58181 , \58182 , \58183 , \58184 , \58185 , \58186 , \58187 , \58188 , \58189 , \58190 ,
         \58191 , \58192 , \58193 , \58194 , \58195 , \58196 , \58197 , \58198 , \58199 , \58200 ,
         \58201 , \58202 , \58203 , \58204 , \58205 , \58206 , \58207 , \58208 , \58209 , \58210 ,
         \58211 , \58212 , \58213 , \58214 , \58215 , \58216 , \58217 , \58218 , \58219 , \58220 ,
         \58221 , \58222 , \58223 , \58224 , \58225 , \58226 , \58227 , \58228 , \58229 , \58230 ,
         \58231 , \58232 , \58233 , \58234 , \58235 , \58236 , \58237 , \58238 , \58239 , \58240 ,
         \58241 , \58242 , \58243 , \58244 , \58245 , \58246 , \58247 , \58248 , \58249 , \58250 ,
         \58251 , \58252 , \58253 , \58254 , \58255 , \58256 , \58257 , \58258 , \58259 , \58260 ,
         \58261 , \58262 , \58263 , \58264 , \58265 , \58266 , \58267 , \58268 , \58269 , \58270 ,
         \58271 , \58272 , \58273 , \58274 , \58275 , \58276 , \58277 , \58278 , \58279 , \58280 ,
         \58281 , \58282 , \58283 , \58284 , \58285 , \58286 , \58287 , \58288 , \58289 , \58290 ,
         \58291 , \58292 , \58293 , \58294 , \58295 , \58296 , \58297 , \58298 , \58299 , \58300 ,
         \58301 , \58302 , \58303 , \58304 , \58305 , \58306 , \58307 , \58308 , \58309 , \58310 ,
         \58311 , \58312 , \58313 , \58314 , \58315 , \58316 , \58317 , \58318 , \58319 , \58320 ,
         \58321 , \58322 , \58323 , \58324 , \58325 , \58326 , \58327 , \58328 , \58329 , \58330 ,
         \58331 , \58332 , \58333 , \58334 , \58335 , \58336 , \58337 , \58338 , \58339 , \58340 ,
         \58341 , \58342 , \58343 , \58344 , \58345 , \58346 , \58347 , \58348 , \58349 , \58350 ,
         \58351 , \58352 , \58353 , \58354 , \58355 , \58356 , \58357 , \58358 , \58359 , \58360 ,
         \58361 , \58362 , \58363 , \58364 , \58365 , \58366 , \58367 , \58368 , \58369 , \58370 ,
         \58371 , \58372 , \58373 , \58374 , \58375 , \58376 , \58377 , \58378 , \58379 , \58380 ,
         \58381 , \58382 , \58383 , \58384 , \58385 , \58386 , \58387 , \58388 , \58389 , \58390 ,
         \58391 , \58392 , \58393 , \58394 , \58395 , \58396 , \58397 , \58398 , \58399 , \58400 ,
         \58401 , \58402 , \58403 , \58404 , \58405 , \58406 , \58407 , \58408 , \58409 , \58410 ,
         \58411 , \58412 , \58413 , \58414 , \58415 , \58416 , \58417 , \58418 , \58419 , \58420 ,
         \58421 , \58422 , \58423 , \58424 , \58425 , \58426 , \58427 , \58428 , \58429 , \58430 ,
         \58431 , \58432 , \58433 , \58434 , \58435 , \58436 , \58437 , \58438 , \58439 , \58440 ,
         \58441 , \58442 , \58443 , \58444 , \58445 , \58446 , \58447 , \58448 , \58449 , \58450 ,
         \58451 , \58452 , \58453 , \58454 , \58455 , \58456 , \58457 , \58458 , \58459 , \58460 ,
         \58461 , \58462 , \58463 , \58464 , \58465 , \58466 , \58467 , \58468 , \58469 , \58470 ,
         \58471 , \58472 , \58473 , \58474 , \58475 , \58476 , \58477 , \58478 , \58479 , \58480 ,
         \58481 , \58482 , \58483 , \58484 , \58485 , \58486 , \58487 , \58488 , \58489 , \58490 ,
         \58491 , \58492 , \58493 , \58494 , \58495 , \58496 , \58497 , \58498 , \58499 , \58500 ,
         \58501 , \58502 , \58503 , \58504 , \58505 , \58506 , \58507 , \58508 , \58509 , \58510 ,
         \58511 , \58512 , \58513 , \58514 , \58515 , \58516 , \58517 , \58518 , \58519 , \58520 ,
         \58521 , \58522 , \58523 , \58524 , \58525 , \58526 , \58527 , \58528 , \58529 , \58530 ,
         \58531 , \58532 , \58533 , \58534 , \58535 , \58536 , \58537 , \58538 , \58539 , \58540 ,
         \58541 , \58542 , \58543 , \58544 , \58545 , \58546 , \58547 , \58548 , \58549 , \58550 ,
         \58551 , \58552 , \58553 , \58554 , \58555 , \58556 , \58557 , \58558 , \58559 , \58560 ,
         \58561 , \58562 , \58563 , \58564 , \58565 , \58566 , \58567 , \58568 , \58569 , \58570 ,
         \58571 , \58572 , \58573 , \58574 , \58575 , \58576 , \58577 , \58578 , \58579 , \58580 ,
         \58581 , \58582 , \58583 , \58584 , \58585 , \58586 , \58587 , \58588 , \58589 , \58590 ,
         \58591 , \58592 , \58593 , \58594 , \58595 , \58596 , \58597 , \58598 , \58599 , \58600 ,
         \58601 , \58602 , \58603 , \58604 , \58605 , \58606 , \58607 , \58608 , \58609 , \58610 ,
         \58611 , \58612 , \58613 , \58614 , \58615 , \58616 , \58617 , \58618 , \58619 , \58620 ,
         \58621 , \58622 , \58623 , \58624 , \58625 , \58626 , \58627 , \58628 , \58629 , \58630 ,
         \58631 , \58632 , \58633 , \58634 , \58635 , \58636 , \58637 , \58638 , \58639 , \58640 ,
         \58641 , \58642 , \58643 , \58644 , \58645 , \58646 , \58647 , \58648 , \58649 , \58650 ,
         \58651 , \58652 , \58653 , \58654 , \58655 , \58656 , \58657 , \58658 , \58659 , \58660 ,
         \58661 , \58662 , \58663 , \58664 , \58665 , \58666 , \58667 , \58668 , \58669 , \58670 ,
         \58671 , \58672 , \58673 , \58674 , \58675 , \58676 , \58677 , \58678 , \58679 , \58680 ,
         \58681 , \58682 , \58683 , \58684 , \58685 , \58686 , \58687 , \58688 , \58689 , \58690 ,
         \58691 , \58692 , \58693 , \58694 , \58695 , \58696 , \58697 , \58698 , \58699 , \58700 ,
         \58701 , \58702 , \58703 , \58704 , \58705 , \58706 , \58707 , \58708 , \58709 , \58710 ,
         \58711 , \58712 , \58713 , \58714 , \58715 , \58716 , \58717 , \58718 , \58719 , \58720 ,
         \58721 , \58722 , \58723 , \58724 , \58725 , \58726 , \58727 , \58728 , \58729 , \58730 ,
         \58731 , \58732 , \58733 , \58734 , \58735 , \58736 , \58737 , \58738 , \58739 , \58740 ,
         \58741 , \58742 , \58743 , \58744 , \58745 , \58746 , \58747 , \58748 , \58749 , \58750 ,
         \58751 , \58752 , \58753 , \58754 , \58755 , \58756 , \58757 , \58758 , \58759 , \58760 ,
         \58761 , \58762 , \58763 , \58764 , \58765 , \58766 , \58767 , \58768 , \58769 , \58770 ,
         \58771 , \58772 , \58773 , \58774 , \58775 , \58776 , \58777 , \58778 , \58779 , \58780 ,
         \58781 , \58782 , \58783 , \58784 , \58785 , \58786 , \58787 , \58788 , \58789 , \58790 ,
         \58791 , \58792 , \58793 , \58794 , \58795 , \58796 , \58797 , \58798 , \58799 , \58800 ,
         \58801 , \58802 , \58803 , \58804 , \58805 , \58806 , \58807 , \58808 , \58809 , \58810 ,
         \58811 , \58812 , \58813 , \58814 , \58815 , \58816 , \58817 , \58818 , \58819 , \58820 ,
         \58821 , \58822 , \58823 , \58824 , \58825 , \58826 , \58827 , \58828 , \58829 , \58830 ,
         \58831 , \58832 , \58833 , \58834 , \58835 , \58836 , \58837 , \58838 , \58839 , \58840 ,
         \58841 , \58842 , \58843 , \58844 , \58845 , \58846 , \58847 , \58848 , \58849 , \58850 ,
         \58851 , \58852 , \58853 , \58854 , \58855 , \58856 , \58857 , \58858 , \58859 , \58860 ,
         \58861 , \58862 , \58863 , \58864 , \58865 , \58866 , \58867 , \58868 , \58869 , \58870 ,
         \58871 , \58872 , \58873 , \58874 , \58875 , \58876 , \58877 , \58878 , \58879 , \58880 ,
         \58881 , \58882 , \58883 , \58884 , \58885 , \58886 , \58887 , \58888 , \58889 , \58890 ,
         \58891 , \58892 , \58893 , \58894 , \58895 , \58896 , \58897 , \58898 , \58899 , \58900 ,
         \58901 , \58902 , \58903 , \58904 , \58905 , \58906 , \58907 , \58908 , \58909 , \58910 ,
         \58911 , \58912 , \58913 , \58914 , \58915 , \58916 , \58917 , \58918 , \58919 , \58920 ,
         \58921 , \58922 , \58923 , \58924 , \58925 , \58926 , \58927 , \58928 , \58929 , \58930 ,
         \58931 , \58932 , \58933 , \58934 , \58935 , \58936 , \58937 , \58938 , \58939 , \58940 ,
         \58941 , \58942 , \58943 , \58944 , \58945 , \58946 , \58947 , \58948 , \58949 , \58950 ,
         \58951 , \58952 , \58953 , \58954 , \58955 , \58956 , \58957 , \58958 , \58959 , \58960 ,
         \58961 , \58962 , \58963 , \58964 , \58965 , \58966 , \58967 , \58968 , \58969 , \58970 ,
         \58971 , \58972 , \58973 , \58974 , \58975 , \58976 , \58977 , \58978 , \58979 , \58980 ,
         \58981 , \58982 , \58983 , \58984 , \58985 , \58986 , \58987 , \58988 , \58989 , \58990 ,
         \58991 , \58992 , \58993 , \58994 , \58995 , \58996 , \58997 , \58998 , \58999 , \59000 ,
         \59001 , \59002 , \59003 , \59004 , \59005 , \59006 , \59007 , \59008 , \59009 , \59010 ,
         \59011 , \59012 , \59013 , \59014 , \59015 , \59016 , \59017 , \59018 , \59019 , \59020 ,
         \59021 , \59022 , \59023 , \59024 , \59025 , \59026 , \59027 , \59028 , \59029 , \59030 ,
         \59031 , \59032 , \59033 , \59034 , \59035 , \59036 , \59037 , \59038 , \59039 , \59040 ,
         \59041 , \59042 , \59043 , \59044 , \59045 , \59046 , \59047 , \59048 , \59049 , \59050 ,
         \59051 , \59052 , \59053 , \59054 , \59055 , \59056 , \59057 , \59058 , \59059 , \59060 ,
         \59061 , \59062 , \59063 , \59064 , \59065 , \59066 , \59067 , \59068 , \59069 , \59070 ,
         \59071 , \59072 , \59073 , \59074 , \59075 , \59076 , \59077 , \59078 , \59079 , \59080 ,
         \59081 , \59082 , \59083 , \59084 , \59085 , \59086 , \59087 , \59088 , \59089 , \59090 ,
         \59091 , \59092 , \59093 , \59094 , \59095 , \59096 , \59097 , \59098 , \59099 , \59100 ,
         \59101 , \59102 , \59103 , \59104 , \59105 , \59106 , \59107 , \59108 , \59109 , \59110 ,
         \59111 , \59112 , \59113 , \59114 , \59115 , \59116 , \59117 , \59118 , \59119 , \59120 ,
         \59121 , \59122 , \59123 , \59124 , \59125 , \59126 , \59127 , \59128 , \59129 , \59130 ,
         \59131 , \59132 , \59133 , \59134 , \59135 , \59136 , \59137 , \59138 , \59139 , \59140 ,
         \59141 , \59142 , \59143 , \59144 , \59145 , \59146 , \59147 , \59148 , \59149 , \59150 ,
         \59151 , \59152 , \59153 , \59154 , \59155 , \59156 , \59157 , \59158 , \59159 , \59160 ,
         \59161 , \59162 , \59163 , \59164 , \59165 , \59166 , \59167 , \59168 , \59169 , \59170 ,
         \59171 , \59172 , \59173 , \59174 , \59175 , \59176 , \59177 , \59178 , \59179 , \59180 ,
         \59181 , \59182 , \59183 , \59184 , \59185 , \59186 , \59187 , \59188 , \59189 , \59190 ,
         \59191 , \59192 , \59193 , \59194 , \59195 , \59196 , \59197 , \59198 , \59199 , \59200 ,
         \59201 , \59202 , \59203 , \59204 , \59205 , \59206 , \59207 , \59208 , \59209 , \59210 ,
         \59211 , \59212 , \59213 , \59214 , \59215 , \59216 , \59217 , \59218 , \59219 , \59220 ,
         \59221 , \59222 , \59223 , \59224 , \59225 , \59226 , \59227 , \59228 , \59229 , \59230 ,
         \59231 , \59232 , \59233 , \59234 , \59235 , \59236 , \59237 , \59238 , \59239 , \59240 ,
         \59241 , \59242 , \59243 , \59244 , \59245 , \59246 , \59247 , \59248 , \59249 , \59250 ,
         \59251 , \59252 , \59253 , \59254 , \59255 , \59256 , \59257 , \59258 , \59259 , \59260 ,
         \59261 , \59262 , \59263 , \59264 , \59265 , \59266 , \59267 , \59268 , \59269 , \59270 ,
         \59271 , \59272 , \59273 , \59274 , \59275 , \59276 , \59277 , \59278 , \59279 , \59280 ,
         \59281 , \59282 , \59283 , \59284 , \59285 , \59286 , \59287 , \59288 , \59289 , \59290 ,
         \59291 , \59292 , \59293 , \59294 , \59295 , \59296 , \59297 , \59298 , \59299 , \59300 ,
         \59301 , \59302 , \59303 , \59304 , \59305 , \59306 , \59307 , \59308 , \59309 , \59310 ,
         \59311 , \59312 , \59313 , \59314 , \59315 , \59316 , \59317 , \59318 , \59319 , \59320 ,
         \59321 , \59322 , \59323 , \59324 , \59325 , \59326 , \59327 , \59328 , \59329 , \59330 ,
         \59331 , \59332 , \59333 , \59334 , \59335 , \59336 , \59337 , \59338 , \59339 , \59340 ,
         \59341 , \59342 , \59343 , \59344 , \59345 , \59346 , \59347 , \59348 , \59349 , \59350 ,
         \59351 , \59352 , \59353 , \59354 , \59355 , \59356 , \59357 , \59358 , \59359 , \59360 ,
         \59361 , \59362 , \59363 , \59364 , \59365 , \59366 , \59367 , \59368 , \59369 , \59370 ,
         \59371 , \59372 , \59373 , \59374 , \59375 , \59376 , \59377 , \59378 , \59379 , \59380 ,
         \59381 , \59382 , \59383 , \59384 , \59385 , \59386 , \59387 , \59388 , \59389 , \59390 ,
         \59391 , \59392 , \59393 , \59394 , \59395 , \59396 , \59397 , \59398 , \59399 , \59400 ,
         \59401 , \59402 , \59403 , \59404 , \59405 , \59406 , \59407 , \59408 , \59409 , \59410 ,
         \59411 , \59412 , \59413 , \59414 , \59415 , \59416 , \59417 , \59418 , \59419 , \59420 ,
         \59421 , \59422 , \59423 , \59424 , \59425 , \59426 , \59427 , \59428 , \59429 , \59430 ,
         \59431 , \59432 , \59433 , \59434 , \59435 , \59436 , \59437 , \59438 , \59439 , \59440 ,
         \59441 , \59442 , \59443 , \59444 , \59445 , \59446 , \59447 , \59448 , \59449 , \59450 ,
         \59451 , \59452 , \59453 , \59454 , \59455 , \59456 , \59457 , \59458 , \59459 , \59460 ,
         \59461 , \59462 , \59463 , \59464 , \59465 , \59466 , \59467 , \59468 , \59469 , \59470 ,
         \59471 , \59472 , \59473 , \59474 , \59475 , \59476 , \59477 , \59478 , \59479 , \59480 ,
         \59481 , \59482 , \59483 , \59484 , \59485 , \59486 , \59487 , \59488 , \59489 , \59490 ,
         \59491 , \59492 , \59493 , \59494 , \59495 , \59496 , \59497 , \59498 , \59499 , \59500 ,
         \59501 , \59502 , \59503 , \59504 , \59505 , \59506 , \59507 , \59508 , \59509 , \59510 ,
         \59511 , \59512 , \59513 , \59514 , \59515 , \59516 , \59517 , \59518 , \59519 , \59520 ,
         \59521 , \59522 , \59523 , \59524 , \59525 , \59526 , \59527 , \59528 , \59529 , \59530 ,
         \59531 , \59532 , \59533 , \59534 , \59535 , \59536 , \59537 , \59538 , \59539 , \59540 ,
         \59541 , \59542 , \59543 , \59544 , \59545 , \59546 , \59547 , \59548 , \59549 , \59550 ,
         \59551 , \59552 , \59553 , \59554 , \59555 , \59556 , \59557 , \59558 , \59559 , \59560 ,
         \59561 , \59562 , \59563 , \59564 , \59565 , \59566 , \59567 , \59568 , \59569 , \59570 ,
         \59571 , \59572 , \59573 , \59574 , \59575 , \59576 , \59577 , \59578 , \59579 , \59580 ,
         \59581 , \59582 , \59583 , \59584 , \59585 , \59586 , \59587 , \59588 , \59589 , \59590 ,
         \59591 , \59592 , \59593 , \59594 , \59595 , \59596 , \59597 , \59598 , \59599 , \59600 ,
         \59601 , \59602 , \59603 , \59604 , \59605 , \59606 , \59607 , \59608 , \59609 , \59610 ,
         \59611 , \59612 , \59613 , \59614 , \59615 , \59616 , \59617 , \59618 , \59619 , \59620 ,
         \59621 , \59622 , \59623 , \59624 , \59625 , \59626 , \59627 , \59628 , \59629 , \59630 ,
         \59631 , \59632 , \59633 , \59634 , \59635 , \59636 , \59637 , \59638 , \59639 , \59640 ,
         \59641 , \59642 , \59643 , \59644 , \59645 , \59646 , \59647 , \59648 , \59649 , \59650 ,
         \59651 , \59652 , \59653 , \59654 , \59655 , \59656 , \59657 , \59658 , \59659 , \59660 ,
         \59661 , \59662 , \59663 , \59664 , \59665 , \59666 , \59667 , \59668 , \59669 , \59670 ,
         \59671 , \59672 , \59673 , \59674 , \59675 , \59676 , \59677 , \59678 , \59679 , \59680 ,
         \59681 , \59682 , \59683 , \59684 , \59685 , \59686 , \59687 , \59688 , \59689 , \59690 ,
         \59691 , \59692 , \59693 , \59694 , \59695 , \59696 , \59697 , \59698 , \59699 , \59700 ,
         \59701 , \59702 , \59703 , \59704 , \59705 , \59706 , \59707 , \59708 , \59709 , \59710 ,
         \59711 , \59712 , \59713 , \59714 , \59715 , \59716 , \59717 , \59718 , \59719 , \59720 ,
         \59721 , \59722 , \59723 , \59724 , \59725 , \59726 , \59727 , \59728 , \59729 , \59730 ,
         \59731 , \59732 , \59733 , \59734 , \59735 , \59736 , \59737 , \59738 , \59739 , \59740 ,
         \59741 , \59742 , \59743 , \59744 , \59745 , \59746 , \59747 , \59748 , \59749 , \59750 ,
         \59751 , \59752 , \59753 , \59754 , \59755 , \59756 , \59757 , \59758 , \59759 , \59760 ,
         \59761 , \59762 , \59763 , \59764 , \59765 , \59766 , \59767 , \59768 , \59769 , \59770 ,
         \59771 , \59772 , \59773 , \59774 , \59775 , \59776 , \59777 , \59778 , \59779 , \59780 ,
         \59781 , \59782 , \59783 , \59784 , \59785 , \59786 , \59787 , \59788 , \59789 , \59790 ,
         \59791 , \59792 , \59793 , \59794 , \59795 , \59796 , \59797 , \59798 , \59799 , \59800 ,
         \59801 , \59802 , \59803 , \59804 , \59805 , \59806 , \59807 , \59808 , \59809 , \59810 ,
         \59811 , \59812 , \59813 , \59814 , \59815 , \59816 , \59817 , \59818 , \59819 , \59820 ,
         \59821 , \59822 , \59823 , \59824 , \59825 , \59826 , \59827 , \59828 , \59829 , \59830 ,
         \59831 , \59832 , \59833 , \59834 , \59835 , \59836 , \59837 , \59838 , \59839 , \59840 ,
         \59841 , \59842 , \59843 , \59844 , \59845 , \59846 , \59847 , \59848 , \59849 , \59850 ,
         \59851 , \59852 , \59853 , \59854 , \59855 , \59856 , \59857 , \59858 , \59859 , \59860 ,
         \59861 , \59862 , \59863 , \59864 , \59865 , \59866 , \59867 , \59868 , \59869 , \59870 ,
         \59871 , \59872 , \59873 , \59874 , \59875 , \59876 , \59877 , \59878 , \59879 , \59880 ,
         \59881 , \59882 , \59883 , \59884 , \59885 , \59886 , \59887 , \59888 , \59889 , \59890 ,
         \59891 , \59892 , \59893 , \59894 , \59895 , \59896 , \59897 , \59898 , \59899 , \59900 ,
         \59901 , \59902 , \59903 , \59904 , \59905 , \59906 , \59907 , \59908 , \59909 , \59910 ,
         \59911 , \59912 , \59913 , \59914 , \59915 , \59916 , \59917 , \59918 , \59919 , \59920 ,
         \59921 , \59922 , \59923 , \59924 , \59925 , \59926 , \59927 , \59928 , \59929 , \59930 ,
         \59931 , \59932 , \59933 , \59934 , \59935 , \59936 , \59937 , \59938 , \59939 , \59940 ,
         \59941 , \59942 , \59943 , \59944 , \59945 , \59946 , \59947 , \59948 , \59949 , \59950 ,
         \59951 , \59952 , \59953 , \59954 , \59955 , \59956 , \59957 , \59958 , \59959 , \59960 ,
         \59961 , \59962 , \59963 , \59964 , \59965 , \59966 , \59967 , \59968 , \59969 , \59970 ,
         \59971 , \59972 , \59973 , \59974 , \59975 , \59976 , \59977 , \59978 , \59979 , \59980 ,
         \59981 , \59982 , \59983 , \59984 , \59985 , \59986 , \59987 , \59988 , \59989 , \59990 ,
         \59991 , \59992 , \59993 , \59994 , \59995 , \59996 , \59997 , \59998 , \59999 , \60000 ,
         \60001 , \60002 , \60003 , \60004 , \60005 , \60006 , \60007 , \60008 , \60009 , \60010 ,
         \60011 , \60012 , \60013 , \60014 , \60015 , \60016 , \60017 , \60018 , \60019 , \60020 ,
         \60021 , \60022 , \60023 , \60024 , \60025 , \60026 , \60027 , \60028 , \60029 , \60030 ,
         \60031 , \60032 , \60033 , \60034 , \60035 , \60036 , \60037 , \60038 , \60039 , \60040 ,
         \60041 , \60042 , \60043 , \60044 , \60045 , \60046 , \60047 , \60048 , \60049 , \60050 ,
         \60051 , \60052 , \60053 , \60054 , \60055 , \60056 , \60057 , \60058 , \60059 , \60060 ,
         \60061 , \60062 , \60063 , \60064 , \60065 , \60066 , \60067 , \60068 , \60069 , \60070 ,
         \60071 , \60072 , \60073 , \60074 , \60075 , \60076 , \60077 , \60078 , \60079 , \60080 ,
         \60081 , \60082 , \60083 , \60084 , \60085 , \60086 , \60087 , \60088 , \60089 , \60090 ,
         \60091 , \60092 , \60093 , \60094 , \60095 , \60096 , \60097 , \60098 , \60099 , \60100 ,
         \60101 , \60102 , \60103 , \60104 , \60105 , \60106 , \60107 , \60108 , \60109 , \60110 ,
         \60111 , \60112 , \60113 , \60114 , \60115 , \60116 , \60117 , \60118 , \60119 , \60120 ,
         \60121 , \60122 , \60123 , \60124 , \60125 , \60126 , \60127 , \60128 , \60129 , \60130 ,
         \60131 , \60132 , \60133 , \60134 , \60135 , \60136 , \60137 , \60138 , \60139 , \60140 ,
         \60141 , \60142 , \60143 , \60144 , \60145 , \60146 , \60147 , \60148 , \60149 , \60150 ,
         \60151 , \60152 , \60153 , \60154 , \60155 , \60156 , \60157 , \60158 , \60159 , \60160 ,
         \60161 , \60162 , \60163 , \60164 , \60165 , \60166 , \60167 , \60168 , \60169 , \60170 ,
         \60171 , \60172 , \60173 , \60174 , \60175 , \60176 , \60177 , \60178 , \60179 , \60180 ,
         \60181 , \60182 , \60183 , \60184 , \60185 , \60186 , \60187 , \60188 , \60189 , \60190 ,
         \60191 , \60192 , \60193 , \60194 , \60195 , \60196 , \60197 , \60198 , \60199 , \60200 ,
         \60201 , \60202 , \60203 , \60204 , \60205 , \60206 , \60207 , \60208 , \60209 , \60210 ,
         \60211 , \60212 , \60213 , \60214 , \60215 , \60216 , \60217 , \60218 , \60219 , \60220 ,
         \60221 , \60222 , \60223 , \60224 , \60225 , \60226 , \60227 , \60228 , \60229 , \60230 ,
         \60231 , \60232 , \60233 , \60234 , \60235 , \60236 , \60237 , \60238 , \60239 , \60240 ,
         \60241 , \60242 , \60243 , \60244 , \60245 , \60246 , \60247 , \60248 , \60249 , \60250 ,
         \60251 , \60252 , \60253 , \60254 , \60255 , \60256 , \60257 , \60258 , \60259 , \60260 ,
         \60261 , \60262 , \60263 , \60264 , \60265 , \60266 , \60267 , \60268 , \60269 , \60270 ,
         \60271 , \60272 , \60273 , \60274 , \60275 , \60276 , \60277 , \60278 , \60279 , \60280 ,
         \60281 , \60282 , \60283 , \60284 , \60285 , \60286 , \60287 , \60288 , \60289 , \60290 ,
         \60291 , \60292 , \60293 , \60294 , \60295 , \60296 , \60297 , \60298 , \60299 , \60300 ,
         \60301 , \60302 , \60303 , \60304 , \60305 , \60306 , \60307 , \60308 , \60309 , \60310 ,
         \60311 , \60312 , \60313 , \60314 , \60315 , \60316 , \60317 , \60318 , \60319 , \60320 ,
         \60321 , \60322 , \60323 , \60324 , \60325 , \60326 , \60327 , \60328 , \60329 , \60330 ,
         \60331 , \60332 , \60333 , \60334 , \60335 , \60336 , \60337 , \60338 , \60339 , \60340 ,
         \60341 , \60342 , \60343 , \60344 , \60345 , \60346 , \60347 , \60348 , \60349 , \60350 ,
         \60351 , \60352 , \60353 , \60354 , \60355 , \60356 , \60357 , \60358 , \60359 , \60360 ,
         \60361 , \60362 , \60363 , \60364 , \60365 , \60366 , \60367 , \60368 , \60369 , \60370 ,
         \60371 , \60372 , \60373 , \60374 , \60375 , \60376 , \60377 , \60378 , \60379 , \60380 ,
         \60381 , \60382 , \60383 , \60384 , \60385 , \60386 , \60387 , \60388 , \60389 , \60390 ,
         \60391 , \60392 , \60393 , \60394 , \60395 , \60396 , \60397 , \60398 , \60399 , \60400 ,
         \60401 , \60402 , \60403 , \60404 , \60405 , \60406 , \60407 , \60408 , \60409 , \60410 ,
         \60411 , \60412 , \60413 , \60414 , \60415 , \60416 , \60417 , \60418 , \60419 , \60420 ,
         \60421 , \60422 , \60423 , \60424 , \60425 , \60426 , \60427 , \60428 , \60429 , \60430 ,
         \60431 , \60432 , \60433 , \60434 , \60435 , \60436 , \60437 , \60438 , \60439 , \60440 ,
         \60441 , \60442 , \60443 , \60444 , \60445 , \60446 , \60447 , \60448 , \60449 , \60450 ,
         \60451 , \60452 , \60453 , \60454 , \60455 , \60456 , \60457 , \60458 , \60459 , \60460 ,
         \60461 , \60462 , \60463 , \60464 , \60465 , \60466 , \60467 , \60468 , \60469 , \60470 ,
         \60471 , \60472 , \60473 , \60474 , \60475 , \60476 , \60477 , \60478 , \60479 , \60480 ,
         \60481 , \60482 , \60483 , \60484 , \60485 , \60486 , \60487 , \60488 , \60489 , \60490 ,
         \60491 , \60492 , \60493 , \60494 , \60495 , \60496 , \60497 , \60498 , \60499 , \60500 ,
         \60501 , \60502 , \60503 , \60504 , \60505 , \60506 , \60507 , \60508 , \60509 , \60510 ,
         \60511 , \60512 , \60513 , \60514 , \60515 , \60516 , \60517 , \60518 , \60519 , \60520 ,
         \60521 , \60522 , \60523 , \60524 , \60525 , \60526 , \60527 , \60528 , \60529 , \60530 ,
         \60531 , \60532 , \60533 , \60534 , \60535 , \60536 , \60537 , \60538 , \60539 , \60540 ,
         \60541 , \60542 , \60543 , \60544 , \60545 , \60546 , \60547 , \60548 , \60549 , \60550 ,
         \60551 , \60552 , \60553 , \60554 , \60555 , \60556 , \60557 , \60558 , \60559 , \60560 ,
         \60561 , \60562 , \60563 , \60564 , \60565 , \60566 , \60567 , \60568 , \60569 , \60570 ,
         \60571 , \60572 , \60573 , \60574 , \60575 , \60576 , \60577 , \60578 , \60579 , \60580 ,
         \60581 , \60582 , \60583 , \60584 , \60585 , \60586 , \60587 , \60588 , \60589 , \60590 ,
         \60591 , \60592 , \60593 , \60594 , \60595 , \60596 , \60597 , \60598 , \60599 , \60600 ,
         \60601 , \60602 , \60603 , \60604 , \60605 , \60606 , \60607 , \60608 , \60609 , \60610 ,
         \60611 , \60612 , \60613 , \60614 , \60615 , \60616 , \60617 , \60618 , \60619 , \60620 ,
         \60621 , \60622 , \60623 , \60624 , \60625 , \60626 , \60627 , \60628 , \60629 , \60630 ,
         \60631 , \60632 , \60633 , \60634 , \60635 , \60636 , \60637 , \60638 , \60639 , \60640 ,
         \60641 , \60642 , \60643 , \60644 , \60645 , \60646 , \60647 , \60648 , \60649 , \60650 ,
         \60651 , \60652 , \60653 , \60654 , \60655 , \60656 , \60657 , \60658 , \60659 , \60660 ,
         \60661 , \60662 , \60663 , \60664 , \60665 , \60666 , \60667 , \60668 , \60669 , \60670 ,
         \60671 , \60672 , \60673 , \60674 , \60675 , \60676 , \60677 , \60678 , \60679 , \60680 ,
         \60681 , \60682 , \60683 , \60684 , \60685 , \60686 , \60687 , \60688 , \60689 , \60690 ,
         \60691 , \60692 , \60693 , \60694 , \60695 , \60696 , \60697 , \60698 , \60699 , \60700 ,
         \60701 , \60702 , \60703 , \60704 , \60705 , \60706 , \60707 , \60708 , \60709 , \60710 ,
         \60711 , \60712 , \60713 , \60714 , \60715 , \60716 , \60717 , \60718 , \60719 , \60720 ,
         \60721 , \60722 , \60723 , \60724 , \60725 , \60726 , \60727 , \60728 , \60729 , \60730 ,
         \60731 , \60732 , \60733 , \60734 , \60735 , \60736 , \60737 , \60738 , \60739 , \60740 ,
         \60741 , \60742 , \60743 , \60744 , \60745 , \60746 , \60747 , \60748 , \60749 , \60750 ,
         \60751 , \60752 , \60753 , \60754 , \60755 , \60756 , \60757 , \60758 , \60759 , \60760 ,
         \60761 , \60762 , \60763 , \60764 , \60765 , \60766 , \60767 , \60768 , \60769 , \60770 ,
         \60771 , \60772 , \60773 , \60774 , \60775 , \60776 , \60777 , \60778 , \60779 , \60780 ,
         \60781 , \60782 , \60783 , \60784 , \60785 , \60786 , \60787 , \60788 , \60789 , \60790 ,
         \60791 , \60792 , \60793 , \60794 , \60795 , \60796 , \60797 , \60798 , \60799 , \60800 ,
         \60801 , \60802 , \60803 , \60804 , \60805 , \60806 , \60807 , \60808 , \60809 , \60810 ,
         \60811 , \60812 , \60813 , \60814 , \60815 , \60816 , \60817 , \60818 , \60819 , \60820 ,
         \60821 , \60822 , \60823 , \60824 , \60825 , \60826 , \60827 , \60828 , \60829 , \60830 ,
         \60831 , \60832 , \60833 , \60834 , \60835 , \60836 , \60837 , \60838 , \60839 , \60840 ,
         \60841 , \60842 , \60843 , \60844 , \60845 , \60846 , \60847 , \60848 , \60849 , \60850 ,
         \60851 , \60852 , \60853 , \60854 , \60855 , \60856 , \60857 , \60858 , \60859 , \60860 ,
         \60861 , \60862 , \60863 , \60864 , \60865 , \60866 , \60867 , \60868 , \60869 , \60870 ,
         \60871 , \60872 , \60873 , \60874 , \60875 , \60876 , \60877 , \60878 , \60879 , \60880 ,
         \60881 , \60882 , \60883 , \60884 , \60885 , \60886 , \60887 , \60888 , \60889 , \60890 ,
         \60891 , \60892 , \60893 , \60894 , \60895 , \60896 , \60897 , \60898 , \60899 , \60900 ,
         \60901 , \60902 , \60903 , \60904 , \60905 , \60906 , \60907 , \60908 , \60909 , \60910 ,
         \60911 , \60912 , \60913 , \60914 , \60915 , \60916 , \60917 , \60918 , \60919 , \60920 ,
         \60921 , \60922 , \60923 , \60924 , \60925 , \60926 , \60927 , \60928 , \60929 , \60930 ,
         \60931 , \60932 , \60933 , \60934 , \60935 , \60936 , \60937 , \60938 , \60939 , \60940 ,
         \60941 , \60942 , \60943 , \60944 , \60945 , \60946 , \60947 , \60948 , \60949 , \60950 ,
         \60951 , \60952 , \60953 , \60954 , \60955 , \60956 , \60957 , \60958 , \60959 , \60960 ,
         \60961 , \60962 , \60963 , \60964 , \60965 , \60966 , \60967 , \60968 , \60969 , \60970 ,
         \60971 , \60972 , \60973 , \60974 , \60975 , \60976 , \60977 , \60978 , \60979 , \60980 ,
         \60981 , \60982 , \60983 , \60984 , \60985 , \60986 , \60987 , \60988 , \60989 , \60990 ,
         \60991 , \60992 , \60993 , \60994 , \60995 , \60996 , \60997 , \60998 , \60999 , \61000 ,
         \61001 , \61002 , \61003 , \61004 , \61005 , \61006 , \61007 , \61008 , \61009 , \61010 ,
         \61011 , \61012 , \61013 , \61014 , \61015 , \61016 , \61017 , \61018 , \61019 , \61020 ,
         \61021 , \61022 , \61023 , \61024 , \61025 , \61026 , \61027 , \61028 , \61029 , \61030 ,
         \61031 , \61032 , \61033 , \61034 , \61035 , \61036 , \61037 , \61038 , \61039 , \61040 ,
         \61041 , \61042 , \61043 , \61044 , \61045 , \61046 , \61047 , \61048 , \61049 , \61050 ,
         \61051 , \61052 , \61053 , \61054 , \61055 , \61056 , \61057 , \61058 , \61059 , \61060 ,
         \61061 , \61062 , \61063 , \61064 , \61065 , \61066 , \61067 , \61068 , \61069 , \61070 ,
         \61071 , \61072 , \61073 , \61074 , \61075 , \61076 , \61077 , \61078 , \61079 , \61080 ,
         \61081 , \61082 , \61083 , \61084 , \61085 , \61086 , \61087 , \61088 , \61089 , \61090 ,
         \61091 , \61092 , \61093 , \61094 , \61095 , \61096 , \61097 , \61098 , \61099 , \61100 ,
         \61101 , \61102 , \61103 , \61104 , \61105 , \61106 , \61107 , \61108 , \61109 , \61110 ,
         \61111 , \61112 , \61113 , \61114 , \61115 , \61116 , \61117 , \61118 , \61119 , \61120 ,
         \61121 , \61122 , \61123 , \61124 , \61125 , \61126 , \61127 , \61128 , \61129 , \61130 ,
         \61131 , \61132 , \61133 , \61134 , \61135 , \61136 , \61137 , \61138 , \61139 , \61140 ,
         \61141 , \61142 , \61143 , \61144 , \61145 , \61146 , \61147 , \61148 , \61149 , \61150 ,
         \61151 , \61152 , \61153 , \61154 , \61155 , \61156 , \61157 , \61158 , \61159 , \61160 ,
         \61161 , \61162 , \61163 , \61164 , \61165 , \61166 , \61167 , \61168 , \61169 , \61170 ,
         \61171 , \61172 , \61173 , \61174 , \61175 , \61176 , \61177 , \61178 , \61179 , \61180 ,
         \61181 , \61182 , \61183 , \61184 , \61185 , \61186 , \61187 , \61188 , \61189 , \61190 ,
         \61191 , \61192 , \61193 , \61194 , \61195 , \61196 , \61197 , \61198 , \61199 , \61200 ,
         \61201 , \61202 , \61203 , \61204 , \61205 , \61206 , \61207 , \61208 , \61209 , \61210 ,
         \61211 , \61212 , \61213 , \61214 , \61215 , \61216 , \61217 , \61218 , \61219 , \61220 ,
         \61221 , \61222 , \61223 , \61224 , \61225 , \61226 , \61227 , \61228 , \61229 , \61230 ,
         \61231 , \61232 , \61233 , \61234 , \61235 , \61236 , \61237 , \61238 , \61239 , \61240 ,
         \61241 , \61242 , \61243 , \61244 , \61245 , \61246 , \61247 , \61248 , \61249 , \61250 ,
         \61251 , \61252 , \61253 , \61254 , \61255 , \61256 , \61257 , \61258 , \61259 , \61260 ,
         \61261 , \61262 , \61263 , \61264 , \61265 , \61266 , \61267 , \61268 , \61269 , \61270 ,
         \61271 , \61272 , \61273 , \61274 , \61275 , \61276 , \61277 , \61278 , \61279 , \61280 ,
         \61281 , \61282 , \61283 , \61284 , \61285 , \61286 , \61287 , \61288 , \61289 , \61290 ,
         \61291 , \61292 , \61293 , \61294 , \61295 , \61296 , \61297 , \61298 , \61299 , \61300 ,
         \61301 , \61302 , \61303 , \61304 , \61305 , \61306 , \61307 , \61308 , \61309 , \61310 ,
         \61311 , \61312 , \61313 , \61314 , \61315 , \61316 , \61317 , \61318 , \61319 , \61320 ,
         \61321 , \61322 , \61323 , \61324 , \61325 , \61326 , \61327 , \61328 , \61329 , \61330 ,
         \61331 , \61332 , \61333 , \61334 , \61335 , \61336 , \61337 , \61338 , \61339 , \61340 ,
         \61341 , \61342 , \61343 , \61344 , \61345 , \61346 , \61347 , \61348 , \61349 , \61350 ,
         \61351 , \61352 , \61353 , \61354 , \61355 , \61356 , \61357 , \61358 , \61359 , \61360 ,
         \61361 , \61362 , \61363 , \61364 , \61365 , \61366 , \61367 , \61368 , \61369 , \61370 ,
         \61371 , \61372 , \61373 , \61374 , \61375 , \61376 , \61377 , \61378 , \61379 , \61380 ,
         \61381 , \61382 , \61383 , \61384 , \61385 , \61386 , \61387 , \61388 , \61389 , \61390 ,
         \61391 , \61392 , \61393 , \61394 , \61395 , \61396 , \61397 , \61398 , \61399 , \61400 ,
         \61401 , \61402 , \61403 , \61404 , \61405 , \61406 , \61407 , \61408 , \61409 , \61410 ,
         \61411 , \61412 , \61413 , \61414 , \61415 , \61416 , \61417 , \61418 , \61419 , \61420 ,
         \61421 , \61422 , \61423 , \61424 , \61425 , \61426 , \61427 , \61428 , \61429 , \61430 ,
         \61431 , \61432 , \61433 , \61434 , \61435 , \61436 , \61437 , \61438 , \61439 , \61440 ,
         \61441 , \61442 , \61443 , \61444 , \61445 , \61446 , \61447 , \61448 , \61449 , \61450 ,
         \61451 , \61452 , \61453 , \61454 , \61455 , \61456 , \61457 , \61458 , \61459 , \61460 ,
         \61461 , \61462 , \61463 , \61464 , \61465 , \61466 , \61467 , \61468 , \61469 , \61470 ,
         \61471 , \61472 , \61473 , \61474 , \61475 , \61476 , \61477 , \61478 , \61479 , \61480 ,
         \61481 , \61482 , \61483 , \61484 , \61485 , \61486 , \61487 , \61488 , \61489 , \61490 ,
         \61491 , \61492 , \61493 , \61494 , \61495 , \61496 , \61497 , \61498 , \61499 , \61500 ,
         \61501 , \61502 , \61503 , \61504 , \61505 , \61506 , \61507 , \61508 , \61509 , \61510 ,
         \61511 , \61512 , \61513 , \61514 , \61515 , \61516 , \61517 , \61518 , \61519 , \61520 ,
         \61521 , \61522 , \61523 , \61524 , \61525 , \61526 , \61527 , \61528 , \61529 , \61530 ,
         \61531 , \61532 , \61533 , \61534 , \61535 , \61536 , \61537 , \61538 , \61539 , \61540 ,
         \61541 , \61542 , \61543 , \61544 , \61545 , \61546 , \61547 , \61548 , \61549 , \61550 ,
         \61551 , \61552 , \61553 , \61554 , \61555 , \61556 , \61557 , \61558 , \61559 , \61560 ,
         \61561 , \61562 , \61563 , \61564 , \61565 , \61566 , \61567 , \61568 , \61569 , \61570 ,
         \61571 , \61572 , \61573 , \61574 , \61575 , \61576 , \61577 , \61578 , \61579 , \61580 ,
         \61581 , \61582 , \61583 , \61584 , \61585 , \61586 , \61587 , \61588 , \61589 , \61590 ,
         \61591 , \61592 , \61593 , \61594 , \61595 , \61596 , \61597 , \61598 , \61599 , \61600 ,
         \61601 , \61602 , \61603 , \61604 , \61605 , \61606 , \61607 , \61608 , \61609 , \61610 ,
         \61611 , \61612 , \61613 , \61614 , \61615 , \61616 , \61617 , \61618 , \61619 , \61620 ,
         \61621 , \61622 , \61623 , \61624 , \61625 , \61626 , \61627 , \61628 , \61629 , \61630 ,
         \61631 , \61632 , \61633 , \61634 , \61635 , \61636 , \61637 , \61638 , \61639 , \61640 ,
         \61641 , \61642 , \61643 , \61644 , \61645 , \61646 , \61647 , \61648 , \61649 , \61650 ,
         \61651 , \61652 , \61653 , \61654 , \61655 , \61656 , \61657 , \61658 , \61659 , \61660 ,
         \61661 , \61662 , \61663 , \61664 , \61665 , \61666 , \61667 , \61668 , \61669 , \61670 ,
         \61671 , \61672 , \61673 , \61674 , \61675 , \61676 , \61677 , \61678 , \61679 , \61680 ,
         \61681 , \61682 , \61683 , \61684 , \61685 , \61686 , \61687 , \61688 , \61689 , \61690 ,
         \61691 , \61692 , \61693 , \61694 , \61695 , \61696 , \61697 , \61698 , \61699 , \61700 ,
         \61701 , \61702 , \61703 , \61704 , \61705 , \61706 , \61707 , \61708 , \61709 , \61710 ,
         \61711 , \61712 , \61713 , \61714 , \61715 , \61716 , \61717 , \61718 , \61719 , \61720 ,
         \61721 , \61722 , \61723 , \61724 , \61725 , \61726 , \61727 , \61728 , \61729 , \61730 ,
         \61731 , \61732 , \61733 , \61734 , \61735 , \61736 , \61737 , \61738 , \61739 , \61740 ,
         \61741 , \61742 , \61743 , \61744 , \61745 , \61746 , \61747 , \61748 , \61749 , \61750 ,
         \61751 , \61752 , \61753 , \61754 , \61755 , \61756 , \61757 , \61758 , \61759 , \61760 ,
         \61761 , \61762 , \61763 , \61764 , \61765 , \61766 , \61767 , \61768 , \61769 , \61770 ,
         \61771 , \61772 , \61773 , \61774 , \61775 , \61776 , \61777 , \61778 , \61779 , \61780 ,
         \61781 , \61782 , \61783 , \61784 , \61785 , \61786 , \61787 , \61788 , \61789 , \61790 ,
         \61791 , \61792 , \61793 , \61794 , \61795 , \61796 , \61797 , \61798 , \61799 , \61800 ,
         \61801 , \61802 , \61803 , \61804 , \61805 , \61806 , \61807 , \61808 , \61809 , \61810 ,
         \61811 , \61812 , \61813 , \61814 , \61815 , \61816 , \61817 , \61818 , \61819 , \61820 ,
         \61821 , \61822 , \61823 , \61824 , \61825 , \61826 , \61827 , \61828 , \61829 , \61830 ,
         \61831 , \61832 , \61833 , \61834 , \61835 , \61836 , \61837 , \61838 , \61839 , \61840 ,
         \61841 , \61842 , \61843 , \61844 , \61845 , \61846 , \61847 , \61848 , \61849 , \61850 ,
         \61851 , \61852 , \61853 , \61854 , \61855 , \61856 , \61857 , \61858 , \61859 , \61860 ,
         \61861 , \61862 , \61863 , \61864 , \61865 , \61866 , \61867 , \61868 , \61869 , \61870 ,
         \61871 , \61872 , \61873 , \61874 , \61875 , \61876 , \61877 , \61878 , \61879 , \61880 ,
         \61881 , \61882 , \61883 , \61884 , \61885 , \61886 , \61887 , \61888 , \61889 , \61890 ,
         \61891 , \61892 , \61893 , \61894 , \61895 , \61896 , \61897 , \61898 , \61899 , \61900 ,
         \61901 , \61902 , \61903 , \61904 , \61905 , \61906 , \61907 , \61908 , \61909 , \61910 ,
         \61911 , \61912 , \61913 , \61914 , \61915 , \61916 , \61917 , \61918 , \61919 , \61920 ,
         \61921 , \61922 , \61923 , \61924 , \61925 , \61926 , \61927 , \61928 , \61929 , \61930 ,
         \61931 , \61932 , \61933 , \61934 , \61935 , \61936 , \61937 , \61938 , \61939 , \61940 ,
         \61941 , \61942 , \61943 , \61944 , \61945 , \61946 , \61947 , \61948 , \61949 , \61950 ,
         \61951 , \61952 , \61953 , \61954 , \61955 , \61956 , \61957 , \61958 , \61959 , \61960 ,
         \61961 , \61962 , \61963 , \61964 , \61965 , \61966 , \61967 , \61968 , \61969 , \61970 ,
         \61971 , \61972 , \61973 , \61974 , \61975 , \61976 , \61977 , \61978 , \61979 , \61980 ,
         \61981 , \61982 , \61983 , \61984 , \61985 , \61986 , \61987 , \61988 , \61989 , \61990 ,
         \61991 , \61992 , \61993 , \61994 , \61995 , \61996 , \61997 , \61998 , \61999 , \62000 ,
         \62001 , \62002 , \62003 , \62004 , \62005 , \62006 , \62007 , \62008 , \62009 , \62010 ,
         \62011 , \62012 , \62013 , \62014 , \62015 , \62016 , \62017 , \62018 , \62019 , \62020 ,
         \62021 , \62022 , \62023 , \62024 , \62025 , \62026 , \62027 , \62028 , \62029 , \62030 ,
         \62031 , \62032 , \62033 , \62034 , \62035 , \62036 , \62037 , \62038 , \62039 , \62040 ,
         \62041 , \62042 , \62043 , \62044 , \62045 , \62046 , \62047 , \62048 , \62049 , \62050 ,
         \62051 , \62052 , \62053 , \62054 , \62055 , \62056 , \62057 , \62058 , \62059 , \62060 ,
         \62061 , \62062 , \62063 , \62064 , \62065 , \62066 , \62067 , \62068 , \62069 , \62070 ,
         \62071 , \62072 , \62073 , \62074 , \62075 , \62076 , \62077 , \62078 , \62079 , \62080 ,
         \62081 , \62082 , \62083 , \62084 , \62085 , \62086 , \62087 , \62088 , \62089 , \62090 ,
         \62091 , \62092 , \62093 , \62094 , \62095 , \62096 , \62097 , \62098 , \62099 , \62100 ,
         \62101 , \62102 , \62103 , \62104 , \62105 , \62106 , \62107 , \62108 , \62109 , \62110 ,
         \62111 , \62112 , \62113 , \62114 , \62115 , \62116 , \62117 , \62118 , \62119 , \62120 ,
         \62121 , \62122 , \62123 , \62124 , \62125 , \62126 , \62127 , \62128 , \62129 , \62130 ,
         \62131 , \62132 , \62133 , \62134 , \62135 , \62136 , \62137 , \62138 , \62139 , \62140 ,
         \62141 , \62142 , \62143 , \62144 , \62145 , \62146 , \62147 , \62148 , \62149 , \62150 ,
         \62151 , \62152 , \62153 , \62154 , \62155 , \62156 , \62157 , \62158 , \62159 , \62160 ,
         \62161 , \62162 , \62163 , \62164 , \62165 , \62166 , \62167 , \62168 , \62169 , \62170 ,
         \62171 , \62172 , \62173 , \62174 , \62175 , \62176 , \62177 , \62178 , \62179 , \62180 ,
         \62181 , \62182 , \62183 , \62184 , \62185 , \62186 , \62187 , \62188 , \62189 , \62190 ,
         \62191 , \62192 , \62193 , \62194 , \62195 , \62196 , \62197 , \62198 , \62199 , \62200 ,
         \62201 , \62202 , \62203 , \62204 , \62205 , \62206 , \62207 , \62208 , \62209 , \62210 ,
         \62211 , \62212 , \62213 , \62214 , \62215 , \62216 , \62217 , \62218 , \62219 , \62220 ,
         \62221 , \62222 , \62223 , \62224 , \62225 , \62226 , \62227 , \62228 , \62229 , \62230 ,
         \62231 , \62232 , \62233 , \62234 , \62235 , \62236 , \62237 , \62238 , \62239 , \62240 ,
         \62241 , \62242 , \62243 , \62244 , \62245 , \62246 , \62247 , \62248 , \62249 , \62250 ,
         \62251 , \62252 , \62253 , \62254 , \62255 , \62256 , \62257 , \62258 , \62259 , \62260 ,
         \62261 , \62262 , \62263 , \62264 , \62265 , \62266 , \62267 , \62268 , \62269 , \62270 ,
         \62271 , \62272 , \62273 , \62274 , \62275 , \62276 , \62277 , \62278 , \62279 , \62280 ,
         \62281 , \62282 , \62283 , \62284 , \62285 , \62286 , \62287 , \62288 , \62289 , \62290 ,
         \62291 , \62292 , \62293 , \62294 , \62295 , \62296 , \62297 , \62298 , \62299 , \62300 ,
         \62301 , \62302 , \62303 , \62304 , \62305 , \62306 , \62307 , \62308 , \62309 , \62310 ,
         \62311 , \62312 , \62313 , \62314 , \62315 , \62316 , \62317 , \62318 , \62319 , \62320 ,
         \62321 , \62322 , \62323 , \62324 , \62325 , \62326 , \62327 , \62328 , \62329 , \62330 ,
         \62331 , \62332 , \62333 , \62334 , \62335 , \62336 , \62337 , \62338 , \62339 , \62340 ,
         \62341 , \62342 , \62343 , \62344 , \62345 , \62346 , \62347 , \62348 , \62349 , \62350 ,
         \62351 , \62352 , \62353 , \62354 , \62355 , \62356 , \62357 , \62358 , \62359 , \62360 ,
         \62361 , \62362 , \62363 , \62364 , \62365 , \62366 , \62367 , \62368 , \62369 , \62370 ,
         \62371 , \62372 , \62373 , \62374 , \62375 , \62376 , \62377 , \62378 , \62379 , \62380 ,
         \62381 , \62382 , \62383 , \62384 , \62385 , \62386 , \62387 , \62388 , \62389 , \62390 ,
         \62391 , \62392 , \62393 , \62394 , \62395 , \62396 , \62397 , \62398 , \62399 , \62400 ,
         \62401 , \62402 , \62403 , \62404 , \62405 , \62406 , \62407 , \62408 , \62409 , \62410 ,
         \62411 , \62412 , \62413 , \62414 , \62415 , \62416 , \62417 , \62418 , \62419 , \62420 ,
         \62421 , \62422 , \62423 , \62424 , \62425 , \62426 , \62427 , \62428 , \62429 , \62430 ,
         \62431 , \62432 , \62433 , \62434 , \62435 , \62436 , \62437 , \62438 , \62439 , \62440 ,
         \62441 , \62442 , \62443 , \62444 , \62445 , \62446 , \62447 , \62448 , \62449 , \62450 ,
         \62451 , \62452 , \62453 , \62454 , \62455 , \62456 , \62457 , \62458 , \62459 , \62460 ,
         \62461 , \62462 , \62463 , \62464 , \62465 , \62466 , \62467 , \62468 , \62469 , \62470 ,
         \62471 , \62472 , \62473 , \62474 , \62475 , \62476 , \62477 , \62478 , \62479 , \62480 ,
         \62481 , \62482 , \62483 , \62484 , \62485 , \62486 , \62487 , \62488 , \62489 , \62490 ,
         \62491 , \62492 , \62493 , \62494 , \62495 , \62496 , \62497 , \62498 , \62499 , \62500 ,
         \62501 , \62502 , \62503 , \62504 , \62505 , \62506 , \62507 , \62508 , \62509 , \62510 ,
         \62511 , \62512 , \62513 , \62514 , \62515 , \62516 , \62517 , \62518 , \62519 , \62520 ,
         \62521 , \62522 , \62523 , \62524 , \62525 , \62526 , \62527 , \62528 , \62529 , \62530 ,
         \62531 , \62532 , \62533 , \62534 , \62535 , \62536 , \62537 , \62538 , \62539 , \62540 ,
         \62541 , \62542 , \62543 , \62544 , \62545 , \62546 , \62547 , \62548 , \62549 , \62550 ,
         \62551 , \62552 , \62553 , \62554 , \62555 , \62556 , \62557 , \62558 , \62559 , \62560 ,
         \62561 , \62562 , \62563 , \62564 , \62565 , \62566 , \62567 , \62568 , \62569 , \62570 ,
         \62571 , \62572 , \62573 , \62574 , \62575 , \62576 , \62577 , \62578 , \62579 , \62580 ,
         \62581 , \62582 , \62583 , \62584 , \62585 , \62586 , \62587 , \62588 , \62589 , \62590 ,
         \62591 , \62592 , \62593 , \62594 , \62595 , \62596 , \62597 , \62598 , \62599 , \62600 ,
         \62601 , \62602 , \62603 , \62604 , \62605 , \62606 , \62607 , \62608 , \62609 , \62610 ,
         \62611 , \62612 , \62613 , \62614 , \62615 , \62616 , \62617 , \62618 , \62619 , \62620 ,
         \62621 , \62622 , \62623 , \62624 , \62625 , \62626 , \62627 , \62628 , \62629 , \62630 ,
         \62631 , \62632 , \62633 , \62634 , \62635 , \62636 , \62637 , \62638 , \62639 , \62640 ,
         \62641 , \62642 , \62643 , \62644 , \62645 , \62646 , \62647 , \62648 , \62649 , \62650 ,
         \62651 , \62652 , \62653 , \62654 , \62655 , \62656 , \62657 , \62658 , \62659 , \62660 ,
         \62661 , \62662 , \62663 , \62664 , \62665 , \62666 , \62667 , \62668 , \62669 , \62670 ,
         \62671 , \62672 , \62673 , \62674 , \62675 , \62676 , \62677 , \62678 , \62679 , \62680 ,
         \62681 , \62682 , \62683 , \62684 , \62685 , \62686 , \62687 , \62688 , \62689 , \62690 ,
         \62691 , \62692 , \62693 , \62694 , \62695 , \62696 , \62697 , \62698 , \62699 , \62700 ,
         \62701 , \62702 , \62703 , \62704 , \62705 , \62706 , \62707 , \62708 , \62709 , \62710 ,
         \62711 , \62712 , \62713 , \62714 , \62715 , \62716 , \62717 , \62718 , \62719 , \62720 ,
         \62721 , \62722 , \62723 , \62724 , \62725 , \62726 , \62727 , \62728 , \62729 , \62730 ,
         \62731 , \62732 , \62733 , \62734 , \62735 , \62736 , \62737 , \62738 , \62739 , \62740 ,
         \62741 , \62742 , \62743 , \62744 , \62745 , \62746 , \62747 , \62748 , \62749 , \62750 ,
         \62751 , \62752 , \62753 , \62754 , \62755 , \62756 , \62757 , \62758 , \62759 , \62760 ,
         \62761 , \62762 , \62763 , \62764 , \62765 , \62766 , \62767 , \62768 , \62769 , \62770 ,
         \62771 , \62772 , \62773 , \62774 , \62775 , \62776 , \62777 , \62778 , \62779 , \62780 ,
         \62781 , \62782 , \62783 , \62784 , \62785 , \62786 , \62787 , \62788 , \62789 , \62790 ,
         \62791 , \62792 , \62793 , \62794 , \62795 , \62796 , \62797 , \62798 , \62799 , \62800 ,
         \62801 , \62802 , \62803 , \62804 , \62805 , \62806 , \62807 , \62808 , \62809 , \62810 ,
         \62811 , \62812 , \62813 , \62814 , \62815 , \62816 , \62817 , \62818 , \62819 , \62820 ,
         \62821 , \62822 , \62823 , \62824 , \62825 , \62826 , \62827 , \62828 , \62829 , \62830 ,
         \62831 , \62832 , \62833 , \62834 , \62835 , \62836 , \62837 , \62838 , \62839 , \62840 ,
         \62841 , \62842 , \62843 , \62844 , \62845 , \62846 , \62847 , \62848 , \62849 , \62850 ,
         \62851 , \62852 , \62853 , \62854 , \62855 , \62856 , \62857 , \62858 , \62859 , \62860 ,
         \62861 , \62862 , \62863 , \62864 , \62865 , \62866 , \62867 , \62868 , \62869 , \62870 ,
         \62871 , \62872 , \62873 , \62874 , \62875 , \62876 , \62877 , \62878 , \62879 , \62880 ,
         \62881 , \62882 , \62883 , \62884 , \62885 , \62886 , \62887 , \62888 , \62889 , \62890 ,
         \62891 , \62892 , \62893 , \62894 , \62895 , \62896 , \62897 , \62898 , \62899 , \62900 ,
         \62901 , \62902 , \62903 , \62904 , \62905 , \62906 , \62907 , \62908 , \62909 , \62910 ,
         \62911 , \62912 , \62913 , \62914 , \62915 , \62916 , \62917 , \62918 , \62919 , \62920 ,
         \62921 , \62922 , \62923 , \62924 , \62925 , \62926 , \62927 , \62928 , \62929 , \62930 ,
         \62931 , \62932 , \62933 , \62934 , \62935 , \62936 , \62937 , \62938 , \62939 , \62940 ,
         \62941 , \62942 , \62943 , \62944 , \62945 , \62946 , \62947 , \62948 , \62949 , \62950 ,
         \62951 , \62952 , \62953 , \62954 , \62955 , \62956 , \62957 , \62958 , \62959 , \62960 ,
         \62961 , \62962 , \62963 , \62964 , \62965 , \62966 , \62967 , \62968 , \62969 , \62970 ,
         \62971 , \62972 , \62973 , \62974 , \62975 , \62976 , \62977 , \62978 , \62979 , \62980 ,
         \62981 , \62982 , \62983 , \62984 , \62985 , \62986 , \62987 , \62988 , \62989 , \62990 ,
         \62991 , \62992 , \62993 , \62994 , \62995 , \62996 , \62997 , \62998 , \62999 , \63000 ,
         \63001 , \63002 , \63003 , \63004 , \63005 , \63006 , \63007 , \63008 , \63009 , \63010 ,
         \63011 , \63012 , \63013 , \63014 , \63015 , \63016 , \63017 , \63018 , \63019 , \63020 ,
         \63021 , \63022 , \63023 , \63024 , \63025 , \63026 , \63027 , \63028 , \63029 , \63030 ,
         \63031 , \63032 , \63033 , \63034 , \63035 , \63036 , \63037 , \63038 , \63039 , \63040 ,
         \63041 , \63042 , \63043 , \63044 , \63045 , \63046 , \63047 , \63048 , \63049 , \63050 ,
         \63051 , \63052 , \63053 , \63054 , \63055 , \63056 , \63057 , \63058 , \63059 , \63060 ,
         \63061 , \63062 , \63063 , \63064 , \63065 , \63066 , \63067 , \63068 , \63069 , \63070 ,
         \63071 , \63072 , \63073 , \63074 , \63075 , \63076 , \63077 , \63078 , \63079 , \63080 ,
         \63081 , \63082 , \63083 , \63084 , \63085 , \63086 , \63087 , \63088 , \63089 , \63090 ,
         \63091 , \63092 , \63093 , \63094 , \63095 , \63096 , \63097 , \63098 , \63099 , \63100 ,
         \63101 , \63102 , \63103 , \63104 , \63105 , \63106 , \63107 , \63108 , \63109 , \63110 ,
         \63111 , \63112 , \63113 , \63114 , \63115 , \63116 , \63117 , \63118 , \63119 , \63120 ,
         \63121 , \63122 , \63123 , \63124 , \63125 , \63126 , \63127 , \63128 , \63129 , \63130 ,
         \63131 , \63132 , \63133 , \63134 , \63135 , \63136 , \63137 , \63138 , \63139 , \63140 ,
         \63141 , \63142 , \63143 , \63144 , \63145 , \63146 , \63147 , \63148 , \63149 , \63150 ,
         \63151 , \63152 , \63153 , \63154 , \63155 , \63156 , \63157 , \63158 , \63159 , \63160 ,
         \63161 , \63162 , \63163 , \63164 , \63165 , \63166 , \63167 , \63168 , \63169 , \63170 ,
         \63171 , \63172 , \63173 , \63174 , \63175 , \63176 , \63177 , \63178 , \63179 , \63180 ,
         \63181 , \63182 , \63183 , \63184 , \63185 , \63186 , \63187 , \63188 , \63189 , \63190 ,
         \63191 , \63192 , \63193 , \63194 , \63195 , \63196 , \63197 , \63198 , \63199 , \63200 ,
         \63201 , \63202 , \63203 , \63204 , \63205 , \63206 , \63207 , \63208 , \63209 , \63210 ,
         \63211 , \63212 , \63213 , \63214 , \63215 , \63216 , \63217 , \63218 , \63219 , \63220 ,
         \63221 , \63222 , \63223 , \63224 , \63225 , \63226 , \63227 , \63228 , \63229 , \63230 ,
         \63231 , \63232 , \63233 , \63234 , \63235 , \63236 , \63237 , \63238 , \63239 , \63240 ,
         \63241 , \63242 , \63243 , \63244 , \63245 , \63246 , \63247 , \63248 , \63249 , \63250 ,
         \63251 , \63252 , \63253 , \63254 , \63255 , \63256 , \63257 , \63258 , \63259 , \63260 ,
         \63261 , \63262 , \63263 , \63264 , \63265 , \63266 , \63267 , \63268 , \63269 , \63270 ,
         \63271 , \63272 , \63273 , \63274 , \63275 , \63276 , \63277 , \63278 , \63279 , \63280 ,
         \63281 , \63282 , \63283 , \63284 , \63285 , \63286 , \63287 , \63288 , \63289 , \63290 ,
         \63291 , \63292 , \63293 , \63294 , \63295 , \63296 , \63297 , \63298 , \63299 , \63300 ,
         \63301 , \63302 , \63303 , \63304 , \63305 , \63306 , \63307 , \63308 , \63309 , \63310 ,
         \63311 , \63312 , \63313 , \63314 , \63315 , \63316 , \63317 , \63318 , \63319 , \63320 ,
         \63321 , \63322 , \63323 , \63324 , \63325 , \63326 , \63327 , \63328 , \63329 , \63330 ,
         \63331 , \63332 , \63333 , \63334 , \63335 , \63336 , \63337 , \63338 , \63339 , \63340 ,
         \63341 , \63342 , \63343 , \63344 , \63345 , \63346 , \63347 , \63348 , \63349 , \63350 ,
         \63351 , \63352 , \63353 , \63354 , \63355 , \63356 , \63357 , \63358 , \63359 , \63360 ,
         \63361 , \63362 , \63363 , \63364 , \63365 , \63366 , \63367 , \63368 , \63369 , \63370 ,
         \63371 , \63372 , \63373 , \63374 , \63375 , \63376 , \63377 , \63378 , \63379 , \63380 ,
         \63381 , \63382 , \63383 , \63384 , \63385 , \63386 , \63387 , \63388 , \63389 , \63390 ,
         \63391 , \63392 , \63393 , \63394 , \63395 , \63396 , \63397 , \63398 , \63399 , \63400 ,
         \63401 , \63402 , \63403 , \63404 , \63405 , \63406 , \63407 , \63408 , \63409 , \63410 ,
         \63411 , \63412 , \63413 , \63414 , \63415 , \63416 , \63417 , \63418 , \63419 , \63420 ,
         \63421 , \63422 , \63423 , \63424 , \63425 , \63426 , \63427 , \63428 , \63429 , \63430 ,
         \63431 , \63432 , \63433 , \63434 , \63435 , \63436 , \63437 , \63438 , \63439 , \63440 ,
         \63441 , \63442 , \63443 , \63444 , \63445 , \63446 , \63447 , \63448 , \63449 , \63450 ,
         \63451 , \63452 , \63453 , \63454 , \63455 , \63456 , \63457 , \63458 , \63459 , \63460 ,
         \63461 , \63462 , \63463 , \63464 , \63465 , \63466 , \63467 , \63468 , \63469 , \63470 ,
         \63471 , \63472 , \63473 , \63474 , \63475 , \63476 , \63477 , \63478 , \63479 , \63480 ,
         \63481 , \63482 , \63483 , \63484 , \63485 , \63486 , \63487 , \63488 , \63489 , \63490 ,
         \63491 , \63492 , \63493 , \63494 , \63495 , \63496 , \63497 , \63498 , \63499 , \63500 ,
         \63501 , \63502 , \63503 , \63504 , \63505 , \63506 , \63507 , \63508 , \63509 , \63510 ,
         \63511 , \63512 , \63513 , \63514 , \63515 , \63516 , \63517 , \63518 , \63519 , \63520 ,
         \63521 , \63522 , \63523 , \63524 , \63525 , \63526 , \63527 , \63528 , \63529 , \63530 ,
         \63531 , \63532 , \63533 , \63534 , \63535 , \63536 , \63537 , \63538 , \63539 , \63540 ,
         \63541 , \63542 , \63543 , \63544 , \63545 , \63546 , \63547 , \63548 , \63549 , \63550 ,
         \63551 , \63552 , \63553 , \63554 , \63555 , \63556 , \63557 , \63558 , \63559 , \63560 ,
         \63561 , \63562 , \63563 , \63564 , \63565 , \63566 , \63567 , \63568 , \63569 , \63570 ,
         \63571 , \63572 , \63573 , \63574 , \63575 , \63576 , \63577 , \63578 , \63579 , \63580 ,
         \63581 , \63582 , \63583 , \63584 , \63585 , \63586 , \63587 , \63588 , \63589 , \63590 ,
         \63591 , \63592 , \63593 , \63594 , \63595 , \63596 , \63597 , \63598 , \63599 , \63600 ,
         \63601 , \63602 , \63603 , \63604 , \63605 , \63606 , \63607 , \63608 , \63609 , \63610 ,
         \63611 , \63612 , \63613 , \63614 , \63615 , \63616 , \63617 , \63618 , \63619 , \63620 ,
         \63621 , \63622 , \63623 , \63624 , \63625 , \63626 , \63627 , \63628 , \63629 , \63630 ,
         \63631 , \63632 , \63633 , \63634 , \63635 , \63636 , \63637 , \63638 , \63639 , \63640 ,
         \63641 , \63642 , \63643 , \63644 , \63645 , \63646 , \63647 , \63648 , \63649 , \63650 ,
         \63651 , \63652 , \63653 , \63654 , \63655 , \63656 , \63657 , \63658 , \63659 , \63660 ,
         \63661 , \63662 , \63663 , \63664 , \63665 , \63666 , \63667 , \63668 , \63669 , \63670 ,
         \63671 , \63672 , \63673 , \63674 , \63675 , \63676 , \63677 , \63678 , \63679 , \63680 ,
         \63681 , \63682 , \63683 , \63684 , \63685 , \63686 , \63687 , \63688 , \63689 , \63690 ,
         \63691 , \63692 , \63693 , \63694 , \63695 , \63696 , \63697 , \63698 , \63699 , \63700 ,
         \63701 , \63702 , \63703 , \63704 , \63705 , \63706 , \63707 , \63708 , \63709 , \63710 ,
         \63711 , \63712 , \63713 , \63714 , \63715 , \63716 , \63717 , \63718 , \63719 , \63720 ,
         \63721 , \63722 , \63723 , \63724 , \63725 , \63726 , \63727 , \63728 , \63729 , \63730 ,
         \63731 , \63732 , \63733 , \63734 , \63735 , \63736 , \63737 , \63738 , \63739 , \63740 ,
         \63741 , \63742 , \63743 , \63744 , \63745 , \63746 , \63747 , \63748 , \63749 , \63750 ,
         \63751 , \63752 , \63753 , \63754 , \63755 , \63756 , \63757 , \63758 , \63759 , \63760 ,
         \63761 , \63762 , \63763 , \63764 , \63765 , \63766 , \63767 , \63768 , \63769 , \63770 ,
         \63771 , \63772 , \63773 , \63774 , \63775 , \63776 , \63777 , \63778 , \63779 , \63780 ,
         \63781 , \63782 , \63783 , \63784 , \63785 , \63786 , \63787 , \63788 , \63789 , \63790 ,
         \63791 , \63792 , \63793 , \63794 , \63795 , \63796 , \63797 , \63798 , \63799 , \63800 ,
         \63801 , \63802 , \63803 , \63804 , \63805 , \63806 , \63807 , \63808 , \63809 , \63810 ,
         \63811 , \63812 , \63813 , \63814 , \63815 , \63816 , \63817 , \63818 , \63819 , \63820 ,
         \63821 , \63822 , \63823 , \63824 , \63825 , \63826 , \63827 , \63828 , \63829 , \63830 ,
         \63831 , \63832 , \63833 , \63834 , \63835 , \63836 , \63837 , \63838 , \63839 , \63840 ,
         \63841 , \63842 , \63843 , \63844 , \63845 , \63846 , \63847 , \63848 , \63849 , \63850 ,
         \63851 , \63852 , \63853 , \63854 , \63855 , \63856 , \63857 , \63858 , \63859 , \63860 ,
         \63861 , \63862 , \63863 , \63864 , \63865 , \63866 , \63867 , \63868 , \63869 , \63870 ,
         \63871 , \63872 , \63873 , \63874 , \63875 , \63876 , \63877 , \63878 , \63879 , \63880 ,
         \63881 , \63882 , \63883 , \63884 , \63885 , \63886 , \63887 , \63888 , \63889 , \63890 ,
         \63891 , \63892 , \63893 , \63894 , \63895 , \63896 , \63897 , \63898 , \63899 , \63900 ,
         \63901 , \63902 , \63903 , \63904 , \63905 , \63906 , \63907 , \63908 , \63909 , \63910 ,
         \63911 , \63912 , \63913 , \63914 , \63915 , \63916 , \63917 , \63918 , \63919 , \63920 ,
         \63921 , \63922 , \63923 , \63924 , \63925 , \63926 , \63927 , \63928 , \63929 , \63930 ,
         \63931 , \63932 , \63933 , \63934 , \63935 , \63936 , \63937 , \63938 , \63939 , \63940 ,
         \63941 , \63942 , \63943 , \63944 , \63945 , \63946 , \63947 , \63948 , \63949 , \63950 ,
         \63951 , \63952 , \63953 , \63954 , \63955 , \63956 , \63957 , \63958 , \63959 , \63960 ,
         \63961 , \63962 , \63963 , \63964 , \63965 , \63966 , \63967 , \63968 , \63969 , \63970 ,
         \63971 , \63972 , \63973 , \63974 , \63975 , \63976 , \63977 , \63978 , \63979 , \63980 ,
         \63981 , \63982 , \63983 , \63984 , \63985 , \63986 , \63987 , \63988 , \63989 , \63990 ,
         \63991 , \63992 , \63993 , \63994 , \63995 , \63996 , \63997 , \63998 , \63999 , \64000 ,
         \64001 , \64002 , \64003 , \64004 , \64005 , \64006 , \64007 , \64008 , \64009 , \64010 ,
         \64011 , \64012 , \64013 , \64014 , \64015 , \64016 , \64017 , \64018 , \64019 , \64020 ,
         \64021 , \64022 , \64023 , \64024 , \64025 , \64026 , \64027 , \64028 , \64029 , \64030 ,
         \64031 , \64032 , \64033 , \64034 , \64035 , \64036 , \64037 , \64038 , \64039 , \64040 ,
         \64041 , \64042 , \64043 , \64044 , \64045 , \64046 , \64047 , \64048 , \64049 , \64050 ,
         \64051 , \64052 , \64053 , \64054 , \64055 , \64056 , \64057 , \64058 , \64059 , \64060 ,
         \64061 , \64062 , \64063 , \64064 , \64065 , \64066 , \64067 , \64068 , \64069 , \64070 ,
         \64071 , \64072 , \64073 , \64074 , \64075 , \64076 , \64077 , \64078 , \64079 , \64080 ,
         \64081 , \64082 , \64083 , \64084 , \64085 , \64086 , \64087 , \64088 , \64089 , \64090 ,
         \64091 , \64092 , \64093 , \64094 , \64095 , \64096 , \64097 , \64098 , \64099 , \64100 ,
         \64101 , \64102 , \64103 , \64104 , \64105 , \64106 , \64107 , \64108 , \64109 , \64110 ,
         \64111 , \64112 , \64113 , \64114 , \64115 , \64116 , \64117 , \64118 , \64119 , \64120 ,
         \64121 , \64122 , \64123 , \64124 , \64125 , \64126 , \64127 , \64128 , \64129 , \64130 ,
         \64131 , \64132 , \64133 , \64134 , \64135 , \64136 , \64137 , \64138 , \64139 , \64140 ,
         \64141 , \64142 , \64143 , \64144 , \64145 , \64146 , \64147 , \64148 , \64149 , \64150 ,
         \64151 , \64152 , \64153 , \64154 , \64155 , \64156 , \64157 , \64158 , \64159 , \64160 ,
         \64161 , \64162 , \64163 , \64164 , \64165 , \64166 , \64167 , \64168 , \64169 , \64170 ,
         \64171 , \64172 , \64173 , \64174 , \64175 , \64176 , \64177 , \64178 , \64179 , \64180 ,
         \64181 , \64182 , \64183 , \64184 , \64185 , \64186 , \64187 , \64188 , \64189 , \64190 ,
         \64191 , \64192 , \64193 , \64194 , \64195 , \64196 , \64197 , \64198 , \64199 , \64200 ,
         \64201 , \64202 , \64203 , \64204 , \64205 , \64206 , \64207 , \64208 , \64209 , \64210 ,
         \64211 , \64212 , \64213 , \64214 , \64215 , \64216 , \64217 , \64218 , \64219 , \64220 ,
         \64221 , \64222 , \64223 , \64224 , \64225 , \64226 , \64227 , \64228 , \64229 , \64230 ,
         \64231 , \64232 , \64233 , \64234 , \64235 , \64236 , \64237 , \64238 , \64239 , \64240 ,
         \64241 , \64242 , \64243 , \64244 , \64245 , \64246 , \64247 , \64248 , \64249 , \64250 ,
         \64251 , \64252 , \64253 , \64254 , \64255 , \64256 , \64257 , \64258 , \64259 , \64260 ,
         \64261 , \64262 , \64263 , \64264 , \64265 , \64266 , \64267 , \64268 , \64269 , \64270 ,
         \64271 , \64272 , \64273 , \64274 , \64275 , \64276 , \64277 , \64278 , \64279 , \64280 ,
         \64281 , \64282 , \64283 , \64284 , \64285 , \64286 , \64287 , \64288 , \64289 , \64290 ,
         \64291 , \64292 , \64293 , \64294 , \64295 , \64296 , \64297 , \64298 , \64299 , \64300 ,
         \64301 , \64302 , \64303 , \64304 , \64305 , \64306 , \64307 , \64308 , \64309 , \64310 ,
         \64311 , \64312 , \64313 , \64314 , \64315 , \64316 , \64317 , \64318 , \64319 , \64320 ,
         \64321 , \64322 , \64323 , \64324 , \64325 , \64326 , \64327 , \64328 , \64329 , \64330 ,
         \64331 , \64332 , \64333 , \64334 , \64335 , \64336 , \64337 , \64338 , \64339 , \64340 ,
         \64341 , \64342 , \64343 , \64344 , \64345 , \64346 , \64347 , \64348 , \64349 , \64350 ,
         \64351 , \64352 , \64353 , \64354 , \64355 , \64356 , \64357 , \64358 , \64359 , \64360 ,
         \64361 , \64362 , \64363 , \64364 , \64365 , \64366 , \64367 , \64368 , \64369 , \64370 ,
         \64371 , \64372 , \64373 , \64374 , \64375 , \64376 , \64377 , \64378 , \64379 , \64380 ,
         \64381 , \64382 , \64383 , \64384 , \64385 , \64386 , \64387 , \64388 , \64389 , \64390 ,
         \64391 , \64392 , \64393 , \64394 , \64395 , \64396 , \64397 , \64398 , \64399 , \64400 ,
         \64401 , \64402 , \64403 , \64404 , \64405 , \64406 , \64407 , \64408 , \64409 , \64410 ,
         \64411 , \64412 , \64413 , \64414 , \64415 , \64416 , \64417 , \64418 , \64419 , \64420 ,
         \64421 , \64422 , \64423 , \64424 , \64425 , \64426 , \64427 , \64428 , \64429 , \64430 ,
         \64431 , \64432 , \64433 , \64434 , \64435 , \64436 , \64437 , \64438 , \64439 , \64440 ,
         \64441 , \64442 , \64443 , \64444 , \64445 , \64446 , \64447 , \64448 , \64449 , \64450 ,
         \64451 , \64452 , \64453 , \64454 , \64455 , \64456 , \64457 , \64458 , \64459 , \64460 ,
         \64461 , \64462 , \64463 , \64464 , \64465 , \64466 , \64467 , \64468 , \64469 , \64470 ,
         \64471 , \64472 , \64473 , \64474 , \64475 , \64476 , \64477 , \64478 , \64479 , \64480 ,
         \64481 , \64482 , \64483 , \64484 , \64485 , \64486 , \64487 , \64488 , \64489 , \64490 ,
         \64491 , \64492 , \64493 , \64494 , \64495 , \64496 , \64497 , \64498 , \64499 , \64500 ,
         \64501 , \64502 , \64503 , \64504 , \64505 , \64506 , \64507 , \64508 , \64509 , \64510 ,
         \64511 , \64512 , \64513 , \64514 , \64515 , \64516 , \64517 , \64518 , \64519 , \64520 ,
         \64521 , \64522 , \64523 , \64524 , \64525 , \64526 , \64527 , \64528 , \64529 , \64530 ,
         \64531 , \64532 , \64533 , \64534 , \64535 , \64536 , \64537 , \64538 , \64539 , \64540 ,
         \64541 , \64542 , \64543 , \64544 , \64545 , \64546 , \64547 , \64548 , \64549 , \64550 ,
         \64551 , \64552 , \64553 , \64554 , \64555 , \64556 , \64557 , \64558 , \64559 , \64560 ,
         \64561 , \64562 , \64563 , \64564 , \64565 , \64566 , \64567 , \64568 , \64569 , \64570 ,
         \64571 , \64572 , \64573 , \64574 , \64575 , \64576 , \64577 , \64578 , \64579 , \64580 ,
         \64581 , \64582 , \64583 , \64584 , \64585 , \64586 , \64587 , \64588 , \64589 , \64590 ,
         \64591 , \64592 , \64593 , \64594 , \64595 , \64596 , \64597 , \64598 , \64599 , \64600 ,
         \64601 , \64602 , \64603 , \64604 , \64605 , \64606 , \64607 , \64608 , \64609 , \64610 ,
         \64611 , \64612 , \64613 , \64614 , \64615 , \64616 , \64617 , \64618 , \64619 , \64620 ,
         \64621 , \64622 , \64623 , \64624 , \64625 , \64626 , \64627 , \64628 , \64629 , \64630 ,
         \64631 , \64632 , \64633 , \64634 , \64635 , \64636 , \64637 , \64638 , \64639 , \64640 ,
         \64641 , \64642 , \64643 , \64644 , \64645 , \64646 , \64647 , \64648 , \64649 , \64650 ,
         \64651 , \64652 , \64653 , \64654 , \64655 , \64656 , \64657 , \64658 , \64659 , \64660 ,
         \64661 , \64662 , \64663 , \64664 , \64665 , \64666 , \64667 , \64668 , \64669 , \64670 ,
         \64671 , \64672 , \64673 , \64674 , \64675 , \64676 , \64677 , \64678 , \64679 , \64680 ,
         \64681 , \64682 , \64683 , \64684 , \64685 , \64686 , \64687 , \64688 , \64689 , \64690 ,
         \64691 , \64692 , \64693 , \64694 , \64695 , \64696 , \64697 , \64698 , \64699 , \64700 ,
         \64701 , \64702 , \64703 , \64704 , \64705 , \64706 , \64707 , \64708 , \64709 , \64710 ,
         \64711 , \64712 , \64713 , \64714 , \64715 , \64716 , \64717 , \64718 , \64719 , \64720 ,
         \64721 , \64722 , \64723 , \64724 , \64725 , \64726 , \64727 , \64728 , \64729 , \64730 ,
         \64731 , \64732 , \64733 , \64734 , \64735 , \64736 , \64737 , \64738 , \64739 , \64740 ,
         \64741 , \64742 , \64743 , \64744 , \64745 , \64746 , \64747 , \64748 , \64749 , \64750 ,
         \64751 , \64752 , \64753 , \64754 , \64755 , \64756 , \64757 , \64758 , \64759 , \64760 ,
         \64761 , \64762 , \64763 , \64764 , \64765 , \64766 , \64767 , \64768 , \64769 , \64770 ,
         \64771 , \64772 , \64773 , \64774 , \64775 , \64776 , \64777 , \64778 , \64779 , \64780 ,
         \64781 , \64782 , \64783 , \64784 , \64785 , \64786 , \64787 , \64788 , \64789 , \64790 ,
         \64791 , \64792 , \64793 , \64794 , \64795 , \64796 , \64797 , \64798 , \64799 , \64800 ,
         \64801 , \64802 , \64803 , \64804 , \64805 , \64806 , \64807 , \64808 , \64809 , \64810 ,
         \64811 , \64812 , \64813 , \64814 , \64815 , \64816 , \64817 , \64818 , \64819 , \64820 ,
         \64821 , \64822 , \64823 , \64824 , \64825 , \64826 , \64827 , \64828 , \64829 , \64830 ,
         \64831 , \64832 , \64833 , \64834 , \64835 , \64836 , \64837 , \64838 , \64839 , \64840 ,
         \64841 , \64842 , \64843 , \64844 , \64845 , \64846 , \64847 , \64848 , \64849 , \64850 ,
         \64851 , \64852 , \64853 , \64854 , \64855 , \64856 , \64857 , \64858 , \64859 , \64860 ,
         \64861 , \64862 , \64863 , \64864 , \64865 , \64866 , \64867 , \64868 , \64869 , \64870 ,
         \64871 , \64872 , \64873 , \64874 , \64875 , \64876 , \64877 , \64878 , \64879 , \64880 ,
         \64881 , \64882 , \64883 , \64884 , \64885 , \64886 , \64887 , \64888 , \64889 , \64890 ,
         \64891 , \64892 , \64893 , \64894 , \64895 , \64896 , \64897 , \64898 , \64899 , \64900 ,
         \64901 , \64902 , \64903 , \64904 , \64905 , \64906 , \64907 , \64908 , \64909 , \64910 ,
         \64911 , \64912 , \64913 , \64914 , \64915 , \64916 , \64917 , \64918 , \64919 , \64920 ,
         \64921 , \64922 , \64923 , \64924 , \64925 , \64926 , \64927 , \64928 , \64929 , \64930 ,
         \64931 , \64932 , \64933 , \64934 , \64935 , \64936 , \64937 , \64938 , \64939 , \64940 ,
         \64941 , \64942 , \64943 , \64944 , \64945 , \64946 , \64947 , \64948 , \64949 , \64950 ,
         \64951 , \64952 , \64953 , \64954 , \64955 , \64956 , \64957 , \64958 , \64959 , \64960 ,
         \64961 , \64962 , \64963 , \64964 , \64965 , \64966 , \64967 , \64968 , \64969 , \64970 ,
         \64971 , \64972 , \64973 , \64974 , \64975 , \64976 , \64977 , \64978 , \64979 , \64980 ,
         \64981 , \64982 , \64983 , \64984 , \64985 , \64986 , \64987 , \64988 , \64989 , \64990 ,
         \64991 , \64992 , \64993 , \64994 , \64995 , \64996 , \64997 , \64998 , \64999 , \65000 ,
         \65001 , \65002 , \65003 , \65004 , \65005 , \65006 , \65007 , \65008 , \65009 , \65010 ,
         \65011 , \65012 , \65013 , \65014 , \65015 , \65016 , \65017 , \65018 , \65019 , \65020_nGff1e ,
         \65021 , \65022 , \65023 , \65024_nGfe5e , \65025 , \65026 , \65027 , \65028 , \65029 , \65030 ,
         \65031 , \65032_nGfcc0 , \65033 , \65034 , \65035 , \65036 , \65037 , \65038 , \65039 , \65040_nGf9d4 ,
         \65041 , \65042 , \65043 , \65044 , \65045 , \65046 , \65047 , \65048_nGf7a2 , \65049 , \65050 ,
         \65051 , \65052 , \65053 , \65054 , \65055 , \65056_nGec11 , \65057 , \65058 , \65059 , \65060 ,
         \65061 , \65062 , \65063 , \65064_nGe638 , \65065 , \65066 , \65067 , \65068_nGe441 , \65069 , \65070 ,
         \65071 , \65072 , \65073 , \65074 , \65075 , \65076_nGe060 , \65077 , \65078 , \65079 , \65080 ,
         \65081 , \65082 , \65083 , \65084_nGd9de , \65085 , \65086 , \65087 , \65088_nGd7a2 , \65089 , \65090 ,
         \65091 , \65092_nGd59f , \65093 , \65094 , \65095 , \65096_nGd368 , \65097 , \65098 , \65099 , \65100 ,
         \65101 , \65102 , \65103 , \65104_nGcebb , \65105 , \65106 , \65107 , \65108_nGcc44 , \65109 , \65110 ,
         \65111 , \65112_nGc9e1 , \65113 , \65114 , \65115 , \65116 , \65117 , \65118 , \65119 , \65120_nGc4a5 ,
         \65121 , \65122 , \65123 , \65124_nGc1e2 , \65125 , \65126 , \65127 , \65128 , \65129 , \65130 ,
         \65131 , \65132_nGbc0f , \65133 , \65134 , \65135 , \65136_nGb8f8 , \65137 , \65138 , \65139 , \65140_nGb5fc ,
         \65141 , \65142 , \65143 , \65144_nGb31e , \65145 , \65146 , \65147 , \65148 , \65149 , \65150 ,
         \65151 , \65152_nGa763 , \65153 , \65154 , \65155 , \65156_nGa455 , \65157 , \65158 , \65159 , \65160_nGa121 ,
         \65161 , \65162 , \65163 , \65164_nG9e06 , \65165 , \65166 , \65167 , \65168_nG9ab5 , \65169 , \65170 ,
         \65171 , \65172 , \65173 , \65174 , \65175 , \65176_nG93cf , \65177 , \65178 , \65179 , \65180 ,
         \65181 , \65182 , \65183 , \65184_nG8c6c , \65185 , \65186 , \65187 , \65188_nG88da , \65189 , \65190 ,
         \65191 , \65192_nG84f5 , \65193 , \65194 , \65195 , \65196_nG80db , \65197 , \65198 , \65199 , \65200_nG7cdd ,
         \65201 , \65202 , \65203 , \65204 , \65205 , \65206 , \65207 , \65208_nG7550 , \65209 , \65210 ,
         \65211 , \65212_nG71d5 , \65213 , \65214 , \65215 , \65216_nG6e56 , \65217 , \65218 , \65219 , \65220_nG6aad ,
         \65221 , \65222 , \65223 , \65224_nG6724 , \65225 , \65226 , \65227 , \65228_nG63c0 , \65229 , \65230 ,
         \65231 , \65232_nG6058 , \65233 , \65234 , \65235 , \65236_nG5ce5 , \65237 , \65238 , \65239 , \65240_nG59a6 ,
         \65241 , \65242 , \65243 , \65244_nG5674 , \65245 , \65246 , \65247 , \65248_nG5358 , \65249 , \65250 ,
         \65251 , \65252_nG5053 , \65253 , \65254 , \65255 , \65256_nG4d41 , \65257 , \65258 , \65259 , \65260_nG4a68 ,
         \65261 , \65262 , \65263 , \65264_nG4793 , \65265 , \65266 , \65267 , \65268_nG44bd , \65269 , \65270 ,
         \65271 , \65272_nG41fa , \65273 , \65274 , \65275 , \65276_nG3f43 , \65277 , \65278 , \65279 , \65280_nG3cb4 ,
         \65281 , \65282 , \65283 , \65284_nG3a4a , \65285 , \65286 , \65287 , \65288_nG37e1 , \65289 , \65290 ,
         \65291 , \65292_nG358f , \65293 , \65294 , \65295 , \65296_nG332f , \65297 , \65298 , \65299 , \65300_nG30bf ,
         \65301 , \65302 , \65303 , \65304_nG2e68 , \65305 , \65306 , \65307 , \65308_nG2bfd , \65309 , \65310 ,
         \65311 , \65312_nG29b2 , \65313 , \65314 , \65315 , \65316_nG276d , \65317 , \65318 , \65319 , \65320_nG2549 ,
         \65321 , \65322 , \65323 , \65324_nG2359 , \65325 , \65326 , \65327 , \65328_nG2175 , \65329 , \65330 ,
         \65331 , \65332_nG1f9c , \65333 , \65334 , \65335 , \65336_nG1dda , \65337 , \65338 , \65339 , \65340_nG1c2e ,
         \65341 , \65342 , \65343 , \65344_nG1a7f , \65345 , \65346 , \65347 , \65348_nG18e2 , \65349 , \65350 ,
         \65351 , \65352_nG173e , \65353 , \65354 , \65355 , \65356_nGff30 , \65357 , \65358 , \65359 , \65360_nGff2d ,
         \65361 , \65362 , \65363 , \65364_nGff2a , \65365 , \65366 , \65367 , \65368_nGff27 , \65369 , \65370 ,
         \65371 , \65372_nGff24 , \65373 , \65374 , \65375 , \65376_nGff21 , \65377 , \65378 , \65379 , \65380_nGec14 ,
         \65381 , \65382 , \65383 , \65384_nGd7a5 , \65385 , \65386 , \65387 , \65388_nGc4a8 , \65389 , \65390 ,
         \65391 , \65392_nGb321 , \65393 , \65394 , \65395 , \65396_nGa458 , \65397 , \65398 , \65399 , \65400_nG93d2 ,
         \65401 , \65402 , \65403 , \65404_nG88dd , \65405 , \65406 , \65407 , \65408_nG7553 , \65409 , \65410 ,
         \65411 , \65412_nG6e59 , \65413 ;
buf \U$labajz6583 ( R_101_8a8e950, \65021 );
buf \U$labajz6584 ( R_102_8a8f868, \65025 );
buf \U$labajz6585 ( R_103_8a8f910, \65033 );
buf \U$labajz6586 ( R_104_8a8f9b8, \65041 );
buf \U$labajz6587 ( R_105_8a8fa60, \65049 );
buf \U$labajz6588 ( R_106_8a8fb08, \65057 );
buf \U$labajz6589 ( R_107_8a8fbb0, \65065 );
buf \U$labajz6590 ( R_108_8a8fc58, \65069 );
buf \U$labajz6591 ( R_109_8a8fd00, \65077 );
buf \U$labajz6592 ( R_10a_8a8fda8, \65085 );
buf \U$labajz6593 ( R_10b_8a8fe50, \65089 );
buf \U$labajz6594 ( R_10c_8a8fef8, \65093 );
buf \U$labajz6595 ( R_10d_8a8ffa0, \65097 );
buf \U$labajz6596 ( R_10e_8a90048, \65105 );
buf \U$labajz6597 ( R_10f_8a900f0, \65109 );
buf \U$labajz6598 ( R_110_8a90198, \65113 );
buf \U$labajz6599 ( R_111_8a90240, \65121 );
buf \U$labajz6600 ( R_112_8a902e8, \65125 );
buf \U$labajz6601 ( R_113_8a90390, \65133 );
buf \U$labajz6602 ( R_114_8a90438, \65137 );
buf \U$labajz6603 ( R_115_8a904e0, \65141 );
buf \U$labajz6604 ( R_116_8a90588, \65145 );
buf \U$labajz6605 ( R_117_8a90630, \65153 );
buf \U$labajz6606 ( R_118_8a906d8, \65157 );
buf \U$labajz6607 ( R_119_8a90780, \65161 );
buf \U$labajz6608 ( R_11a_8a90828, \65165 );
buf \U$labajz6609 ( R_11b_8a908d0, \65169 );
buf \U$labajz6610 ( R_11c_8a90978, \65177 );
buf \U$labajz6611 ( R_11d_8a90a20, \65185 );
buf \U$labajz6612 ( R_11e_8a90ac8, \65189 );
buf \U$labajz6613 ( R_11f_8a90b70, \65193 );
buf \U$labajz6614 ( R_120_8a90c18, \65197 );
buf \U$labajz6615 ( R_121_8a90cc0, \65201 );
buf \U$labajz6616 ( R_122_8a90d68, \65209 );
buf \U$labajz6617 ( R_123_8a90e10, \65213 );
buf \U$labajz6618 ( R_124_8a90eb8, \65217 );
buf \U$labajz6619 ( R_125_8a90f60, \65221 );
buf \U$labajz6620 ( R_126_8a91008, \65225 );
buf \U$labajz6621 ( R_127_8a910b0, \65229 );
buf \U$labajz6622 ( R_128_8a91158, \65233 );
buf \U$labajz6623 ( R_129_8a91200, \65237 );
buf \U$labajz6624 ( R_12a_8a912a8, \65241 );
buf \U$labajz6625 ( R_12b_8a91350, \65245 );
buf \U$labajz6626 ( R_12c_8a913f8, \65249 );
buf \U$labajz6627 ( R_12d_8a914a0, \65253 );
buf \U$labajz6628 ( R_12e_8a91548, \65257 );
buf \U$labajz6629 ( R_12f_8a915f0, \65261 );
buf \U$labajz6630 ( R_130_8a91698, \65265 );
buf \U$labajz6631 ( R_131_8a91740, \65269 );
buf \U$labajz6632 ( R_132_8a917e8, \65273 );
buf \U$labajz6633 ( R_133_8a91890, \65277 );
buf \U$labajz6634 ( R_134_8a91938, \65281 );
buf \U$labajz6635 ( R_135_8a919e0, \65285 );
buf \U$labajz6636 ( R_136_8a91a88, \65289 );
buf \U$labajz6637 ( R_137_8a91b30, \65293 );
buf \U$labajz6638 ( R_138_8a91bd8, \65297 );
buf \U$labajz6639 ( R_139_8a91c80, \65301 );
buf \U$labajz6640 ( R_13a_8a91d28, \65305 );
buf \U$labajz6641 ( R_13b_8a91dd0, \65309 );
buf \U$labajz6642 ( R_13c_8a91e78, \65313 );
buf \U$labajz6643 ( R_13d_8a91f20, \65317 );
buf \U$labajz6644 ( R_13e_8a91fc8, \65321 );
buf \U$labajz6645 ( R_13f_8a92070, \65325 );
buf \U$labajz6646 ( R_140_8a92118, \65329 );
buf \U$labajz6647 ( R_141_8a921c0, \65333 );
buf \U$labajz6648 ( R_142_8a92268, \65337 );
buf \U$labajz6649 ( R_143_8a92310, \65341 );
buf \U$labajz6650 ( R_144_8a923b8, \65345 );
buf \U$labajz6651 ( R_145_8a92460, \65349 );
buf \U$labajz6652 ( R_146_8a92508, \65353 );
buf \U$labajz6653 ( R_147_8a925b0, \65357 );
buf \U$labajz6654 ( R_148_8a92658, \65361 );
buf \U$labajz6655 ( R_149_8a92700, \65365 );
buf \U$labajz6656 ( R_14a_8a927a8, \65369 );
buf \U$labajz6657 ( R_14b_8a92850, \65373 );
buf \U$labajz6658 ( R_14c_8a928f8, \65377 );
buf \U$labajz6659 ( R_14d_8a929a0, \65381 );
buf \U$labajz6660 ( R_14e_8a92a48, \65385 );
buf \U$labajz6661 ( R_14f_8a92af0, \65389 );
buf \U$labajz6662 ( R_150_8a92b98, \65393 );
buf \U$labajz6663 ( R_151_8a92c40, \65397 );
buf \U$labajz6664 ( R_152_8a92ce8, \65401 );
buf \U$labajz6665 ( R_153_8a92d90, \65405 );
buf \U$labajz6666 ( R_154_8a92e38, \65409 );
buf \U$labajz6667 ( R_155_8a92ee0, \65413 );
nand \U$1 ( \344 , RI9871f50_143, RI9871e60_141);
and \U$2 ( \345 , \344 , RI9871ed8_142);
not \U$3 ( \346 , \345 );
and \U$4 ( \347 , RI9871ed8_142, RI9871f50_143);
not \U$5 ( \348 , RI9871e60_141);
nor \U$6 ( \349 , \348 , RI9871f50_143);
not \U$7 ( \350 , RI9871f50_143);
nor \U$8 ( \351 , \350 , RI9871e60_141);
or \U$9 ( \352 , \349 , \351 );
nor \U$10 ( \353 , RI9871ed8_142, RI9871f50_143);
nor \U$11 ( \354 , \347 , \352 , \353 );
and \U$12 ( \355 , \354 , RI986f520_53);
and \U$13 ( \356 , RI986f610_55, \352 );
nor \U$14 ( \357 , \355 , \356 );
not \U$15 ( \358 , \357 );
or \U$16 ( \359 , \346 , \358 );
not \U$17 ( \360 , \345 );
not \U$18 ( \361 , \360 );
or \U$19 ( \362 , \357 , \361 );
nand \U$20 ( \363 , \359 , \362 );
nand \U$21 ( \364 , RI9872220_149, RI9872130_147);
and \U$22 ( \365 , \364 , RI9871d70_139);
not \U$23 ( \366 , \365 );
not \U$24 ( \367 , \366 );
not \U$25 ( \368 , \367 );
and \U$26 ( \369 , RI9871d70_139, RI9872220_149);
not \U$27 ( \370 , RI9872130_147);
nor \U$28 ( \371 , \370 , RI9872220_149);
not \U$29 ( \372 , RI9872220_149);
nor \U$30 ( \373 , \372 , RI9872130_147);
or \U$31 ( \374 , \371 , \373 );
nor \U$32 ( \375 , RI9871d70_139, RI9872220_149);
nor \U$33 ( \376 , \369 , \374 , \375 );
and \U$34 ( \377 , \376 , RI986ddb0_3);
and \U$35 ( \378 , RI986dcc0_1, \374 );
nor \U$36 ( \379 , \377 , \378 );
not \U$37 ( \380 , \379 );
or \U$38 ( \381 , \368 , \380 );
or \U$39 ( \382 , \379 , \367 );
nand \U$40 ( \383 , \381 , \382 );
xor \U$41 ( \384 , \363 , \383 );
nand \U$42 ( \385 , RI9871de8_140, RI9871d70_139);
and \U$43 ( \386 , \385 , RI9871e60_141);
not \U$44 ( \387 , \386 );
and \U$45 ( \388 , RI9871e60_141, RI9871de8_140);
not \U$46 ( \389 , RI9871d70_139);
nor \U$47 ( \390 , \389 , RI9871de8_140);
not \U$48 ( \391 , RI9871de8_140);
nor \U$49 ( \392 , \391 , RI9871d70_139);
or \U$50 ( \393 , \390 , \392 );
nor \U$51 ( \394 , RI9871e60_141, RI9871de8_140);
nor \U$52 ( \395 , \388 , \393 , \394 );
and \U$53 ( \396 , \395 , RI986df90_7);
and \U$54 ( \397 , RI986dea0_5, \393 );
nor \U$55 ( \398 , \396 , \397 );
not \U$56 ( \399 , \398 );
or \U$57 ( \400 , \387 , \399 );
or \U$58 ( \401 , \398 , \386 );
nand \U$59 ( \402 , \400 , \401 );
and \U$60 ( \403 , \384 , \402 );
and \U$61 ( \404 , \363 , \383 );
or \U$62 ( \405 , \403 , \404 );
not \U$63 ( \406 , RI986f8e0_61);
not \U$64 ( \407 , RI9871fc8_144);
nor \U$65 ( \408 , \406 , \407 );
and \U$66 ( \409 , RI9871fc8_144, RI9872040_145);
not \U$67 ( \410 , RI9871ed8_142);
nor \U$68 ( \411 , \410 , RI9872040_145);
not \U$69 ( \412 , RI9872040_145);
nor \U$70 ( \413 , \412 , RI9871ed8_142);
or \U$71 ( \414 , \411 , \413 );
nor \U$72 ( \415 , RI9871fc8_144, RI9872040_145);
nor \U$73 ( \416 , \409 , \414 , \415 );
and \U$74 ( \417 , \416 , RI986f430_51);
and \U$75 ( \418 , RI986f340_49, \414 );
nor \U$76 ( \419 , \417 , \418 );
nand \U$77 ( \420 , RI9872040_145, RI9871ed8_142);
and \U$78 ( \421 , \420 , RI9871fc8_144);
not \U$79 ( \422 , \421 );
and \U$80 ( \423 , \419 , \422 );
not \U$81 ( \424 , \419 );
and \U$82 ( \425 , \424 , \421 );
nor \U$83 ( \426 , \423 , \425 );
and \U$84 ( \427 , \408 , \426 );
and \U$85 ( \428 , \405 , \427 );
not \U$86 ( \429 , \405 );
not \U$87 ( \430 , \427 );
and \U$88 ( \431 , \429 , \430 );
and \U$89 ( \432 , RI9871c80_137, RI9871cf8_138);
not \U$90 ( \433 , RI9871b18_134);
nor \U$91 ( \434 , \433 , RI9871cf8_138);
and \U$92 ( \435 , \433 , RI9871cf8_138);
or \U$93 ( \436 , \434 , \435 );
nor \U$94 ( \437 , RI9871c80_137, RI9871cf8_138);
nor \U$95 ( \438 , \432 , \436 , \437 );
and \U$96 ( \439 , \438 , RI986e260_13);
and \U$97 ( \440 , RI986e350_15, \436 );
nor \U$98 ( \441 , \439 , \440 );
nand \U$99 ( \442 , RI9871cf8_138, RI9871b18_134);
and \U$100 ( \443 , \442 , RI9871c80_137);
not \U$101 ( \444 , \443 );
and \U$102 ( \445 , \441 , \444 );
not \U$103 ( \446 , \441 );
and \U$104 ( \447 , \446 , \443 );
nor \U$105 ( \448 , \445 , \447 );
not \U$106 ( \449 , \448 );
nand \U$107 ( \450 , RI9871c08_136, RI9871b90_135);
and \U$108 ( \451 , \450 , RI9871b18_134);
nand \U$109 ( \452 , \449 , \451 );
nand \U$110 ( \453 , RI98721a8_148, RI9871c80_137);
and \U$111 ( \454 , \453 , RI9872130_147);
not \U$112 ( \455 , \454 );
not \U$113 ( \456 , \455 );
not \U$114 ( \457 , \456 );
and \U$115 ( \458 , RI9872130_147, RI98721a8_148);
not \U$116 ( \459 , RI9871c80_137);
nor \U$117 ( \460 , \459 , RI98721a8_148);
not \U$118 ( \461 , RI98721a8_148);
nor \U$119 ( \462 , \461 , RI9871c80_137);
or \U$120 ( \463 , \460 , \462 );
nor \U$121 ( \464 , RI9872130_147, RI98721a8_148);
nor \U$122 ( \465 , \458 , \463 , \464 );
and \U$123 ( \466 , \465 , RI986e170_11);
and \U$124 ( \467 , RI986e080_9, \463 );
nor \U$125 ( \468 , \466 , \467 );
not \U$126 ( \469 , \468 );
or \U$127 ( \470 , \457 , \469 );
or \U$128 ( \471 , \468 , \456 );
nand \U$129 ( \472 , \470 , \471 );
and \U$130 ( \473 , \452 , \472 );
not \U$131 ( \474 , \451 );
and \U$132 ( \475 , \474 , \448 );
nor \U$133 ( \476 , \473 , \475 );
nor \U$134 ( \477 , \431 , \476 );
nor \U$135 ( \478 , \428 , \477 );
nand \U$136 ( \479 , RI9871fc8_144, RI986f430_51);
not \U$137 ( \480 , \386 );
and \U$138 ( \481 , \395 , RI986dea0_5);
and \U$139 ( \482 , RI986ddb0_3, \393 );
nor \U$140 ( \483 , \481 , \482 );
not \U$141 ( \484 , \483 );
or \U$142 ( \485 , \480 , \484 );
not \U$143 ( \486 , \386 );
not \U$144 ( \487 , \486 );
or \U$145 ( \488 , \483 , \487 );
nand \U$146 ( \489 , \485 , \488 );
not \U$147 ( \490 , \361 );
and \U$148 ( \491 , \354 , RI986f610_55);
and \U$149 ( \492 , RI986df90_7, \352 );
nor \U$150 ( \493 , \491 , \492 );
not \U$151 ( \494 , \493 );
or \U$152 ( \495 , \490 , \494 );
or \U$153 ( \496 , \493 , \361 );
nand \U$154 ( \497 , \495 , \496 );
xor \U$155 ( \498 , \489 , \497 );
and \U$156 ( \499 , \416 , RI986f340_49);
and \U$157 ( \500 , RI986f520_53, \414 );
nor \U$158 ( \501 , \499 , \500 );
and \U$159 ( \502 , \501 , \422 );
not \U$160 ( \503 , \501 );
and \U$161 ( \504 , \503 , \421 );
nor \U$162 ( \505 , \502 , \504 );
xor \U$163 ( \506 , \498 , \505 );
xor \U$164 ( \507 , \479 , \506 );
and \U$165 ( \508 , \376 , RI986dcc0_1);
and \U$166 ( \509 , RI986e170_11, \374 );
nor \U$167 ( \510 , \508 , \509 );
not \U$168 ( \511 , \510 );
not \U$169 ( \512 , \367 );
and \U$170 ( \513 , \511 , \512 );
and \U$171 ( \514 , \510 , \365 );
nor \U$172 ( \515 , \513 , \514 );
not \U$173 ( \516 , \515 );
nand \U$174 ( \517 , RI986e350_15, \438 );
and \U$175 ( \518 , \517 , \443 );
not \U$176 ( \519 , \517 );
and \U$177 ( \520 , \519 , \444 );
nor \U$178 ( \521 , \518 , \520 );
and \U$179 ( \522 , \465 , RI986e080_9);
and \U$180 ( \523 , RI986e260_13, \463 );
nor \U$181 ( \524 , \522 , \523 );
not \U$182 ( \525 , \524 );
not \U$183 ( \526 , \456 );
and \U$184 ( \527 , \525 , \526 );
and \U$185 ( \528 , \524 , \456 );
nor \U$186 ( \529 , \527 , \528 );
xor \U$187 ( \530 , \521 , \529 );
not \U$188 ( \531 , \530 );
or \U$189 ( \532 , \516 , \531 );
or \U$190 ( \533 , \530 , \515 );
nand \U$191 ( \534 , \532 , \533 );
and \U$192 ( \535 , \507 , \534 );
and \U$193 ( \536 , \479 , \506 );
nor \U$194 ( \537 , \535 , \536 );
xor \U$195 ( \538 , \478 , \537 );
and \U$196 ( \539 , \416 , RI986f520_53);
and \U$197 ( \540 , RI986f610_55, \414 );
nor \U$198 ( \541 , \539 , \540 );
and \U$199 ( \542 , \541 , \421 );
not \U$200 ( \543 , \541 );
and \U$201 ( \544 , \543 , \422 );
nor \U$202 ( \545 , \542 , \544 );
and \U$203 ( \546 , \395 , RI986ddb0_3);
and \U$204 ( \547 , RI986dcc0_1, \393 );
nor \U$205 ( \548 , \546 , \547 );
not \U$206 ( \549 , \548 );
not \U$207 ( \550 , \386 );
and \U$208 ( \551 , \549 , \550 );
and \U$209 ( \552 , \548 , \487 );
nor \U$210 ( \553 , \551 , \552 );
xor \U$211 ( \554 , \545 , \553 );
and \U$212 ( \555 , \354 , RI986df90_7);
and \U$213 ( \556 , RI986dea0_5, \352 );
nor \U$214 ( \557 , \555 , \556 );
not \U$215 ( \558 , \557 );
not \U$216 ( \559 , \361 );
and \U$217 ( \560 , \558 , \559 );
and \U$218 ( \561 , \557 , \361 );
nor \U$219 ( \562 , \560 , \561 );
xor \U$220 ( \563 , \554 , \562 );
nand \U$221 ( \564 , RI986f340_49, RI9871fc8_144);
and \U$222 ( \565 , \465 , RI986e260_13);
and \U$223 ( \566 , RI986e350_15, \463 );
nor \U$224 ( \567 , \565 , \566 );
not \U$225 ( \568 , \567 );
not \U$226 ( \569 , \454 );
and \U$227 ( \570 , \568 , \569 );
and \U$228 ( \571 , \567 , \456 );
nor \U$229 ( \572 , \570 , \571 );
xor \U$230 ( \573 , \572 , \443 );
and \U$231 ( \574 , \376 , RI986e170_11);
and \U$232 ( \575 , RI986e080_9, \374 );
nor \U$233 ( \576 , \574 , \575 );
not \U$234 ( \577 , \576 );
not \U$235 ( \578 , \365 );
and \U$236 ( \579 , \577 , \578 );
and \U$237 ( \580 , \576 , \365 );
nor \U$238 ( \581 , \579 , \580 );
xor \U$239 ( \582 , \573 , \581 );
xor \U$240 ( \583 , \564 , \582 );
xor \U$241 ( \584 , \563 , \583 );
and \U$242 ( \585 , \538 , \584 );
and \U$243 ( \586 , \478 , \537 );
nor \U$244 ( \587 , \585 , \586 );
not \U$245 ( \588 , \587 );
xor \U$246 ( \589 , \489 , \497 );
and \U$247 ( \590 , \589 , \505 );
and \U$248 ( \591 , \489 , \497 );
nor \U$249 ( \592 , \590 , \591 );
xor \U$250 ( \593 , \592 , \479 );
not \U$251 ( \594 , \529 );
not \U$252 ( \595 , \515 );
and \U$253 ( \596 , \594 , \595 );
and \U$254 ( \597 , \529 , \515 );
nor \U$255 ( \598 , \597 , \521 );
nor \U$256 ( \599 , \596 , \598 );
and \U$257 ( \600 , \593 , \599 );
and \U$258 ( \601 , \592 , \479 );
or \U$259 ( \602 , \600 , \601 );
and \U$260 ( \603 , \416 , RI986f610_55);
and \U$261 ( \604 , RI986df90_7, \414 );
nor \U$262 ( \605 , \603 , \604 );
and \U$263 ( \606 , \605 , \421 );
not \U$264 ( \607 , \605 );
and \U$265 ( \608 , \607 , \422 );
nor \U$266 ( \609 , \606 , \608 );
nand \U$267 ( \610 , RI9871fc8_144, RI986f520_53);
xor \U$268 ( \611 , \609 , \610 );
and \U$269 ( \612 , \354 , RI986dea0_5);
and \U$270 ( \613 , RI986ddb0_3, \352 );
nor \U$271 ( \614 , \612 , \613 );
not \U$272 ( \615 , \614 );
not \U$273 ( \616 , \345 );
and \U$274 ( \617 , \615 , \616 );
and \U$275 ( \618 , \614 , \345 );
nor \U$276 ( \619 , \617 , \618 );
xor \U$277 ( \620 , \611 , \619 );
xor \U$278 ( \621 , \602 , \620 );
xor \U$279 ( \622 , \545 , \553 );
xor \U$280 ( \623 , \622 , \562 );
and \U$281 ( \624 , \564 , \623 );
xor \U$282 ( \625 , \545 , \553 );
xor \U$283 ( \626 , \625 , \562 );
and \U$284 ( \627 , \582 , \626 );
and \U$285 ( \628 , \564 , \582 );
or \U$286 ( \629 , \624 , \627 , \628 );
xor \U$287 ( \630 , \621 , \629 );
not \U$288 ( \631 , \630 );
or \U$289 ( \632 , \588 , \631 );
or \U$290 ( \633 , \630 , \587 );
nand \U$291 ( \634 , \632 , \633 );
not \U$292 ( \635 , \634 );
xor \U$293 ( \636 , \545 , \553 );
and \U$294 ( \637 , \636 , \562 );
and \U$295 ( \638 , \545 , \553 );
or \U$296 ( \639 , \637 , \638 );
xor \U$297 ( \640 , \572 , \443 );
and \U$298 ( \641 , \640 , \581 );
and \U$299 ( \642 , \572 , \443 );
or \U$300 ( \643 , \641 , \642 );
or \U$301 ( \644 , \639 , \643 );
nand \U$302 ( \645 , \643 , \639 );
nand \U$303 ( \646 , \644 , \645 );
not \U$304 ( \647 , \646 );
not \U$305 ( \648 , \456 );
nand \U$306 ( \649 , RI986e350_15, \465 );
not \U$307 ( \650 , \649 );
or \U$308 ( \651 , \648 , \650 );
or \U$309 ( \652 , \649 , \456 );
nand \U$310 ( \653 , \651 , \652 );
not \U$311 ( \654 , \653 );
and \U$312 ( \655 , \376 , RI986e080_9);
and \U$313 ( \656 , RI986e260_13, \374 );
nor \U$314 ( \657 , \655 , \656 );
not \U$315 ( \658 , \657 );
not \U$316 ( \659 , \367 );
and \U$317 ( \660 , \658 , \659 );
and \U$318 ( \661 , \657 , \365 );
nor \U$319 ( \662 , \660 , \661 );
not \U$320 ( \663 , \662 );
or \U$321 ( \664 , \654 , \663 );
or \U$322 ( \665 , \662 , \653 );
nand \U$323 ( \666 , \664 , \665 );
not \U$324 ( \667 , \666 );
and \U$325 ( \668 , \395 , RI986dcc0_1);
and \U$326 ( \669 , RI986e170_11, \393 );
nor \U$327 ( \670 , \668 , \669 );
not \U$328 ( \671 , \670 );
not \U$329 ( \672 , \386 );
and \U$330 ( \673 , \671 , \672 );
and \U$331 ( \674 , \670 , \386 );
nor \U$332 ( \675 , \673 , \674 );
not \U$333 ( \676 , \675 );
and \U$334 ( \677 , \667 , \676 );
and \U$335 ( \678 , \666 , \675 );
nor \U$336 ( \679 , \677 , \678 );
not \U$337 ( \680 , \679 );
and \U$338 ( \681 , \647 , \680 );
and \U$339 ( \682 , \646 , \679 );
nor \U$340 ( \683 , \681 , \682 );
not \U$341 ( \684 , \683 );
and \U$342 ( \685 , \635 , \684 );
and \U$343 ( \686 , \634 , \683 );
nor \U$344 ( \687 , \685 , \686 );
not \U$345 ( \688 , \687 );
xor \U$346 ( \689 , \478 , \537 );
xor \U$347 ( \690 , \689 , \584 );
xor \U$348 ( \691 , \592 , \479 );
xor \U$349 ( \692 , \691 , \599 );
or \U$350 ( \693 , \690 , \692 );
not \U$351 ( \694 , \692 );
not \U$352 ( \695 , \690 );
or \U$353 ( \696 , \694 , \695 );
not \U$354 ( \697 , \472 );
and \U$355 ( \698 , \448 , \451 );
not \U$356 ( \699 , \448 );
and \U$357 ( \700 , \699 , \474 );
nor \U$358 ( \701 , \698 , \700 );
not \U$359 ( \702 , \701 );
or \U$360 ( \703 , \697 , \702 );
or \U$361 ( \704 , \701 , \472 );
nand \U$362 ( \705 , \703 , \704 );
xor \U$363 ( \706 , \408 , \426 );
xor \U$364 ( \707 , \705 , \706 );
xor \U$365 ( \708 , \363 , \383 );
xor \U$366 ( \709 , \708 , \402 );
and \U$367 ( \710 , \707 , \709 );
and \U$368 ( \711 , \705 , \706 );
or \U$369 ( \712 , \710 , \711 );
and \U$370 ( \713 , \376 , RI986dea0_5);
and \U$371 ( \714 , RI986ddb0_3, \374 );
nor \U$372 ( \715 , \713 , \714 );
not \U$373 ( \716 , \715 );
not \U$374 ( \717 , \365 );
and \U$375 ( \718 , \716 , \717 );
and \U$376 ( \719 , \715 , \367 );
nor \U$377 ( \720 , \718 , \719 );
and \U$378 ( \721 , \395 , RI986f610_55);
and \U$379 ( \722 , RI986df90_7, \393 );
nor \U$380 ( \723 , \721 , \722 );
not \U$381 ( \724 , \723 );
not \U$382 ( \725 , \487 );
and \U$383 ( \726 , \724 , \725 );
and \U$384 ( \727 , \723 , \386 );
nor \U$385 ( \728 , \726 , \727 );
xor \U$386 ( \729 , \720 , \728 );
and \U$387 ( \730 , \354 , RI986f340_49);
and \U$388 ( \731 , RI986f520_53, \352 );
nor \U$389 ( \732 , \730 , \731 );
not \U$390 ( \733 , \732 );
not \U$391 ( \734 , \345 );
and \U$392 ( \735 , \733 , \734 );
and \U$393 ( \736 , \732 , \361 );
nor \U$394 ( \737 , \735 , \736 );
and \U$395 ( \738 , \729 , \737 );
and \U$396 ( \739 , \720 , \728 );
nor \U$397 ( \740 , \738 , \739 );
nand \U$398 ( \741 , RI986f9d0_63, RI9871fc8_144);
and \U$399 ( \742 , \416 , RI986f8e0_61);
and \U$400 ( \743 , RI986f430_51, \414 );
nor \U$401 ( \744 , \742 , \743 );
and \U$402 ( \745 , \744 , \421 );
not \U$403 ( \746 , \744 );
and \U$404 ( \747 , \746 , \422 );
nor \U$405 ( \748 , \745 , \747 );
nand \U$406 ( \749 , \741 , \748 );
xor \U$407 ( \750 , \740 , \749 );
and \U$408 ( \751 , \438 , RI986e080_9);
and \U$409 ( \752 , RI986e260_13, \436 );
nor \U$410 ( \753 , \751 , \752 );
and \U$411 ( \754 , \753 , \443 );
not \U$412 ( \755 , \753 );
and \U$413 ( \756 , \755 , \444 );
nor \U$414 ( \757 , \754 , \756 );
and \U$415 ( \758 , \465 , RI986dcc0_1);
and \U$416 ( \759 , RI986e170_11, \463 );
nor \U$417 ( \760 , \758 , \759 );
not \U$418 ( \761 , \760 );
not \U$419 ( \762 , \456 );
and \U$420 ( \763 , \761 , \762 );
and \U$421 ( \764 , \760 , \454 );
nor \U$422 ( \765 , \763 , \764 );
or \U$423 ( \766 , \757 , \765 );
not \U$424 ( \767 , \765 );
not \U$425 ( \768 , \757 );
or \U$426 ( \769 , \767 , \768 );
and \U$427 ( \770 , RI9871b18_134, RI9871b90_135);
not \U$428 ( \771 , RI9871c08_136);
and \U$429 ( \772 , \771 , RI9871b90_135);
nor \U$430 ( \773 , \771 , RI9871b90_135);
or \U$431 ( \774 , \772 , \773 );
nor \U$432 ( \775 , RI9871b18_134, RI9871b90_135);
nor \U$433 ( \776 , \770 , \774 , \775 );
nand \U$434 ( \777 , RI986e350_15, \776 );
and \U$435 ( \778 , \777 , \474 );
not \U$436 ( \779 , \777 );
and \U$437 ( \780 , \779 , \451 );
nor \U$438 ( \781 , \778 , \780 );
nand \U$439 ( \782 , \769 , \781 );
nand \U$440 ( \783 , \766 , \782 );
and \U$441 ( \784 , \750 , \783 );
and \U$442 ( \785 , \740 , \749 );
or \U$443 ( \786 , \784 , \785 );
xor \U$444 ( \787 , \712 , \786 );
xor \U$445 ( \788 , \479 , \506 );
xor \U$446 ( \789 , \788 , \534 );
and \U$447 ( \790 , \787 , \789 );
and \U$448 ( \791 , \712 , \786 );
or \U$449 ( \792 , \790 , \791 );
nand \U$450 ( \793 , \696 , \792 );
nand \U$451 ( \794 , \693 , \793 );
nand \U$452 ( \795 , \688 , \794 );
not \U$453 ( \796 , \795 );
not \U$454 ( \797 , RI986f610_55);
nor \U$455 ( \798 , \797 , \407 );
not \U$456 ( \799 , \798 );
and \U$457 ( \800 , \796 , \799 );
and \U$458 ( \801 , \795 , \798 );
nor \U$459 ( \802 , \800 , \801 );
not \U$460 ( \803 , \802 );
and \U$461 ( \804 , \465 , RI986e0f8_10);
and \U$462 ( \805 , RI986e2d8_14, \463 );
nor \U$463 ( \806 , \804 , \805 );
not \U$464 ( \807 , \806 );
not \U$465 ( \808 , \456 );
and \U$466 ( \809 , \807 , \808 );
and \U$467 ( \810 , \806 , \454 );
nor \U$468 ( \811 , \809 , \810 );
nand \U$469 ( \812 , RI986e3c8_16, \438 );
and \U$470 ( \813 , \812 , \443 );
not \U$471 ( \814 , \812 );
and \U$472 ( \815 , \814 , \444 );
nor \U$473 ( \816 , \813 , \815 );
xor \U$474 ( \817 , \811 , \816 );
and \U$475 ( \818 , \376 , RI986dd38_2);
and \U$476 ( \819 , RI986e1e8_12, \374 );
nor \U$477 ( \820 , \818 , \819 );
not \U$478 ( \821 , \820 );
not \U$479 ( \822 , \365 );
and \U$480 ( \823 , \821 , \822 );
and \U$481 ( \824 , \820 , \367 );
nor \U$482 ( \825 , \823 , \824 );
xor \U$483 ( \826 , \817 , \825 );
not \U$484 ( \827 , \826 );
nand \U$485 ( \828 , RI986f4a8_52, RI9871fc8_144);
not \U$486 ( \829 , \828 );
not \U$487 ( \830 , \829 );
and \U$488 ( \831 , \827 , \830 );
and \U$489 ( \832 , \826 , \829 );
and \U$490 ( \833 , \416 , RI986f3b8_50);
and \U$491 ( \834 , RI986f598_54, \414 );
nor \U$492 ( \835 , \833 , \834 );
and \U$493 ( \836 , \835 , \421 );
not \U$494 ( \837 , \835 );
and \U$495 ( \838 , \837 , \422 );
nor \U$496 ( \839 , \836 , \838 );
and \U$497 ( \840 , \395 , RI986df18_6);
and \U$498 ( \841 , RI986de28_4, \393 );
nor \U$499 ( \842 , \840 , \841 );
not \U$500 ( \843 , \842 );
not \U$501 ( \844 , \487 );
and \U$502 ( \845 , \843 , \844 );
and \U$503 ( \846 , \842 , \386 );
nor \U$504 ( \847 , \845 , \846 );
xor \U$505 ( \848 , \839 , \847 );
and \U$506 ( \849 , \354 , RI986f688_56);
and \U$507 ( \850 , RI986e008_8, \352 );
nor \U$508 ( \851 , \849 , \850 );
not \U$509 ( \852 , \851 );
not \U$510 ( \853 , \345 );
and \U$511 ( \854 , \852 , \853 );
and \U$512 ( \855 , \851 , \345 );
nor \U$513 ( \856 , \854 , \855 );
xor \U$514 ( \857 , \848 , \856 );
nor \U$515 ( \858 , \832 , \857 );
nor \U$516 ( \859 , \831 , \858 );
not \U$517 ( \860 , \487 );
and \U$518 ( \861 , \395 , RI986e008_8);
and \U$519 ( \862 , RI986df18_6, \393 );
nor \U$520 ( \863 , \861 , \862 );
not \U$521 ( \864 , \863 );
or \U$522 ( \865 , \860 , \864 );
or \U$523 ( \866 , \863 , \386 );
nand \U$524 ( \867 , \865 , \866 );
not \U$525 ( \868 , \365 );
and \U$526 ( \869 , \376 , RI986de28_4);
and \U$527 ( \870 , RI986dd38_2, \374 );
nor \U$528 ( \871 , \869 , \870 );
not \U$529 ( \872 , \871 );
or \U$530 ( \873 , \868 , \872 );
or \U$531 ( \874 , \871 , \365 );
nand \U$532 ( \875 , \873 , \874 );
xor \U$533 ( \876 , \867 , \875 );
not \U$534 ( \877 , \345 );
and \U$535 ( \878 , \354 , RI986f598_54);
and \U$536 ( \879 , RI986f688_56, \352 );
nor \U$537 ( \880 , \878 , \879 );
not \U$538 ( \881 , \880 );
or \U$539 ( \882 , \877 , \881 );
or \U$540 ( \883 , \880 , \345 );
nand \U$541 ( \884 , \882 , \883 );
and \U$542 ( \885 , \876 , \884 );
and \U$543 ( \886 , \867 , \875 );
or \U$544 ( \887 , \885 , \886 );
and \U$545 ( \888 , \438 , RI986e2d8_14);
and \U$546 ( \889 , RI986e3c8_16, \436 );
nor \U$547 ( \890 , \888 , \889 );
and \U$548 ( \891 , \890 , \444 );
not \U$549 ( \892 , \890 );
and \U$550 ( \893 , \892 , \443 );
nor \U$551 ( \894 , \891 , \893 );
xor \U$552 ( \895 , \894 , \474 );
not \U$553 ( \896 , \456 );
and \U$554 ( \897 , \465 , RI986e1e8_12);
and \U$555 ( \898 , RI986e0f8_10, \463 );
nor \U$556 ( \899 , \897 , \898 );
not \U$557 ( \900 , \899 );
or \U$558 ( \901 , \896 , \900 );
or \U$559 ( \902 , \899 , \454 );
nand \U$560 ( \903 , \901 , \902 );
and \U$561 ( \904 , \895 , \903 );
and \U$562 ( \905 , \894 , \474 );
or \U$563 ( \906 , \904 , \905 );
xor \U$564 ( \907 , \887 , \906 );
not \U$565 ( \908 , RI986f958_62);
nor \U$566 ( \909 , \908 , \407 );
and \U$567 ( \910 , \416 , RI986f4a8_52);
and \U$568 ( \911 , RI986f3b8_50, \414 );
nor \U$569 ( \912 , \910 , \911 );
and \U$570 ( \913 , \912 , \422 );
not \U$571 ( \914 , \912 );
and \U$572 ( \915 , \914 , \421 );
nor \U$573 ( \916 , \913 , \915 );
and \U$574 ( \917 , \909 , \916 );
and \U$575 ( \918 , \907 , \917 );
and \U$576 ( \919 , \887 , \906 );
nor \U$577 ( \920 , \918 , \919 );
xor \U$578 ( \921 , \859 , \920 );
and \U$579 ( \922 , \376 , RI986e1e8_12);
and \U$580 ( \923 , RI986e0f8_10, \374 );
nor \U$581 ( \924 , \922 , \923 );
not \U$582 ( \925 , \924 );
not \U$583 ( \926 , \365 );
and \U$584 ( \927 , \925 , \926 );
and \U$585 ( \928 , \924 , \367 );
nor \U$586 ( \929 , \927 , \928 );
xor \U$587 ( \930 , \929 , \443 );
and \U$588 ( \931 , \465 , RI986e2d8_14);
and \U$589 ( \932 , RI986e3c8_16, \463 );
nor \U$590 ( \933 , \931 , \932 );
not \U$591 ( \934 , \933 );
not \U$592 ( \935 , \454 );
and \U$593 ( \936 , \934 , \935 );
and \U$594 ( \937 , \933 , \456 );
nor \U$595 ( \938 , \936 , \937 );
xor \U$596 ( \939 , \930 , \938 );
nand \U$597 ( \940 , RI986f3b8_50, RI9871fc8_144);
and \U$598 ( \941 , \416 , RI986f598_54);
and \U$599 ( \942 , RI986f688_56, \414 );
nor \U$600 ( \943 , \941 , \942 );
and \U$601 ( \944 , \943 , \421 );
not \U$602 ( \945 , \943 );
and \U$603 ( \946 , \945 , \422 );
nor \U$604 ( \947 , \944 , \946 );
and \U$605 ( \948 , \395 , RI986de28_4);
and \U$606 ( \949 , RI986dd38_2, \393 );
nor \U$607 ( \950 , \948 , \949 );
not \U$608 ( \951 , \950 );
not \U$609 ( \952 , \487 );
and \U$610 ( \953 , \951 , \952 );
and \U$611 ( \954 , \950 , \386 );
nor \U$612 ( \955 , \953 , \954 );
xor \U$613 ( \956 , \947 , \955 );
and \U$614 ( \957 , \354 , RI986e008_8);
and \U$615 ( \958 , RI986df18_6, \352 );
nor \U$616 ( \959 , \957 , \958 );
not \U$617 ( \960 , \959 );
not \U$618 ( \961 , \345 );
and \U$619 ( \962 , \960 , \961 );
and \U$620 ( \963 , \959 , \345 );
nor \U$621 ( \964 , \962 , \963 );
xor \U$622 ( \965 , \956 , \964 );
xor \U$623 ( \966 , \940 , \965 );
xor \U$624 ( \967 , \939 , \966 );
and \U$625 ( \968 , \921 , \967 );
and \U$626 ( \969 , \859 , \920 );
or \U$627 ( \970 , \968 , \969 );
xor \U$628 ( \971 , \929 , \443 );
and \U$629 ( \972 , \971 , \938 );
and \U$630 ( \973 , \929 , \443 );
or \U$631 ( \974 , \972 , \973 );
xor \U$632 ( \975 , \947 , \955 );
and \U$633 ( \976 , \975 , \964 );
and \U$634 ( \977 , \947 , \955 );
or \U$635 ( \978 , \976 , \977 );
or \U$636 ( \979 , \974 , \978 );
nand \U$637 ( \980 , \974 , \978 );
nand \U$638 ( \981 , \979 , \980 );
not \U$639 ( \982 , \981 );
and \U$640 ( \983 , \376 , RI986e0f8_10);
and \U$641 ( \984 , RI986e2d8_14, \374 );
nor \U$642 ( \985 , \983 , \984 );
not \U$643 ( \986 , \985 );
not \U$644 ( \987 , \367 );
and \U$645 ( \988 , \986 , \987 );
and \U$646 ( \989 , \985 , \365 );
nor \U$647 ( \990 , \988 , \989 );
nand \U$648 ( \991 , RI986e3c8_16, \465 );
not \U$649 ( \992 , \991 );
not \U$650 ( \993 , \456 );
and \U$651 ( \994 , \992 , \993 );
and \U$652 ( \995 , \991 , \456 );
nor \U$653 ( \996 , \994 , \995 );
xor \U$654 ( \997 , \990 , \996 );
and \U$655 ( \998 , \395 , RI986dd38_2);
and \U$656 ( \999 , RI986e1e8_12, \393 );
nor \U$657 ( \1000 , \998 , \999 );
not \U$658 ( \1001 , \1000 );
not \U$659 ( \1002 , \386 );
and \U$660 ( \1003 , \1001 , \1002 );
and \U$661 ( \1004 , \1000 , \487 );
nor \U$662 ( \1005 , \1003 , \1004 );
xor \U$663 ( \1006 , \997 , \1005 );
not \U$664 ( \1007 , \1006 );
and \U$665 ( \1008 , \982 , \1007 );
and \U$666 ( \1009 , \981 , \1006 );
nor \U$667 ( \1010 , \1008 , \1009 );
xor \U$668 ( \1011 , \970 , \1010 );
xor \U$669 ( \1012 , \839 , \847 );
and \U$670 ( \1013 , \1012 , \856 );
and \U$671 ( \1014 , \839 , \847 );
or \U$672 ( \1015 , \1013 , \1014 );
xor \U$673 ( \1016 , \1015 , \828 );
xor \U$674 ( \1017 , \811 , \816 );
and \U$675 ( \1018 , \1017 , \825 );
and \U$676 ( \1019 , \811 , \816 );
or \U$677 ( \1020 , \1018 , \1019 );
and \U$678 ( \1021 , \1016 , \1020 );
and \U$679 ( \1022 , \1015 , \828 );
or \U$680 ( \1023 , \1021 , \1022 );
and \U$681 ( \1024 , \416 , RI986f688_56);
and \U$682 ( \1025 , RI986e008_8, \414 );
nor \U$683 ( \1026 , \1024 , \1025 );
and \U$684 ( \1027 , \1026 , \421 );
not \U$685 ( \1028 , \1026 );
and \U$686 ( \1029 , \1028 , \422 );
nor \U$687 ( \1030 , \1027 , \1029 );
not \U$688 ( \1031 , \1030 );
not \U$689 ( \1032 , \345 );
and \U$690 ( \1033 , \354 , RI986df18_6);
and \U$691 ( \1034 , RI986de28_4, \352 );
nor \U$692 ( \1035 , \1033 , \1034 );
not \U$693 ( \1036 , \1035 );
or \U$694 ( \1037 , \1032 , \1036 );
or \U$695 ( \1038 , \1035 , \361 );
nand \U$696 ( \1039 , \1037 , \1038 );
not \U$697 ( \1040 , \1039 );
or \U$698 ( \1041 , \1031 , \1040 );
or \U$699 ( \1042 , \1030 , \1039 );
nand \U$700 ( \1043 , \1041 , \1042 );
not \U$701 ( \1044 , \1043 );
nand \U$702 ( \1045 , RI986f598_54, RI9871fc8_144);
not \U$703 ( \1046 , \1045 );
and \U$704 ( \1047 , \1044 , \1046 );
and \U$705 ( \1048 , \1043 , \1045 );
nor \U$706 ( \1049 , \1047 , \1048 );
xor \U$707 ( \1050 , \1023 , \1049 );
xor \U$708 ( \1051 , \929 , \443 );
xor \U$709 ( \1052 , \1051 , \938 );
and \U$710 ( \1053 , \940 , \1052 );
xor \U$711 ( \1054 , \929 , \443 );
xor \U$712 ( \1055 , \1054 , \938 );
and \U$713 ( \1056 , \965 , \1055 );
and \U$714 ( \1057 , \940 , \965 );
or \U$715 ( \1058 , \1053 , \1056 , \1057 );
xor \U$716 ( \1059 , \1050 , \1058 );
and \U$717 ( \1060 , \1011 , \1059 );
and \U$718 ( \1061 , \970 , \1010 );
or \U$719 ( \1062 , \1060 , \1061 );
not \U$720 ( \1063 , \1062 );
not \U$721 ( \1064 , \687 );
not \U$722 ( \1065 , \794 );
and \U$723 ( \1066 , \1064 , \1065 );
and \U$724 ( \1067 , \687 , \794 );
nor \U$725 ( \1068 , \1066 , \1067 );
not \U$726 ( \1069 , \692 );
not \U$727 ( \1070 , \792 );
or \U$728 ( \1071 , \1069 , \1070 );
or \U$729 ( \1072 , \792 , \692 );
nand \U$730 ( \1073 , \1071 , \1072 );
not \U$731 ( \1074 , \1073 );
not \U$732 ( \1075 , \690 );
and \U$733 ( \1076 , \1074 , \1075 );
and \U$734 ( \1077 , \1073 , \690 );
nor \U$735 ( \1078 , \1076 , \1077 );
not \U$736 ( \1079 , \1078 );
not \U$737 ( \1080 , \781 );
not \U$738 ( \1081 , \757 );
or \U$739 ( \1082 , \1080 , \1081 );
or \U$740 ( \1083 , \757 , \781 );
nand \U$741 ( \1084 , \1082 , \1083 );
not \U$742 ( \1085 , \1084 );
not \U$743 ( \1086 , \765 );
and \U$744 ( \1087 , \1085 , \1086 );
and \U$745 ( \1088 , \1084 , \765 );
nor \U$746 ( \1089 , \1087 , \1088 );
xor \U$747 ( \1090 , \720 , \728 );
xor \U$748 ( \1091 , \1090 , \737 );
or \U$749 ( \1092 , \1089 , \1091 );
not \U$750 ( \1093 , \1091 );
not \U$751 ( \1094 , \1089 );
or \U$752 ( \1095 , \1093 , \1094 );
or \U$753 ( \1096 , \748 , \741 );
nand \U$754 ( \1097 , \1096 , \749 );
nand \U$755 ( \1098 , \1095 , \1097 );
nand \U$756 ( \1099 , \1092 , \1098 );
and \U$757 ( \1100 , \354 , RI986f430_51);
and \U$758 ( \1101 , RI986f340_49, \352 );
nor \U$759 ( \1102 , \1100 , \1101 );
not \U$760 ( \1103 , \1102 );
not \U$761 ( \1104 , \345 );
and \U$762 ( \1105 , \1103 , \1104 );
and \U$763 ( \1106 , \1102 , \361 );
nor \U$764 ( \1107 , \1105 , \1106 );
nand \U$765 ( \1108 , RI986f700_57, RI9871fc8_144);
xor \U$766 ( \1109 , \1107 , \1108 );
and \U$767 ( \1110 , \416 , RI986f9d0_63);
and \U$768 ( \1111 , RI986f8e0_61, \414 );
nor \U$769 ( \1112 , \1110 , \1111 );
and \U$770 ( \1113 , \1112 , \421 );
not \U$771 ( \1114 , \1112 );
and \U$772 ( \1115 , \1114 , \422 );
nor \U$773 ( \1116 , \1113 , \1115 );
and \U$774 ( \1117 , \1109 , \1116 );
and \U$775 ( \1118 , \1107 , \1108 );
or \U$776 ( \1119 , \1117 , \1118 );
and \U$777 ( \1120 , \438 , RI986e170_11);
and \U$778 ( \1121 , RI986e080_9, \436 );
nor \U$779 ( \1122 , \1120 , \1121 );
and \U$780 ( \1123 , \1122 , \443 );
not \U$781 ( \1124 , \1122 );
and \U$782 ( \1125 , \1124 , \444 );
nor \U$783 ( \1126 , \1123 , \1125 );
nand \U$784 ( \1127 , RI98718c0_129, RI98720b8_146);
and \U$785 ( \1128 , \1127 , RI9871c08_136);
xor \U$786 ( \1129 , \1126 , \1128 );
and \U$787 ( \1130 , \776 , RI986e260_13);
and \U$788 ( \1131 , RI986e350_15, \774 );
nor \U$789 ( \1132 , \1130 , \1131 );
and \U$790 ( \1133 , \1132 , \451 );
not \U$791 ( \1134 , \1132 );
and \U$792 ( \1135 , \1134 , \474 );
nor \U$793 ( \1136 , \1133 , \1135 );
and \U$794 ( \1137 , \1129 , \1136 );
and \U$795 ( \1138 , \1126 , \1128 );
or \U$796 ( \1139 , \1137 , \1138 );
xor \U$797 ( \1140 , \1119 , \1139 );
and \U$798 ( \1141 , \465 , RI986ddb0_3);
and \U$799 ( \1142 , RI986dcc0_1, \463 );
nor \U$800 ( \1143 , \1141 , \1142 );
not \U$801 ( \1144 , \1143 );
not \U$802 ( \1145 , \456 );
and \U$803 ( \1146 , \1144 , \1145 );
and \U$804 ( \1147 , \1143 , \454 );
nor \U$805 ( \1148 , \1146 , \1147 );
and \U$806 ( \1149 , \376 , RI986df90_7);
and \U$807 ( \1150 , RI986dea0_5, \374 );
nor \U$808 ( \1151 , \1149 , \1150 );
not \U$809 ( \1152 , \1151 );
not \U$810 ( \1153 , \367 );
and \U$811 ( \1154 , \1152 , \1153 );
and \U$812 ( \1155 , \1151 , \367 );
nor \U$813 ( \1156 , \1154 , \1155 );
xor \U$814 ( \1157 , \1148 , \1156 );
and \U$815 ( \1158 , \395 , RI986f520_53);
and \U$816 ( \1159 , RI986f610_55, \393 );
nor \U$817 ( \1160 , \1158 , \1159 );
not \U$818 ( \1161 , \1160 );
not \U$819 ( \1162 , \487 );
and \U$820 ( \1163 , \1161 , \1162 );
and \U$821 ( \1164 , \1160 , \386 );
nor \U$822 ( \1165 , \1163 , \1164 );
and \U$823 ( \1166 , \1157 , \1165 );
and \U$824 ( \1167 , \1148 , \1156 );
or \U$825 ( \1168 , \1166 , \1167 );
and \U$826 ( \1169 , \1140 , \1168 );
and \U$827 ( \1170 , \1119 , \1139 );
nor \U$828 ( \1171 , \1169 , \1170 );
xor \U$829 ( \1172 , \1099 , \1171 );
xor \U$830 ( \1173 , \705 , \706 );
xor \U$831 ( \1174 , \1173 , \709 );
and \U$832 ( \1175 , \1172 , \1174 );
and \U$833 ( \1176 , \1099 , \1171 );
or \U$834 ( \1177 , \1175 , \1176 );
not \U$835 ( \1178 , \427 );
not \U$836 ( \1179 , \476 );
not \U$837 ( \1180 , \405 );
and \U$838 ( \1181 , \1179 , \1180 );
and \U$839 ( \1182 , \476 , \405 );
nor \U$840 ( \1183 , \1181 , \1182 );
not \U$841 ( \1184 , \1183 );
or \U$842 ( \1185 , \1178 , \1184 );
or \U$843 ( \1186 , \1183 , \427 );
nand \U$844 ( \1187 , \1185 , \1186 );
xor \U$845 ( \1188 , \1177 , \1187 );
xor \U$846 ( \1189 , \712 , \786 );
xor \U$847 ( \1190 , \1189 , \789 );
and \U$848 ( \1191 , \1188 , \1190 );
and \U$849 ( \1192 , \1177 , \1187 );
or \U$850 ( \1193 , \1191 , \1192 );
nand \U$851 ( \1194 , \1079 , \1193 );
or \U$852 ( \1195 , \1068 , \1194 );
xnor \U$853 ( \1196 , \1194 , \1068 );
and \U$854 ( \1197 , \416 , RI986e710_23);
and \U$855 ( \1198 , RI986e620_21, \414 );
nor \U$856 ( \1199 , \1197 , \1198 );
and \U$857 ( \1200 , \1199 , \421 );
not \U$858 ( \1201 , \1199 );
and \U$859 ( \1202 , \1201 , \422 );
nor \U$860 ( \1203 , \1200 , \1202 );
not \U$861 ( \1204 , \1203 );
nand \U$862 ( \1205 , RI986e530_19, RI9871fc8_144);
and \U$863 ( \1206 , \416 , RI986e440_17);
and \U$864 ( \1207 , RI986e710_23, \414 );
nor \U$865 ( \1208 , \1206 , \1207 );
and \U$866 ( \1209 , \1208 , \421 );
not \U$867 ( \1210 , \1208 );
and \U$868 ( \1211 , \1210 , \422 );
nor \U$869 ( \1212 , \1209 , \1211 );
nand \U$870 ( \1213 , \1205 , \1212 );
not \U$871 ( \1214 , \1213 );
or \U$872 ( \1215 , \1204 , \1214 );
or \U$873 ( \1216 , \1213 , \1203 );
nand \U$874 ( \1217 , \1215 , \1216 );
not \U$875 ( \1218 , \1217 );
nand \U$876 ( \1219 , RI986e440_17, RI9871fc8_144);
not \U$877 ( \1220 , \1219 );
and \U$878 ( \1221 , \1218 , \1220 );
and \U$879 ( \1222 , \1217 , \1219 );
nor \U$880 ( \1223 , \1221 , \1222 );
and \U$881 ( \1224 , \395 , RI986f700_57);
and \U$882 ( \1225 , RI986f9d0_63, \393 );
nor \U$883 ( \1226 , \1224 , \1225 );
not \U$884 ( \1227 , \1226 );
not \U$885 ( \1228 , \386 );
and \U$886 ( \1229 , \1227 , \1228 );
and \U$887 ( \1230 , \1226 , \386 );
nor \U$888 ( \1231 , \1229 , \1230 );
and \U$889 ( \1232 , \354 , RI986e620_21);
and \U$890 ( \1233 , RI986f7f0_59, \352 );
nor \U$891 ( \1234 , \1232 , \1233 );
not \U$892 ( \1235 , \1234 );
not \U$893 ( \1236 , \361 );
and \U$894 ( \1237 , \1235 , \1236 );
and \U$895 ( \1238 , \1234 , \345 );
nor \U$896 ( \1239 , \1237 , \1238 );
or \U$897 ( \1240 , \1231 , \1239 );
not \U$898 ( \1241 , \1239 );
not \U$899 ( \1242 , \1231 );
or \U$900 ( \1243 , \1241 , \1242 );
not \U$901 ( \1244 , \365 );
and \U$902 ( \1245 , \376 , RI986f8e0_61);
and \U$903 ( \1246 , RI986f430_51, \374 );
nor \U$904 ( \1247 , \1245 , \1246 );
not \U$905 ( \1248 , \1247 );
or \U$906 ( \1249 , \1244 , \1248 );
or \U$907 ( \1250 , \1247 , \367 );
nand \U$908 ( \1251 , \1249 , \1250 );
nand \U$909 ( \1252 , \1243 , \1251 );
nand \U$910 ( \1253 , \1240 , \1252 );
not \U$911 ( \1254 , \1253 );
and \U$912 ( \1255 , \776 , RI986dea0_5);
and \U$913 ( \1256 , RI986ddb0_3, \774 );
nor \U$914 ( \1257 , \1255 , \1256 );
and \U$915 ( \1258 , \1257 , \474 );
not \U$916 ( \1259 , \1257 );
and \U$917 ( \1260 , \1259 , \451 );
nor \U$918 ( \1261 , \1258 , \1260 );
and \U$919 ( \1262 , \438 , RI986f610_55);
and \U$920 ( \1263 , RI986df90_7, \436 );
nor \U$921 ( \1264 , \1262 , \1263 );
and \U$922 ( \1265 , \1264 , \444 );
not \U$923 ( \1266 , \1264 );
and \U$924 ( \1267 , \1266 , \443 );
nor \U$925 ( \1268 , \1265 , \1267 );
xor \U$926 ( \1269 , \1261 , \1268 );
not \U$927 ( \1270 , \454 );
and \U$928 ( \1271 , \465 , RI986f340_49);
and \U$929 ( \1272 , RI986f520_53, \463 );
nor \U$930 ( \1273 , \1271 , \1272 );
not \U$931 ( \1274 , \1273 );
or \U$932 ( \1275 , \1270 , \1274 );
or \U$933 ( \1276 , \1273 , \456 );
nand \U$934 ( \1277 , \1275 , \1276 );
and \U$935 ( \1278 , \1269 , \1277 );
and \U$936 ( \1279 , \1261 , \1268 );
nor \U$937 ( \1280 , \1278 , \1279 );
not \U$938 ( \1281 , \1280 );
or \U$939 ( \1282 , \1254 , \1281 );
or \U$940 ( \1283 , \1280 , \1253 );
nand \U$941 ( \1284 , \1282 , \1283 );
not \U$942 ( \1285 , \1284 );
and \U$943 ( \1286 , RI9871c08_136, RI98720b8_146);
not \U$944 ( \1287 , RI98720b8_146);
nor \U$945 ( \1288 , \1287 , RI98718c0_129);
not \U$946 ( \1289 , RI98718c0_129);
nor \U$947 ( \1290 , \1289 , RI98720b8_146);
or \U$948 ( \1291 , \1288 , \1290 );
nor \U$949 ( \1292 , RI9871c08_136, RI98720b8_146);
nor \U$950 ( \1293 , \1286 , \1291 , \1292 );
and \U$951 ( \1294 , \1293 , RI986dcc0_1);
and \U$952 ( \1295 , RI986e170_11, \1291 );
nor \U$953 ( \1296 , \1294 , \1295 );
not \U$954 ( \1297 , \1296 );
not \U$955 ( \1298 , \1128 );
and \U$956 ( \1299 , \1297 , \1298 );
not \U$957 ( \1300 , \1128 );
not \U$958 ( \1301 , \1300 );
and \U$959 ( \1302 , \1296 , \1301 );
nor \U$960 ( \1303 , \1299 , \1302 );
and \U$961 ( \1304 , RI98719b0_131, RI9871a28_132);
not \U$962 ( \1305 , RI9871a28_132);
nor \U$963 ( \1306 , \1305 , RI9871aa0_133);
not \U$964 ( \1307 , RI9871aa0_133);
nor \U$965 ( \1308 , \1307 , RI9871a28_132);
or \U$966 ( \1309 , \1306 , \1308 );
nor \U$967 ( \1310 , RI98719b0_131, RI9871a28_132);
nor \U$968 ( \1311 , \1304 , \1309 , \1310 );
nand \U$969 ( \1312 , RI986e350_15, \1311 );
and \U$970 ( \1313 , RI9871a28_132, RI9871aa0_133);
not \U$971 ( \1314 , RI98719b0_131);
nor \U$972 ( \1315 , \1313 , \1314 );
and \U$973 ( \1316 , \1312 , \1315 );
not \U$974 ( \1317 , \1312 );
buf \U$975 ( \1318 , \1315 );
not \U$976 ( \1319 , \1318 );
and \U$977 ( \1320 , \1317 , \1319 );
nor \U$978 ( \1321 , \1316 , \1320 );
xor \U$979 ( \1322 , \1303 , \1321 );
and \U$980 ( \1323 , RI98718c0_129, RI9871938_130);
and \U$981 ( \1324 , RI9871938_130, \1314 );
not \U$982 ( \1325 , RI9871938_130);
and \U$983 ( \1326 , \1325 , RI98719b0_131);
or \U$984 ( \1327 , \1324 , \1326 );
nor \U$985 ( \1328 , RI98718c0_129, RI9871938_130);
nor \U$986 ( \1329 , \1323 , \1327 , \1328 );
and \U$987 ( \1330 , \1329 , RI986e080_9);
and \U$988 ( \1331 , RI986e260_13, \1327 );
nor \U$989 ( \1332 , \1330 , \1331 );
not \U$990 ( \1333 , RI98719b0_131);
not \U$991 ( \1334 , RI9871938_130);
or \U$992 ( \1335 , \1333 , \1334 );
nand \U$993 ( \1336 , \1335 , RI98718c0_129);
not \U$994 ( \1337 , \1336 );
and \U$995 ( \1338 , \1332 , \1337 );
not \U$996 ( \1339 , \1332 );
and \U$997 ( \1340 , \1339 , \1336 );
nor \U$998 ( \1341 , \1338 , \1340 );
and \U$999 ( \1342 , \1322 , \1341 );
and \U$1000 ( \1343 , \1303 , \1321 );
or \U$1001 ( \1344 , \1342 , \1343 );
not \U$1002 ( \1345 , \1344 );
and \U$1003 ( \1346 , \1285 , \1345 );
and \U$1004 ( \1347 , \1284 , \1344 );
nor \U$1005 ( \1348 , \1346 , \1347 );
xor \U$1006 ( \1349 , \1223 , \1348 );
not \U$1007 ( \1350 , \1315 );
and \U$1008 ( \1351 , \1329 , RI986e260_13);
and \U$1009 ( \1352 , RI986e350_15, \1327 );
nor \U$1010 ( \1353 , \1351 , \1352 );
and \U$1011 ( \1354 , \1353 , \1336 );
not \U$1012 ( \1355 , \1353 );
and \U$1013 ( \1356 , \1355 , \1337 );
nor \U$1014 ( \1357 , \1354 , \1356 );
not \U$1015 ( \1358 , \1357 );
or \U$1016 ( \1359 , \1350 , \1358 );
or \U$1017 ( \1360 , \1357 , \1318 );
nand \U$1018 ( \1361 , \1359 , \1360 );
not \U$1019 ( \1362 , \1361 );
and \U$1020 ( \1363 , \1293 , RI986e170_11);
and \U$1021 ( \1364 , RI986e080_9, \1291 );
nor \U$1022 ( \1365 , \1363 , \1364 );
not \U$1023 ( \1366 , \1365 );
not \U$1024 ( \1367 , \1128 );
and \U$1025 ( \1368 , \1366 , \1367 );
and \U$1026 ( \1369 , \1365 , \1301 );
nor \U$1027 ( \1370 , \1368 , \1369 );
not \U$1028 ( \1371 , \1370 );
and \U$1029 ( \1372 , \1362 , \1371 );
and \U$1030 ( \1373 , \1361 , \1370 );
nor \U$1031 ( \1374 , \1372 , \1373 );
and \U$1032 ( \1375 , \438 , RI986df90_7);
and \U$1033 ( \1376 , RI986dea0_5, \436 );
nor \U$1034 ( \1377 , \1375 , \1376 );
and \U$1035 ( \1378 , \1377 , \443 );
not \U$1036 ( \1379 , \1377 );
and \U$1037 ( \1380 , \1379 , \444 );
nor \U$1038 ( \1381 , \1378 , \1380 );
not \U$1039 ( \1382 , \1381 );
and \U$1040 ( \1383 , \776 , RI986ddb0_3);
and \U$1041 ( \1384 , RI986dcc0_1, \774 );
nor \U$1042 ( \1385 , \1383 , \1384 );
and \U$1043 ( \1386 , \1385 , \474 );
not \U$1044 ( \1387 , \1385 );
and \U$1045 ( \1388 , \1387 , \451 );
nor \U$1046 ( \1389 , \1386 , \1388 );
not \U$1047 ( \1390 , \1389 );
or \U$1048 ( \1391 , \1382 , \1390 );
or \U$1049 ( \1392 , \1381 , \1389 );
nand \U$1050 ( \1393 , \1391 , \1392 );
not \U$1051 ( \1394 , \1393 );
and \U$1052 ( \1395 , \465 , RI986f520_53);
and \U$1053 ( \1396 , RI986f610_55, \463 );
nor \U$1054 ( \1397 , \1395 , \1396 );
not \U$1055 ( \1398 , \1397 );
not \U$1056 ( \1399 , \454 );
and \U$1057 ( \1400 , \1398 , \1399 );
and \U$1058 ( \1401 , \1397 , \456 );
nor \U$1059 ( \1402 , \1400 , \1401 );
not \U$1060 ( \1403 , \1402 );
and \U$1061 ( \1404 , \1394 , \1403 );
and \U$1062 ( \1405 , \1393 , \1402 );
nor \U$1063 ( \1406 , \1404 , \1405 );
xor \U$1064 ( \1407 , \1374 , \1406 );
and \U$1065 ( \1408 , \395 , RI986f9d0_63);
and \U$1066 ( \1409 , RI986f8e0_61, \393 );
nor \U$1067 ( \1410 , \1408 , \1409 );
not \U$1068 ( \1411 , \1410 );
not \U$1069 ( \1412 , \487 );
and \U$1070 ( \1413 , \1411 , \1412 );
and \U$1071 ( \1414 , \1410 , \487 );
nor \U$1072 ( \1415 , \1413 , \1414 );
not \U$1073 ( \1416 , \1415 );
not \U$1074 ( \1417 , \365 );
and \U$1075 ( \1418 , \376 , RI986f430_51);
and \U$1076 ( \1419 , RI986f340_49, \374 );
nor \U$1077 ( \1420 , \1418 , \1419 );
not \U$1078 ( \1421 , \1420 );
or \U$1079 ( \1422 , \1417 , \1421 );
or \U$1080 ( \1423 , \1420 , \365 );
nand \U$1081 ( \1424 , \1422 , \1423 );
not \U$1082 ( \1425 , \1424 );
or \U$1083 ( \1426 , \1416 , \1425 );
or \U$1084 ( \1427 , \1415 , \1424 );
nand \U$1085 ( \1428 , \1426 , \1427 );
not \U$1086 ( \1429 , \1428 );
and \U$1087 ( \1430 , \354 , RI986f7f0_59);
and \U$1088 ( \1431 , RI986f700_57, \352 );
nor \U$1089 ( \1432 , \1430 , \1431 );
not \U$1090 ( \1433 , \1432 );
not \U$1091 ( \1434 , \361 );
and \U$1092 ( \1435 , \1433 , \1434 );
and \U$1093 ( \1436 , \1432 , \361 );
nor \U$1094 ( \1437 , \1435 , \1436 );
not \U$1095 ( \1438 , \1437 );
and \U$1096 ( \1439 , \1429 , \1438 );
and \U$1097 ( \1440 , \1428 , \1437 );
nor \U$1098 ( \1441 , \1439 , \1440 );
xor \U$1099 ( \1442 , \1407 , \1441 );
and \U$1100 ( \1443 , \1349 , \1442 );
and \U$1101 ( \1444 , \1223 , \1348 );
nor \U$1102 ( \1445 , \1443 , \1444 );
xor \U$1103 ( \1446 , \1261 , \1268 );
xor \U$1104 ( \1447 , \1446 , \1277 );
not \U$1105 ( \1448 , \1447 );
xor \U$1106 ( \1449 , \1303 , \1321 );
xor \U$1107 ( \1450 , \1449 , \1341 );
nor \U$1108 ( \1451 , \1448 , \1450 );
not \U$1109 ( \1452 , \1451 );
and \U$1110 ( \1453 , \1311 , RI986e260_13);
and \U$1111 ( \1454 , RI986e350_15, \1309 );
nor \U$1112 ( \1455 , \1453 , \1454 );
and \U$1113 ( \1456 , \1455 , \1315 );
not \U$1114 ( \1457 , \1455 );
not \U$1115 ( \1458 , \1315 );
and \U$1116 ( \1459 , \1457 , \1458 );
nor \U$1117 ( \1460 , \1456 , \1459 );
nand \U$1118 ( \1461 , RI9872310_151, RI9872298_150);
and \U$1119 ( \1462 , \1461 , RI9871aa0_133);
xor \U$1120 ( \1463 , \1460 , \1462 );
and \U$1121 ( \1464 , \1329 , RI986e170_11);
and \U$1122 ( \1465 , RI986e080_9, \1327 );
nor \U$1123 ( \1466 , \1464 , \1465 );
and \U$1124 ( \1467 , \1466 , \1337 );
not \U$1125 ( \1468 , \1466 );
and \U$1126 ( \1469 , \1468 , \1336 );
nor \U$1127 ( \1470 , \1467 , \1469 );
and \U$1128 ( \1471 , \1463 , \1470 );
and \U$1129 ( \1472 , \1460 , \1462 );
or \U$1130 ( \1473 , \1471 , \1472 );
and \U$1131 ( \1474 , \376 , RI986f9d0_63);
and \U$1132 ( \1475 , RI986f8e0_61, \374 );
nor \U$1133 ( \1476 , \1474 , \1475 );
not \U$1134 ( \1477 , \1476 );
not \U$1135 ( \1478 , \365 );
and \U$1136 ( \1479 , \1477 , \1478 );
and \U$1137 ( \1480 , \1476 , \367 );
nor \U$1138 ( \1481 , \1479 , \1480 );
and \U$1139 ( \1482 , \465 , RI986f430_51);
and \U$1140 ( \1483 , RI986f340_49, \463 );
nor \U$1141 ( \1484 , \1482 , \1483 );
not \U$1142 ( \1485 , \1484 );
not \U$1143 ( \1486 , \456 );
and \U$1144 ( \1487 , \1485 , \1486 );
and \U$1145 ( \1488 , \1484 , \456 );
nor \U$1146 ( \1489 , \1487 , \1488 );
xor \U$1147 ( \1490 , \1481 , \1489 );
and \U$1148 ( \1491 , \395 , RI986f7f0_59);
and \U$1149 ( \1492 , RI986f700_57, \393 );
nor \U$1150 ( \1493 , \1491 , \1492 );
not \U$1151 ( \1494 , \1493 );
not \U$1152 ( \1495 , \487 );
and \U$1153 ( \1496 , \1494 , \1495 );
and \U$1154 ( \1497 , \1493 , \386 );
nor \U$1155 ( \1498 , \1496 , \1497 );
and \U$1156 ( \1499 , \1490 , \1498 );
and \U$1157 ( \1500 , \1481 , \1489 );
or \U$1158 ( \1501 , \1499 , \1500 );
xor \U$1159 ( \1502 , \1473 , \1501 );
and \U$1160 ( \1503 , \776 , RI986df90_7);
and \U$1161 ( \1504 , RI986dea0_5, \774 );
nor \U$1162 ( \1505 , \1503 , \1504 );
and \U$1163 ( \1506 , \1505 , \451 );
not \U$1164 ( \1507 , \1505 );
and \U$1165 ( \1508 , \1507 , \474 );
nor \U$1166 ( \1509 , \1506 , \1508 );
not \U$1167 ( \1510 , \1509 );
and \U$1168 ( \1511 , \438 , RI986f520_53);
and \U$1169 ( \1512 , RI986f610_55, \436 );
nor \U$1170 ( \1513 , \1511 , \1512 );
and \U$1171 ( \1514 , \1513 , \443 );
not \U$1172 ( \1515 , \1513 );
and \U$1173 ( \1516 , \1515 , \444 );
nor \U$1174 ( \1517 , \1514 , \1516 );
not \U$1175 ( \1518 , \1517 );
and \U$1176 ( \1519 , \1510 , \1518 );
and \U$1177 ( \1520 , \1517 , \1509 );
and \U$1178 ( \1521 , \1293 , RI986ddb0_3);
and \U$1179 ( \1522 , RI986dcc0_1, \1291 );
nor \U$1180 ( \1523 , \1521 , \1522 );
not \U$1181 ( \1524 , \1523 );
not \U$1182 ( \1525 , \1301 );
and \U$1183 ( \1526 , \1524 , \1525 );
and \U$1184 ( \1527 , \1523 , \1128 );
nor \U$1185 ( \1528 , \1526 , \1527 );
nor \U$1186 ( \1529 , \1520 , \1528 );
nor \U$1187 ( \1530 , \1519 , \1529 );
and \U$1188 ( \1531 , \1502 , \1530 );
and \U$1189 ( \1532 , \1473 , \1501 );
nor \U$1190 ( \1533 , \1531 , \1532 );
not \U$1191 ( \1534 , \1533 );
or \U$1192 ( \1535 , \1452 , \1534 );
or \U$1193 ( \1536 , \1533 , \1451 );
not \U$1194 ( \1537 , \1231 );
not \U$1195 ( \1538 , \1251 );
or \U$1196 ( \1539 , \1537 , \1538 );
or \U$1197 ( \1540 , \1231 , \1251 );
nand \U$1198 ( \1541 , \1539 , \1540 );
not \U$1199 ( \1542 , \1541 );
not \U$1200 ( \1543 , \1239 );
and \U$1201 ( \1544 , \1542 , \1543 );
and \U$1202 ( \1545 , \1541 , \1239 );
nor \U$1203 ( \1546 , \1544 , \1545 );
and \U$1204 ( \1547 , \416 , RI986e530_19);
and \U$1205 ( \1548 , RI986e440_17, \414 );
nor \U$1206 ( \1549 , \1547 , \1548 );
and \U$1207 ( \1550 , \1549 , \421 );
not \U$1208 ( \1551 , \1549 );
and \U$1209 ( \1552 , \1551 , \422 );
nor \U$1210 ( \1553 , \1550 , \1552 );
nand \U$1211 ( \1554 , RI986f160_45, RI9871fc8_144);
xor \U$1212 ( \1555 , \1553 , \1554 );
and \U$1213 ( \1556 , \354 , RI986e710_23);
and \U$1214 ( \1557 , RI986e620_21, \352 );
nor \U$1215 ( \1558 , \1556 , \1557 );
not \U$1216 ( \1559 , \1558 );
not \U$1217 ( \1560 , \361 );
and \U$1218 ( \1561 , \1559 , \1560 );
and \U$1219 ( \1562 , \1558 , \345 );
nor \U$1220 ( \1563 , \1561 , \1562 );
and \U$1221 ( \1564 , \1555 , \1563 );
and \U$1222 ( \1565 , \1553 , \1554 );
or \U$1223 ( \1566 , \1564 , \1565 );
or \U$1224 ( \1567 , \1546 , \1566 );
not \U$1225 ( \1568 , \1566 );
not \U$1226 ( \1569 , \1546 );
or \U$1227 ( \1570 , \1568 , \1569 );
or \U$1228 ( \1571 , \1212 , \1205 );
nand \U$1229 ( \1572 , \1571 , \1213 );
nand \U$1230 ( \1573 , \1570 , \1572 );
nand \U$1231 ( \1574 , \1567 , \1573 );
nand \U$1232 ( \1575 , \1536 , \1574 );
nand \U$1233 ( \1576 , \1535 , \1575 );
xor \U$1234 ( \1577 , \1445 , \1576 );
not \U$1235 ( \1578 , \361 );
and \U$1236 ( \1579 , \354 , RI986f700_57);
and \U$1237 ( \1580 , RI986f9d0_63, \352 );
nor \U$1238 ( \1581 , \1579 , \1580 );
not \U$1239 ( \1582 , \1581 );
or \U$1240 ( \1583 , \1578 , \1582 );
or \U$1241 ( \1584 , \1581 , \361 );
nand \U$1242 ( \1585 , \1583 , \1584 );
not \U$1243 ( \1586 , \1585 );
and \U$1244 ( \1587 , \395 , RI986f8e0_61);
and \U$1245 ( \1588 , RI986f430_51, \393 );
nor \U$1246 ( \1589 , \1587 , \1588 );
not \U$1247 ( \1590 , \1589 );
not \U$1248 ( \1591 , \386 );
and \U$1249 ( \1592 , \1590 , \1591 );
and \U$1250 ( \1593 , \1589 , \386 );
nor \U$1251 ( \1594 , \1592 , \1593 );
not \U$1252 ( \1595 , \1594 );
or \U$1253 ( \1596 , \1586 , \1595 );
or \U$1254 ( \1597 , \1594 , \1585 );
nand \U$1255 ( \1598 , \1596 , \1597 );
not \U$1256 ( \1599 , \1598 );
and \U$1257 ( \1600 , \416 , RI986e620_21);
and \U$1258 ( \1601 , RI986f7f0_59, \414 );
nor \U$1259 ( \1602 , \1600 , \1601 );
and \U$1260 ( \1603 , \1602 , \421 );
not \U$1261 ( \1604 , \1602 );
and \U$1262 ( \1605 , \1604 , \422 );
nor \U$1263 ( \1606 , \1603 , \1605 );
not \U$1264 ( \1607 , \1606 );
and \U$1265 ( \1608 , \1599 , \1607 );
and \U$1266 ( \1609 , \1598 , \1606 );
nor \U$1267 ( \1610 , \1608 , \1609 );
nand \U$1268 ( \1611 , RI986e710_23, RI9871fc8_144);
or \U$1269 ( \1612 , \1610 , \1611 );
nand \U$1270 ( \1613 , \1611 , \1610 );
nand \U$1271 ( \1614 , \1612 , \1613 );
not \U$1272 ( \1615 , \454 );
and \U$1273 ( \1616 , \465 , RI986f610_55);
and \U$1274 ( \1617 , RI986df90_7, \463 );
nor \U$1275 ( \1618 , \1616 , \1617 );
not \U$1276 ( \1619 , \1618 );
or \U$1277 ( \1620 , \1615 , \1619 );
or \U$1278 ( \1621 , \1618 , \456 );
nand \U$1279 ( \1622 , \1620 , \1621 );
and \U$1280 ( \1623 , \438 , RI986dea0_5);
and \U$1281 ( \1624 , RI986ddb0_3, \436 );
nor \U$1282 ( \1625 , \1623 , \1624 );
and \U$1283 ( \1626 , \1625 , \444 );
not \U$1284 ( \1627 , \1625 );
and \U$1285 ( \1628 , \1627 , \443 );
nor \U$1286 ( \1629 , \1626 , \1628 );
xor \U$1287 ( \1630 , \1622 , \1629 );
not \U$1288 ( \1631 , \365 );
and \U$1289 ( \1632 , \376 , RI986f340_49);
and \U$1290 ( \1633 , RI986f520_53, \374 );
nor \U$1291 ( \1634 , \1632 , \1633 );
not \U$1292 ( \1635 , \1634 );
or \U$1293 ( \1636 , \1631 , \1635 );
or \U$1294 ( \1637 , \1634 , \365 );
nand \U$1295 ( \1638 , \1636 , \1637 );
xor \U$1296 ( \1639 , \1630 , \1638 );
and \U$1297 ( \1640 , \776 , RI986dcc0_1);
and \U$1298 ( \1641 , RI986e170_11, \774 );
nor \U$1299 ( \1642 , \1640 , \1641 );
and \U$1300 ( \1643 , \1642 , \474 );
not \U$1301 ( \1644 , \1642 );
and \U$1302 ( \1645 , \1644 , \451 );
nor \U$1303 ( \1646 , \1643 , \1645 );
nand \U$1304 ( \1647 , RI986e350_15, \1329 );
and \U$1305 ( \1648 , \1647 , \1336 );
not \U$1306 ( \1649 , \1647 );
and \U$1307 ( \1650 , \1649 , \1337 );
nor \U$1308 ( \1651 , \1648 , \1650 );
xor \U$1309 ( \1652 , \1646 , \1651 );
not \U$1310 ( \1653 , \1128 );
and \U$1311 ( \1654 , \1293 , RI986e080_9);
and \U$1312 ( \1655 , RI986e260_13, \1291 );
nor \U$1313 ( \1656 , \1654 , \1655 );
not \U$1314 ( \1657 , \1656 );
or \U$1315 ( \1658 , \1653 , \1657 );
or \U$1316 ( \1659 , \1656 , \1301 );
nand \U$1317 ( \1660 , \1658 , \1659 );
xor \U$1318 ( \1661 , \1652 , \1660 );
xor \U$1319 ( \1662 , \1639 , \1661 );
xor \U$1320 ( \1663 , \1614 , \1662 );
or \U$1321 ( \1664 , \1415 , \1437 );
not \U$1322 ( \1665 , \1437 );
not \U$1323 ( \1666 , \1415 );
or \U$1324 ( \1667 , \1665 , \1666 );
nand \U$1325 ( \1668 , \1667 , \1424 );
nand \U$1326 ( \1669 , \1664 , \1668 );
or \U$1327 ( \1670 , \1370 , \1318 );
not \U$1328 ( \1671 , \1318 );
not \U$1329 ( \1672 , \1370 );
or \U$1330 ( \1673 , \1671 , \1672 );
nand \U$1331 ( \1674 , \1673 , \1357 );
nand \U$1332 ( \1675 , \1670 , \1674 );
xor \U$1333 ( \1676 , \1669 , \1675 );
or \U$1334 ( \1677 , \1381 , \1402 );
not \U$1335 ( \1678 , \1402 );
not \U$1336 ( \1679 , \1381 );
or \U$1337 ( \1680 , \1678 , \1679 );
nand \U$1338 ( \1681 , \1680 , \1389 );
nand \U$1339 ( \1682 , \1677 , \1681 );
xor \U$1340 ( \1683 , \1676 , \1682 );
xor \U$1341 ( \1684 , \1663 , \1683 );
and \U$1342 ( \1685 , \1577 , \1684 );
and \U$1343 ( \1686 , \1445 , \1576 );
or \U$1344 ( \1687 , \1685 , \1686 );
and \U$1345 ( \1688 , \1639 , \1661 );
xor \U$1346 ( \1689 , \1688 , \1613 );
xor \U$1347 ( \1690 , \1669 , \1675 );
and \U$1348 ( \1691 , \1690 , \1682 );
and \U$1349 ( \1692 , \1669 , \1675 );
or \U$1350 ( \1693 , \1691 , \1692 );
xor \U$1351 ( \1694 , \1689 , \1693 );
xor \U$1352 ( \1695 , \1687 , \1694 );
xor \U$1353 ( \1696 , \1614 , \1662 );
and \U$1354 ( \1697 , \1696 , \1683 );
and \U$1355 ( \1698 , \1614 , \1662 );
or \U$1356 ( \1699 , \1697 , \1698 );
not \U$1357 ( \1700 , \1253 );
or \U$1358 ( \1701 , \1344 , \1700 );
and \U$1359 ( \1702 , \1700 , \1344 );
nor \U$1360 ( \1703 , \1702 , \1280 );
not \U$1361 ( \1704 , \1703 );
nand \U$1362 ( \1705 , \1701 , \1704 );
or \U$1363 ( \1706 , \1203 , \1219 );
not \U$1364 ( \1707 , \1219 );
not \U$1365 ( \1708 , \1203 );
or \U$1366 ( \1709 , \1707 , \1708 );
nand \U$1367 ( \1710 , \1709 , \1213 );
nand \U$1368 ( \1711 , \1706 , \1710 );
xor \U$1369 ( \1712 , \1705 , \1711 );
xor \U$1370 ( \1713 , \1374 , \1406 );
and \U$1371 ( \1714 , \1713 , \1441 );
and \U$1372 ( \1715 , \1374 , \1406 );
nor \U$1373 ( \1716 , \1714 , \1715 );
and \U$1374 ( \1717 , \1712 , \1716 );
and \U$1375 ( \1718 , \1705 , \1711 );
or \U$1376 ( \1719 , \1717 , \1718 );
xor \U$1377 ( \1720 , \1699 , \1719 );
xor \U$1378 ( \1721 , \1622 , \1629 );
and \U$1379 ( \1722 , \1721 , \1638 );
and \U$1380 ( \1723 , \1622 , \1629 );
or \U$1381 ( \1724 , \1722 , \1723 );
or \U$1382 ( \1725 , \1594 , \1606 );
not \U$1383 ( \1726 , \1606 );
not \U$1384 ( \1727 , \1594 );
or \U$1385 ( \1728 , \1726 , \1727 );
nand \U$1386 ( \1729 , \1728 , \1585 );
nand \U$1387 ( \1730 , \1725 , \1729 );
xor \U$1388 ( \1731 , \1724 , \1730 );
xor \U$1389 ( \1732 , \1646 , \1651 );
and \U$1390 ( \1733 , \1732 , \1660 );
and \U$1391 ( \1734 , \1646 , \1651 );
or \U$1392 ( \1735 , \1733 , \1734 );
xor \U$1393 ( \1736 , \1731 , \1735 );
and \U$1394 ( \1737 , \776 , RI986e170_11);
and \U$1395 ( \1738 , RI986e080_9, \774 );
nor \U$1396 ( \1739 , \1737 , \1738 );
and \U$1397 ( \1740 , \1739 , \474 );
not \U$1398 ( \1741 , \1739 );
and \U$1399 ( \1742 , \1741 , \451 );
nor \U$1400 ( \1743 , \1740 , \1742 );
not \U$1401 ( \1744 , \1743 );
not \U$1402 ( \1745 , \1301 );
and \U$1403 ( \1746 , \1293 , RI986e260_13);
and \U$1404 ( \1747 , RI986e350_15, \1291 );
nor \U$1405 ( \1748 , \1746 , \1747 );
not \U$1406 ( \1749 , \1748 );
or \U$1407 ( \1750 , \1745 , \1749 );
or \U$1408 ( \1751 , \1748 , \1128 );
nand \U$1409 ( \1752 , \1750 , \1751 );
and \U$1410 ( \1753 , \1752 , \1337 );
nor \U$1411 ( \1754 , \1752 , \1337 );
nor \U$1412 ( \1755 , \1753 , \1754 );
not \U$1413 ( \1756 , \1755 );
or \U$1414 ( \1757 , \1744 , \1756 );
or \U$1415 ( \1758 , \1755 , \1743 );
nand \U$1416 ( \1759 , \1757 , \1758 );
and \U$1417 ( \1760 , \438 , RI986ddb0_3);
and \U$1418 ( \1761 , RI986dcc0_1, \436 );
nor \U$1419 ( \1762 , \1760 , \1761 );
and \U$1420 ( \1763 , \1762 , \444 );
not \U$1421 ( \1764 , \1762 );
and \U$1422 ( \1765 , \1764 , \443 );
nor \U$1423 ( \1766 , \1763 , \1765 );
not \U$1424 ( \1767 , \456 );
and \U$1425 ( \1768 , \465 , RI986df90_7);
and \U$1426 ( \1769 , RI986dea0_5, \463 );
nor \U$1427 ( \1770 , \1768 , \1769 );
not \U$1428 ( \1771 , \1770 );
or \U$1429 ( \1772 , \1767 , \1771 );
or \U$1430 ( \1773 , \1770 , \456 );
nand \U$1431 ( \1774 , \1772 , \1773 );
xor \U$1432 ( \1775 , \1766 , \1774 );
not \U$1433 ( \1776 , \365 );
and \U$1434 ( \1777 , \376 , RI986f520_53);
and \U$1435 ( \1778 , RI986f610_55, \374 );
nor \U$1436 ( \1779 , \1777 , \1778 );
not \U$1437 ( \1780 , \1779 );
or \U$1438 ( \1781 , \1776 , \1780 );
or \U$1439 ( \1782 , \1779 , \365 );
nand \U$1440 ( \1783 , \1781 , \1782 );
xor \U$1441 ( \1784 , \1775 , \1783 );
not \U$1442 ( \1785 , RI986e620_21);
nor \U$1443 ( \1786 , \1785 , \407 );
xor \U$1444 ( \1787 , \1784 , \1786 );
and \U$1445 ( \1788 , \416 , RI986f7f0_59);
and \U$1446 ( \1789 , RI986f700_57, \414 );
nor \U$1447 ( \1790 , \1788 , \1789 );
and \U$1448 ( \1791 , \1790 , \421 );
not \U$1449 ( \1792 , \1790 );
and \U$1450 ( \1793 , \1792 , \422 );
nor \U$1451 ( \1794 , \1791 , \1793 );
not \U$1452 ( \1795 , \1794 );
and \U$1453 ( \1796 , \395 , RI986f430_51);
and \U$1454 ( \1797 , RI986f340_49, \393 );
nor \U$1455 ( \1798 , \1796 , \1797 );
not \U$1456 ( \1799 , \1798 );
not \U$1457 ( \1800 , \386 );
and \U$1458 ( \1801 , \1799 , \1800 );
and \U$1459 ( \1802 , \1798 , \386 );
nor \U$1460 ( \1803 , \1801 , \1802 );
and \U$1461 ( \1804 , \354 , RI986f9d0_63);
and \U$1462 ( \1805 , RI986f8e0_61, \352 );
nor \U$1463 ( \1806 , \1804 , \1805 );
not \U$1464 ( \1807 , \1806 );
not \U$1465 ( \1808 , \361 );
and \U$1466 ( \1809 , \1807 , \1808 );
and \U$1467 ( \1810 , \1806 , \361 );
nor \U$1468 ( \1811 , \1809 , \1810 );
xor \U$1469 ( \1812 , \1803 , \1811 );
not \U$1470 ( \1813 , \1812 );
or \U$1471 ( \1814 , \1795 , \1813 );
or \U$1472 ( \1815 , \1812 , \1794 );
nand \U$1473 ( \1816 , \1814 , \1815 );
xor \U$1474 ( \1817 , \1787 , \1816 );
xor \U$1475 ( \1818 , \1759 , \1817 );
xor \U$1476 ( \1819 , \1736 , \1818 );
xor \U$1477 ( \1820 , \1720 , \1819 );
and \U$1478 ( \1821 , \1695 , \1820 );
and \U$1479 ( \1822 , \1687 , \1694 );
or \U$1480 ( \1823 , \1821 , \1822 );
not \U$1481 ( \1824 , \1823 );
xor \U$1482 ( \1825 , \1699 , \1719 );
and \U$1483 ( \1826 , \1825 , \1819 );
and \U$1484 ( \1827 , \1699 , \1719 );
or \U$1485 ( \1828 , \1826 , \1827 );
xor \U$1486 ( \1829 , \1688 , \1613 );
and \U$1487 ( \1830 , \1829 , \1693 );
and \U$1488 ( \1831 , \1688 , \1613 );
or \U$1489 ( \1832 , \1830 , \1831 );
and \U$1490 ( \1833 , \354 , RI986f8e0_61);
and \U$1491 ( \1834 , RI986f430_51, \352 );
nor \U$1492 ( \1835 , \1833 , \1834 );
not \U$1493 ( \1836 , \1835 );
not \U$1494 ( \1837 , \345 );
and \U$1495 ( \1838 , \1836 , \1837 );
and \U$1496 ( \1839 , \1835 , \345 );
nor \U$1497 ( \1840 , \1838 , \1839 );
nand \U$1498 ( \1841 , RI986f7f0_59, RI9871fc8_144);
xor \U$1499 ( \1842 , \1840 , \1841 );
and \U$1500 ( \1843 , \416 , RI986f700_57);
and \U$1501 ( \1844 , RI986f9d0_63, \414 );
nor \U$1502 ( \1845 , \1843 , \1844 );
and \U$1503 ( \1846 , \1845 , \421 );
not \U$1504 ( \1847 , \1845 );
and \U$1505 ( \1848 , \1847 , \422 );
nor \U$1506 ( \1849 , \1846 , \1848 );
xor \U$1507 ( \1850 , \1842 , \1849 );
and \U$1508 ( \1851 , \376 , RI986f610_55);
and \U$1509 ( \1852 , RI986df90_7, \374 );
nor \U$1510 ( \1853 , \1851 , \1852 );
not \U$1511 ( \1854 , \1853 );
not \U$1512 ( \1855 , \365 );
and \U$1513 ( \1856 , \1854 , \1855 );
and \U$1514 ( \1857 , \1853 , \365 );
nor \U$1515 ( \1858 , \1856 , \1857 );
and \U$1516 ( \1859 , \465 , RI986dea0_5);
and \U$1517 ( \1860 , RI986ddb0_3, \463 );
nor \U$1518 ( \1861 , \1859 , \1860 );
not \U$1519 ( \1862 , \1861 );
not \U$1520 ( \1863 , \454 );
and \U$1521 ( \1864 , \1862 , \1863 );
and \U$1522 ( \1865 , \1861 , \456 );
nor \U$1523 ( \1866 , \1864 , \1865 );
xor \U$1524 ( \1867 , \1858 , \1866 );
and \U$1525 ( \1868 , \395 , RI986f340_49);
and \U$1526 ( \1869 , RI986f520_53, \393 );
nor \U$1527 ( \1870 , \1868 , \1869 );
not \U$1528 ( \1871 , \1870 );
not \U$1529 ( \1872 , \487 );
and \U$1530 ( \1873 , \1871 , \1872 );
and \U$1531 ( \1874 , \1870 , \487 );
nor \U$1532 ( \1875 , \1873 , \1874 );
xor \U$1533 ( \1876 , \1867 , \1875 );
or \U$1534 ( \1877 , \1850 , \1876 );
nand \U$1535 ( \1878 , \1850 , \1876 );
nand \U$1536 ( \1879 , \1877 , \1878 );
xor \U$1537 ( \1880 , \1832 , \1879 );
xor \U$1538 ( \1881 , \1724 , \1730 );
xor \U$1539 ( \1882 , \1881 , \1735 );
and \U$1540 ( \1883 , \1759 , \1882 );
xor \U$1541 ( \1884 , \1724 , \1730 );
xor \U$1542 ( \1885 , \1884 , \1735 );
and \U$1543 ( \1886 , \1817 , \1885 );
and \U$1544 ( \1887 , \1759 , \1817 );
or \U$1545 ( \1888 , \1883 , \1886 , \1887 );
xor \U$1546 ( \1889 , \1880 , \1888 );
xnor \U$1547 ( \1890 , \1828 , \1889 );
not \U$1548 ( \1891 , \1890 );
not \U$1549 ( \1892 , \1803 );
not \U$1550 ( \1893 , \1794 );
and \U$1551 ( \1894 , \1892 , \1893 );
and \U$1552 ( \1895 , \1803 , \1794 );
nor \U$1553 ( \1896 , \1895 , \1811 );
nor \U$1554 ( \1897 , \1894 , \1896 );
not \U$1555 ( \1898 , \1752 );
nand \U$1556 ( \1899 , \1898 , \1337 );
and \U$1557 ( \1900 , \1899 , \1743 );
and \U$1558 ( \1901 , \1336 , \1752 );
nor \U$1559 ( \1902 , \1900 , \1901 );
xor \U$1560 ( \1903 , \1897 , \1902 );
xor \U$1561 ( \1904 , \1766 , \1774 );
and \U$1562 ( \1905 , \1904 , \1783 );
and \U$1563 ( \1906 , \1766 , \1774 );
nor \U$1564 ( \1907 , \1905 , \1906 );
xor \U$1565 ( \1908 , \1903 , \1907 );
not \U$1566 ( \1909 , \1908 );
and \U$1567 ( \1910 , \438 , RI986dcc0_1);
and \U$1568 ( \1911 , RI986e170_11, \436 );
nor \U$1569 ( \1912 , \1910 , \1911 );
and \U$1570 ( \1913 , \1912 , \443 );
not \U$1571 ( \1914 , \1912 );
and \U$1572 ( \1915 , \1914 , \444 );
nor \U$1573 ( \1916 , \1913 , \1915 );
not \U$1574 ( \1917 , \1916 );
nand \U$1575 ( \1918 , RI986e350_15, \1293 );
not \U$1576 ( \1919 , \1918 );
not \U$1577 ( \1920 , \1301 );
and \U$1578 ( \1921 , \1919 , \1920 );
and \U$1579 ( \1922 , \1918 , \1301 );
nor \U$1580 ( \1923 , \1921 , \1922 );
and \U$1581 ( \1924 , \776 , RI986e080_9);
and \U$1582 ( \1925 , RI986e260_13, \774 );
nor \U$1583 ( \1926 , \1924 , \1925 );
and \U$1584 ( \1927 , \1926 , \451 );
not \U$1585 ( \1928 , \1926 );
and \U$1586 ( \1929 , \1928 , \474 );
nor \U$1587 ( \1930 , \1927 , \1929 );
xor \U$1588 ( \1931 , \1923 , \1930 );
not \U$1589 ( \1932 , \1931 );
or \U$1590 ( \1933 , \1917 , \1932 );
or \U$1591 ( \1934 , \1931 , \1916 );
nand \U$1592 ( \1935 , \1933 , \1934 );
xor \U$1593 ( \1936 , \1724 , \1730 );
and \U$1594 ( \1937 , \1936 , \1735 );
and \U$1595 ( \1938 , \1724 , \1730 );
or \U$1596 ( \1939 , \1937 , \1938 );
not \U$1597 ( \1940 , \1939 );
xor \U$1598 ( \1941 , \1784 , \1786 );
and \U$1599 ( \1942 , \1941 , \1816 );
and \U$1600 ( \1943 , \1784 , \1786 );
nor \U$1601 ( \1944 , \1942 , \1943 );
not \U$1602 ( \1945 , \1944 );
or \U$1603 ( \1946 , \1940 , \1945 );
or \U$1604 ( \1947 , \1944 , \1939 );
nand \U$1605 ( \1948 , \1946 , \1947 );
xor \U$1606 ( \1949 , \1935 , \1948 );
not \U$1607 ( \1950 , \1949 );
or \U$1608 ( \1951 , \1909 , \1950 );
or \U$1609 ( \1952 , \1949 , \1908 );
nand \U$1610 ( \1953 , \1951 , \1952 );
not \U$1611 ( \1954 , \1953 );
and \U$1612 ( \1955 , \1891 , \1954 );
and \U$1613 ( \1956 , \1890 , \1953 );
nor \U$1614 ( \1957 , \1955 , \1956 );
nor \U$1615 ( \1958 , \1824 , \1957 );
not \U$1616 ( \1959 , \1908 );
nand \U$1617 ( \1960 , \1959 , \1949 );
not \U$1618 ( \1961 , \1960 );
xor \U$1619 ( \1962 , \1832 , \1879 );
and \U$1620 ( \1963 , \1962 , \1888 );
and \U$1621 ( \1964 , \1832 , \1879 );
or \U$1622 ( \1965 , \1963 , \1964 );
not \U$1623 ( \1966 , \1965 );
or \U$1624 ( \1967 , \1961 , \1966 );
or \U$1625 ( \1968 , \1965 , \1960 );
nand \U$1626 ( \1969 , \1967 , \1968 );
not \U$1627 ( \1970 , \1969 );
and \U$1628 ( \1971 , \1939 , \1935 );
not \U$1629 ( \1972 , \1939 );
not \U$1630 ( \1973 , \1935 );
and \U$1631 ( \1974 , \1972 , \1973 );
nor \U$1632 ( \1975 , \1974 , \1944 );
nor \U$1633 ( \1976 , \1971 , \1975 );
xor \U$1634 ( \1977 , \1858 , \1866 );
and \U$1635 ( \1978 , \1977 , \1875 );
and \U$1636 ( \1979 , \1858 , \1866 );
or \U$1637 ( \1980 , \1978 , \1979 );
xor \U$1638 ( \1981 , \1840 , \1841 );
and \U$1639 ( \1982 , \1981 , \1849 );
and \U$1640 ( \1983 , \1840 , \1841 );
or \U$1641 ( \1984 , \1982 , \1983 );
xor \U$1642 ( \1985 , \1980 , \1984 );
not \U$1643 ( \1986 , \1930 );
not \U$1644 ( \1987 , \1916 );
and \U$1645 ( \1988 , \1986 , \1987 );
and \U$1646 ( \1989 , \1916 , \1930 );
nor \U$1647 ( \1990 , \1989 , \1923 );
nor \U$1648 ( \1991 , \1988 , \1990 );
xor \U$1649 ( \1992 , \1985 , \1991 );
xor \U$1650 ( \1993 , \1976 , \1992 );
xor \U$1651 ( \1994 , \1897 , \1902 );
and \U$1652 ( \1995 , \1994 , \1907 );
and \U$1653 ( \1996 , \1897 , \1902 );
or \U$1654 ( \1997 , \1995 , \1996 );
not \U$1655 ( \1998 , \1878 );
xor \U$1656 ( \1999 , \1997 , \1998 );
xor \U$1657 ( \2000 , \1126 , \1128 );
xor \U$1658 ( \2001 , \2000 , \1136 );
xor \U$1659 ( \2002 , \1107 , \1108 );
xor \U$1660 ( \2003 , \2002 , \1116 );
xor \U$1661 ( \2004 , \1148 , \1156 );
xor \U$1662 ( \2005 , \2004 , \1165 );
xor \U$1663 ( \2006 , \2003 , \2005 );
xor \U$1664 ( \2007 , \2001 , \2006 );
xor \U$1665 ( \2008 , \1999 , \2007 );
xor \U$1666 ( \2009 , \1993 , \2008 );
not \U$1667 ( \2010 , \2009 );
and \U$1668 ( \2011 , \1970 , \2010 );
and \U$1669 ( \2012 , \1969 , \2009 );
nor \U$1670 ( \2013 , \2011 , \2012 );
not \U$1671 ( \2014 , \2013 );
not \U$1672 ( \2015 , \1953 );
not \U$1673 ( \2016 , \1889 );
or \U$1674 ( \2017 , \2015 , \2016 );
or \U$1675 ( \2018 , \1889 , \1953 );
nand \U$1676 ( \2019 , \2018 , \1828 );
nand \U$1677 ( \2020 , \2017 , \2019 );
not \U$1678 ( \2021 , \2020 );
or \U$1679 ( \2022 , \2014 , \2021 );
or \U$1680 ( \2023 , \2020 , \2013 );
nand \U$1681 ( \2024 , \2022 , \2023 );
and \U$1682 ( \2025 , \1958 , \2024 );
xor \U$1683 ( \2026 , \2024 , \1958 );
not \U$1684 ( \2027 , RI98726d0_159);
not \U$1685 ( \2028 , RI9872748_160);
or \U$1686 ( \2029 , \2027 , \2028 );
nand \U$1687 ( \2030 , \2029 , RI9872310_151);
not \U$1688 ( \2031 , \2030 );
not \U$1689 ( \2032 , \2031 );
not \U$1690 ( \2033 , \1462 );
not \U$1691 ( \2034 , \2033 );
not \U$1692 ( \2035 , \2034 );
and \U$1693 ( \2036 , RI9871aa0_133, RI9872298_150);
not \U$1694 ( \2037 , RI9872310_151);
and \U$1695 ( \2038 , \2037 , RI9872298_150);
nor \U$1696 ( \2039 , \2037 , RI9872298_150);
or \U$1697 ( \2040 , \2038 , \2039 );
nor \U$1698 ( \2041 , RI9871aa0_133, RI9872298_150);
nor \U$1699 ( \2042 , \2036 , \2040 , \2041 );
and \U$1700 ( \2043 , \2042 , RI986e260_13);
and \U$1701 ( \2044 , RI986e350_15, \2040 );
nor \U$1702 ( \2045 , \2043 , \2044 );
not \U$1703 ( \2046 , \2045 );
or \U$1704 ( \2047 , \2035 , \2046 );
or \U$1705 ( \2048 , \2045 , \2034 );
nand \U$1706 ( \2049 , \2047 , \2048 );
not \U$1707 ( \2050 , \2049 );
or \U$1708 ( \2051 , \2032 , \2050 );
or \U$1709 ( \2052 , \2049 , \2031 );
nand \U$1710 ( \2053 , \2051 , \2052 );
not \U$1711 ( \2054 , \2053 );
and \U$1712 ( \2055 , \1311 , RI986e170_11);
and \U$1713 ( \2056 , RI986e080_9, \1309 );
nor \U$1714 ( \2057 , \2055 , \2056 );
and \U$1715 ( \2058 , \2057 , \1315 );
not \U$1716 ( \2059 , \2057 );
and \U$1717 ( \2060 , \2059 , \1458 );
nor \U$1718 ( \2061 , \2058 , \2060 );
not \U$1719 ( \2062 , \2061 );
and \U$1720 ( \2063 , \2054 , \2062 );
and \U$1721 ( \2064 , \2053 , \2061 );
nor \U$1722 ( \2065 , \2063 , \2064 );
nand \U$1723 ( \2066 , RI986f070_43, RI9871fc8_144);
nand \U$1724 ( \2067 , RI986ef80_41, RI9871fc8_144);
xor \U$1725 ( \2068 , \2066 , \2067 );
and \U$1726 ( \2069 , \354 , RI986f160_45);
and \U$1727 ( \2070 , RI986e530_19, \352 );
nor \U$1728 ( \2071 , \2069 , \2070 );
not \U$1729 ( \2072 , \2071 );
not \U$1730 ( \2073 , \345 );
and \U$1731 ( \2074 , \2072 , \2073 );
and \U$1732 ( \2075 , \2071 , \345 );
nor \U$1733 ( \2076 , \2074 , \2075 );
not \U$1734 ( \2077 , \2076 );
and \U$1735 ( \2078 , \416 , RI986ef80_41);
and \U$1736 ( \2079 , RI986f250_47, \414 );
nor \U$1737 ( \2080 , \2078 , \2079 );
and \U$1738 ( \2081 , \2080 , \421 );
not \U$1739 ( \2082 , \2080 );
and \U$1740 ( \2083 , \2082 , \422 );
nor \U$1741 ( \2084 , \2081 , \2083 );
not \U$1742 ( \2085 , \2084 );
and \U$1743 ( \2086 , \2077 , \2085 );
and \U$1744 ( \2087 , \2084 , \2076 );
and \U$1745 ( \2088 , \395 , RI986e440_17);
and \U$1746 ( \2089 , RI986e710_23, \393 );
nor \U$1747 ( \2090 , \2088 , \2089 );
not \U$1748 ( \2091 , \2090 );
not \U$1749 ( \2092 , \487 );
and \U$1750 ( \2093 , \2091 , \2092 );
and \U$1751 ( \2094 , \2090 , \386 );
nor \U$1752 ( \2095 , \2093 , \2094 );
nor \U$1753 ( \2096 , \2087 , \2095 );
nor \U$1754 ( \2097 , \2086 , \2096 );
xor \U$1755 ( \2098 , \2068 , \2097 );
xor \U$1756 ( \2099 , \2065 , \2098 );
and \U$1757 ( \2100 , \465 , RI986f9d0_63);
and \U$1758 ( \2101 , RI986f8e0_61, \463 );
nor \U$1759 ( \2102 , \2100 , \2101 );
not \U$1760 ( \2103 , \2102 );
not \U$1761 ( \2104 , \456 );
and \U$1762 ( \2105 , \2103 , \2104 );
and \U$1763 ( \2106 , \2102 , \454 );
nor \U$1764 ( \2107 , \2105 , \2106 );
not \U$1765 ( \2108 , \2107 );
and \U$1766 ( \2109 , \438 , RI986f430_51);
and \U$1767 ( \2110 , RI986f340_49, \436 );
nor \U$1768 ( \2111 , \2109 , \2110 );
and \U$1769 ( \2112 , \2111 , \444 );
not \U$1770 ( \2113 , \2111 );
and \U$1771 ( \2114 , \2113 , \443 );
nor \U$1772 ( \2115 , \2112 , \2114 );
not \U$1773 ( \2116 , \2115 );
or \U$1774 ( \2117 , \2108 , \2116 );
or \U$1775 ( \2118 , \2107 , \2115 );
nand \U$1776 ( \2119 , \2117 , \2118 );
not \U$1777 ( \2120 , \2119 );
and \U$1778 ( \2121 , \376 , RI986f7f0_59);
and \U$1779 ( \2122 , RI986f700_57, \374 );
nor \U$1780 ( \2123 , \2121 , \2122 );
not \U$1781 ( \2124 , \2123 );
not \U$1782 ( \2125 , \365 );
and \U$1783 ( \2126 , \2124 , \2125 );
and \U$1784 ( \2127 , \2123 , \365 );
nor \U$1785 ( \2128 , \2126 , \2127 );
not \U$1786 ( \2129 , \2128 );
and \U$1787 ( \2130 , \2120 , \2129 );
and \U$1788 ( \2131 , \2119 , \2128 );
nor \U$1789 ( \2132 , \2130 , \2131 );
and \U$1790 ( \2133 , \416 , RI986f250_47);
and \U$1791 ( \2134 , RI986f160_45, \414 );
nor \U$1792 ( \2135 , \2133 , \2134 );
and \U$1793 ( \2136 , \2135 , \421 );
not \U$1794 ( \2137 , \2135 );
and \U$1795 ( \2138 , \2137 , \422 );
nor \U$1796 ( \2139 , \2136 , \2138 );
and \U$1797 ( \2140 , \395 , RI986e710_23);
and \U$1798 ( \2141 , RI986e620_21, \393 );
nor \U$1799 ( \2142 , \2140 , \2141 );
not \U$1800 ( \2143 , \2142 );
not \U$1801 ( \2144 , \386 );
and \U$1802 ( \2145 , \2143 , \2144 );
and \U$1803 ( \2146 , \2142 , \386 );
nor \U$1804 ( \2147 , \2145 , \2146 );
xor \U$1805 ( \2148 , \2139 , \2147 );
and \U$1806 ( \2149 , \354 , RI986e530_19);
and \U$1807 ( \2150 , RI986e440_17, \352 );
nor \U$1808 ( \2151 , \2149 , \2150 );
not \U$1809 ( \2152 , \2151 );
not \U$1810 ( \2153 , \345 );
and \U$1811 ( \2154 , \2152 , \2153 );
and \U$1812 ( \2155 , \2151 , \345 );
nor \U$1813 ( \2156 , \2154 , \2155 );
xor \U$1814 ( \2157 , \2148 , \2156 );
xor \U$1815 ( \2158 , \2132 , \2157 );
and \U$1816 ( \2159 , \1293 , RI986df90_7);
and \U$1817 ( \2160 , RI986dea0_5, \1291 );
nor \U$1818 ( \2161 , \2159 , \2160 );
not \U$1819 ( \2162 , \2161 );
not \U$1820 ( \2163 , \1301 );
and \U$1821 ( \2164 , \2162 , \2163 );
and \U$1822 ( \2165 , \2161 , \1301 );
nor \U$1823 ( \2166 , \2164 , \2165 );
and \U$1824 ( \2167 , \1329 , RI986ddb0_3);
and \U$1825 ( \2168 , RI986dcc0_1, \1327 );
nor \U$1826 ( \2169 , \2167 , \2168 );
and \U$1827 ( \2170 , \2169 , \1337 );
not \U$1828 ( \2171 , \2169 );
and \U$1829 ( \2172 , \2171 , \1336 );
nor \U$1830 ( \2173 , \2170 , \2172 );
xor \U$1831 ( \2174 , \2166 , \2173 );
and \U$1832 ( \2175 , \776 , RI986f520_53);
and \U$1833 ( \2176 , RI986f610_55, \774 );
nor \U$1834 ( \2177 , \2175 , \2176 );
and \U$1835 ( \2178 , \2177 , \451 );
not \U$1836 ( \2179 , \2177 );
and \U$1837 ( \2180 , \2179 , \474 );
nor \U$1838 ( \2181 , \2178 , \2180 );
xor \U$1839 ( \2182 , \2174 , \2181 );
xor \U$1840 ( \2183 , \2158 , \2182 );
xor \U$1841 ( \2184 , \2099 , \2183 );
not \U$1842 ( \2185 , \2184 );
and \U$1843 ( \2186 , \395 , RI986e530_19);
and \U$1844 ( \2187 , RI986e440_17, \393 );
nor \U$1845 ( \2188 , \2186 , \2187 );
not \U$1846 ( \2189 , \2188 );
not \U$1847 ( \2190 , \487 );
and \U$1848 ( \2191 , \2189 , \2190 );
and \U$1849 ( \2192 , \2188 , \487 );
nor \U$1850 ( \2193 , \2191 , \2192 );
and \U$1851 ( \2194 , \354 , RI986f250_47);
and \U$1852 ( \2195 , RI986f160_45, \352 );
nor \U$1853 ( \2196 , \2194 , \2195 );
not \U$1854 ( \2197 , \2196 );
not \U$1855 ( \2198 , \361 );
and \U$1856 ( \2199 , \2197 , \2198 );
and \U$1857 ( \2200 , \2196 , \345 );
nor \U$1858 ( \2201 , \2199 , \2200 );
or \U$1859 ( \2202 , \2193 , \2201 );
not \U$1860 ( \2203 , \2201 );
not \U$1861 ( \2204 , \2193 );
or \U$1862 ( \2205 , \2203 , \2204 );
not \U$1863 ( \2206 , \365 );
and \U$1864 ( \2207 , \376 , RI986e710_23);
and \U$1865 ( \2208 , RI986e620_21, \374 );
nor \U$1866 ( \2209 , \2207 , \2208 );
not \U$1867 ( \2210 , \2209 );
or \U$1868 ( \2211 , \2206 , \2210 );
or \U$1869 ( \2212 , \2209 , \367 );
nand \U$1870 ( \2213 , \2211 , \2212 );
nand \U$1871 ( \2214 , \2205 , \2213 );
nand \U$1872 ( \2215 , \2202 , \2214 );
xor \U$1873 ( \2216 , \2215 , \2066 );
not \U$1874 ( \2217 , \2084 );
xor \U$1875 ( \2218 , \2095 , \2076 );
not \U$1876 ( \2219 , \2218 );
or \U$1877 ( \2220 , \2217 , \2219 );
or \U$1878 ( \2221 , \2218 , \2084 );
nand \U$1879 ( \2222 , \2220 , \2221 );
and \U$1880 ( \2223 , \2216 , \2222 );
and \U$1881 ( \2224 , \2215 , \2066 );
or \U$1882 ( \2225 , \2223 , \2224 );
and \U$1883 ( \2226 , \438 , RI986f9d0_63);
and \U$1884 ( \2227 , RI986f8e0_61, \436 );
nor \U$1885 ( \2228 , \2226 , \2227 );
and \U$1886 ( \2229 , \2228 , \443 );
not \U$1887 ( \2230 , \2228 );
and \U$1888 ( \2231 , \2230 , \444 );
nor \U$1889 ( \2232 , \2229 , \2231 );
and \U$1890 ( \2233 , \465 , RI986f7f0_59);
and \U$1891 ( \2234 , RI986f700_57, \463 );
nor \U$1892 ( \2235 , \2233 , \2234 );
not \U$1893 ( \2236 , \2235 );
not \U$1894 ( \2237 , \454 );
and \U$1895 ( \2238 , \2236 , \2237 );
and \U$1896 ( \2239 , \2235 , \454 );
nor \U$1897 ( \2240 , \2238 , \2239 );
or \U$1898 ( \2241 , \2232 , \2240 );
not \U$1899 ( \2242 , \2240 );
not \U$1900 ( \2243 , \2232 );
or \U$1901 ( \2244 , \2242 , \2243 );
and \U$1902 ( \2245 , \776 , RI986f430_51);
and \U$1903 ( \2246 , RI986f340_49, \774 );
nor \U$1904 ( \2247 , \2245 , \2246 );
and \U$1905 ( \2248 , \2247 , \474 );
not \U$1906 ( \2249 , \2247 );
and \U$1907 ( \2250 , \2249 , \451 );
nor \U$1908 ( \2251 , \2248 , \2250 );
nand \U$1909 ( \2252 , \2244 , \2251 );
nand \U$1910 ( \2253 , \2241 , \2252 );
and \U$1911 ( \2254 , \2042 , RI986e170_11);
and \U$1912 ( \2255 , RI986e080_9, \2040 );
nor \U$1913 ( \2256 , \2254 , \2255 );
not \U$1914 ( \2257 , \2256 );
not \U$1915 ( \2258 , \1462 );
and \U$1916 ( \2259 , \2257 , \2258 );
and \U$1917 ( \2260 , \2256 , \2034 );
nor \U$1918 ( \2261 , \2259 , \2260 );
nand \U$1919 ( \2262 , RI98725e0_157, RI9872658_158);
and \U$1920 ( \2263 , \2262 , RI98726d0_159);
or \U$1921 ( \2264 , \2261 , \2263 );
not \U$1922 ( \2265 , \2263 );
not \U$1923 ( \2266 , \2261 );
or \U$1924 ( \2267 , \2265 , \2266 );
and \U$1925 ( \2268 , RI9872310_151, RI9872748_160);
not \U$1926 ( \2269 , RI98726d0_159);
and \U$1927 ( \2270 , \2269 , RI9872748_160);
nor \U$1928 ( \2271 , \2269 , RI9872748_160);
or \U$1929 ( \2272 , \2270 , \2271 );
nor \U$1930 ( \2273 , RI9872310_151, RI9872748_160);
nor \U$1931 ( \2274 , \2268 , \2272 , \2273 );
and \U$1932 ( \2275 , \2274 , RI986e260_13);
and \U$1933 ( \2276 , RI986e350_15, \2272 );
nor \U$1934 ( \2277 , \2275 , \2276 );
and \U$1935 ( \2278 , \2277 , \2030 );
not \U$1936 ( \2279 , \2277 );
and \U$1937 ( \2280 , \2279 , \2031 );
nor \U$1938 ( \2281 , \2278 , \2280 );
nand \U$1939 ( \2282 , \2267 , \2281 );
nand \U$1940 ( \2283 , \2264 , \2282 );
xor \U$1941 ( \2284 , \2253 , \2283 );
and \U$1942 ( \2285 , \1293 , RI986f520_53);
and \U$1943 ( \2286 , RI986f610_55, \1291 );
nor \U$1944 ( \2287 , \2285 , \2286 );
not \U$1945 ( \2288 , \2287 );
not \U$1946 ( \2289 , \1301 );
and \U$1947 ( \2290 , \2288 , \2289 );
and \U$1948 ( \2291 , \2287 , \1301 );
nor \U$1949 ( \2292 , \2290 , \2291 );
and \U$1950 ( \2293 , \1329 , RI986df90_7);
and \U$1951 ( \2294 , RI986dea0_5, \1327 );
nor \U$1952 ( \2295 , \2293 , \2294 );
and \U$1953 ( \2296 , \2295 , \1337 );
not \U$1954 ( \2297 , \2295 );
and \U$1955 ( \2298 , \2297 , \1336 );
nor \U$1956 ( \2299 , \2296 , \2298 );
or \U$1957 ( \2300 , \2292 , \2299 );
not \U$1958 ( \2301 , \2299 );
not \U$1959 ( \2302 , \2292 );
or \U$1960 ( \2303 , \2301 , \2302 );
and \U$1961 ( \2304 , \1311 , RI986ddb0_3);
and \U$1962 ( \2305 , RI986dcc0_1, \1309 );
nor \U$1963 ( \2306 , \2304 , \2305 );
and \U$1964 ( \2307 , \2306 , \1458 );
not \U$1965 ( \2308 , \2306 );
and \U$1966 ( \2309 , \2308 , \1318 );
nor \U$1967 ( \2310 , \2307 , \2309 );
nand \U$1968 ( \2311 , \2303 , \2310 );
nand \U$1969 ( \2312 , \2300 , \2311 );
and \U$1970 ( \2313 , \2284 , \2312 );
and \U$1971 ( \2314 , \2253 , \2283 );
or \U$1972 ( \2315 , \2313 , \2314 );
xor \U$1973 ( \2316 , \2225 , \2315 );
and \U$1974 ( \2317 , \776 , RI986f340_49);
and \U$1975 ( \2318 , RI986f520_53, \774 );
nor \U$1976 ( \2319 , \2317 , \2318 );
and \U$1977 ( \2320 , \2319 , \451 );
not \U$1978 ( \2321 , \2319 );
and \U$1979 ( \2322 , \2321 , \474 );
nor \U$1980 ( \2323 , \2320 , \2322 );
not \U$1981 ( \2324 , \2323 );
and \U$1982 ( \2325 , \1293 , RI986f610_55);
and \U$1983 ( \2326 , RI986df90_7, \1291 );
nor \U$1984 ( \2327 , \2325 , \2326 );
not \U$1985 ( \2328 , \2327 );
not \U$1986 ( \2329 , \1301 );
and \U$1987 ( \2330 , \2328 , \2329 );
and \U$1988 ( \2331 , \2327 , \1301 );
nor \U$1989 ( \2332 , \2330 , \2331 );
and \U$1990 ( \2333 , \1329 , RI986dea0_5);
and \U$1991 ( \2334 , RI986ddb0_3, \1327 );
nor \U$1992 ( \2335 , \2333 , \2334 );
and \U$1993 ( \2336 , \2335 , \1337 );
not \U$1994 ( \2337 , \2335 );
and \U$1995 ( \2338 , \2337 , \1336 );
nor \U$1996 ( \2339 , \2336 , \2338 );
xor \U$1997 ( \2340 , \2332 , \2339 );
not \U$1998 ( \2341 , \2340 );
or \U$1999 ( \2342 , \2324 , \2341 );
or \U$2000 ( \2343 , \2340 , \2323 );
nand \U$2001 ( \2344 , \2342 , \2343 );
and \U$2002 ( \2345 , \1311 , RI986dcc0_1);
and \U$2003 ( \2346 , RI986e170_11, \1309 );
nor \U$2004 ( \2347 , \2345 , \2346 );
and \U$2005 ( \2348 , \2347 , \1315 );
not \U$2006 ( \2349 , \2347 );
and \U$2007 ( \2350 , \2349 , \1458 );
nor \U$2008 ( \2351 , \2348 , \2350 );
not \U$2009 ( \2352 , \2351 );
nand \U$2010 ( \2353 , RI986e350_15, \2274 );
and \U$2011 ( \2354 , \2353 , \2031 );
not \U$2012 ( \2355 , \2353 );
and \U$2013 ( \2356 , \2355 , \2030 );
nor \U$2014 ( \2357 , \2354 , \2356 );
and \U$2015 ( \2358 , \2042 , RI986e080_9);
and \U$2016 ( \2359 , RI986e260_13, \2040 );
nor \U$2017 ( \2360 , \2358 , \2359 );
not \U$2018 ( \2361 , \2360 );
not \U$2019 ( \2362 , \1462 );
and \U$2020 ( \2363 , \2361 , \2362 );
and \U$2021 ( \2364 , \2360 , \2034 );
nor \U$2022 ( \2365 , \2363 , \2364 );
xor \U$2023 ( \2366 , \2357 , \2365 );
not \U$2024 ( \2367 , \2366 );
or \U$2025 ( \2368 , \2352 , \2367 );
or \U$2026 ( \2369 , \2366 , \2351 );
nand \U$2027 ( \2370 , \2368 , \2369 );
xor \U$2028 ( \2371 , \2344 , \2370 );
and \U$2029 ( \2372 , \376 , RI986e620_21);
and \U$2030 ( \2373 , RI986f7f0_59, \374 );
nor \U$2031 ( \2374 , \2372 , \2373 );
not \U$2032 ( \2375 , \2374 );
not \U$2033 ( \2376 , \367 );
and \U$2034 ( \2377 , \2375 , \2376 );
and \U$2035 ( \2378 , \2374 , \367 );
nor \U$2036 ( \2379 , \2377 , \2378 );
not \U$2037 ( \2380 , \2379 );
and \U$2038 ( \2381 , \465 , RI986f700_57);
and \U$2039 ( \2382 , RI986f9d0_63, \463 );
nor \U$2040 ( \2383 , \2381 , \2382 );
not \U$2041 ( \2384 , \2383 );
not \U$2042 ( \2385 , \456 );
and \U$2043 ( \2386 , \2384 , \2385 );
and \U$2044 ( \2387 , \2383 , \454 );
nor \U$2045 ( \2388 , \2386 , \2387 );
and \U$2046 ( \2389 , \438 , RI986f8e0_61);
and \U$2047 ( \2390 , RI986f430_51, \436 );
nor \U$2048 ( \2391 , \2389 , \2390 );
and \U$2049 ( \2392 , \2391 , \443 );
not \U$2050 ( \2393 , \2391 );
and \U$2051 ( \2394 , \2393 , \444 );
nor \U$2052 ( \2395 , \2392 , \2394 );
xor \U$2053 ( \2396 , \2388 , \2395 );
not \U$2054 ( \2397 , \2396 );
or \U$2055 ( \2398 , \2380 , \2397 );
or \U$2056 ( \2399 , \2396 , \2379 );
nand \U$2057 ( \2400 , \2398 , \2399 );
and \U$2058 ( \2401 , \2371 , \2400 );
and \U$2059 ( \2402 , \2344 , \2370 );
or \U$2060 ( \2403 , \2401 , \2402 );
xor \U$2061 ( \2404 , \2316 , \2403 );
nand \U$2062 ( \2405 , \2185 , \2404 );
not \U$2063 ( \2406 , \2323 );
not \U$2064 ( \2407 , \2332 );
and \U$2065 ( \2408 , \2406 , \2407 );
and \U$2066 ( \2409 , \2332 , \2323 );
nor \U$2067 ( \2410 , \2409 , \2339 );
nor \U$2068 ( \2411 , \2408 , \2410 );
not \U$2069 ( \2412 , \2388 );
not \U$2070 ( \2413 , \2379 );
and \U$2071 ( \2414 , \2412 , \2413 );
and \U$2072 ( \2415 , \2388 , \2379 );
nor \U$2073 ( \2416 , \2415 , \2395 );
nor \U$2074 ( \2417 , \2414 , \2416 );
xor \U$2075 ( \2418 , \2411 , \2417 );
not \U$2076 ( \2419 , \2351 );
not \U$2077 ( \2420 , \2365 );
and \U$2078 ( \2421 , \2419 , \2420 );
and \U$2079 ( \2422 , \2365 , \2351 );
nor \U$2080 ( \2423 , \2422 , \2357 );
nor \U$2081 ( \2424 , \2421 , \2423 );
and \U$2082 ( \2425 , \2418 , \2424 );
and \U$2083 ( \2426 , \2411 , \2417 );
or \U$2084 ( \2427 , \2425 , \2426 );
xor \U$2085 ( \2428 , \2066 , \2067 );
and \U$2086 ( \2429 , \2428 , \2097 );
and \U$2087 ( \2430 , \2066 , \2067 );
or \U$2088 ( \2431 , \2429 , \2430 );
xor \U$2089 ( \2432 , \2427 , \2431 );
xor \U$2090 ( \2433 , \2132 , \2157 );
and \U$2091 ( \2434 , \2433 , \2182 );
and \U$2092 ( \2435 , \2132 , \2157 );
or \U$2093 ( \2436 , \2434 , \2435 );
xor \U$2094 ( \2437 , \2432 , \2436 );
xor \U$2095 ( \2438 , \2405 , \2437 );
and \U$2096 ( \2439 , \2042 , RI986dcc0_1);
and \U$2097 ( \2440 , RI986e170_11, \2040 );
nor \U$2098 ( \2441 , \2439 , \2440 );
not \U$2099 ( \2442 , \2441 );
not \U$2100 ( \2443 , \1462 );
and \U$2101 ( \2444 , \2442 , \2443 );
and \U$2102 ( \2445 , \2441 , \2034 );
nor \U$2103 ( \2446 , \2444 , \2445 );
not \U$2104 ( \2447 , \2446 );
and \U$2105 ( \2448 , \2274 , RI986e080_9);
and \U$2106 ( \2449 , RI986e260_13, \2272 );
nor \U$2107 ( \2450 , \2448 , \2449 );
and \U$2108 ( \2451 , \2450 , \2031 );
not \U$2109 ( \2452 , \2450 );
and \U$2110 ( \2453 , \2452 , \2030 );
nor \U$2111 ( \2454 , \2451 , \2453 );
not \U$2112 ( \2455 , \2454 );
and \U$2113 ( \2456 , \2447 , \2455 );
and \U$2114 ( \2457 , \2454 , \2446 );
and \U$2115 ( \2458 , RI98726d0_159, RI9872658_158);
not \U$2116 ( \2459 , RI98725e0_157);
and \U$2117 ( \2460 , \2459 , RI9872658_158);
nor \U$2118 ( \2461 , \2459 , RI9872658_158);
or \U$2119 ( \2462 , \2460 , \2461 );
nor \U$2120 ( \2463 , RI98726d0_159, RI9872658_158);
nor \U$2121 ( \2464 , \2458 , \2462 , \2463 );
nand \U$2122 ( \2465 , RI986e350_15, \2464 );
and \U$2123 ( \2466 , \2465 , \2263 );
not \U$2124 ( \2467 , \2465 );
not \U$2125 ( \2468 , \2263 );
and \U$2126 ( \2469 , \2467 , \2468 );
nor \U$2127 ( \2470 , \2466 , \2469 );
nor \U$2128 ( \2471 , \2457 , \2470 );
nor \U$2129 ( \2472 , \2456 , \2471 );
and \U$2130 ( \2473 , \776 , RI986f8e0_61);
and \U$2131 ( \2474 , RI986f430_51, \774 );
nor \U$2132 ( \2475 , \2473 , \2474 );
and \U$2133 ( \2476 , \2475 , \474 );
not \U$2134 ( \2477 , \2475 );
and \U$2135 ( \2478 , \2477 , \451 );
nor \U$2136 ( \2479 , \2476 , \2478 );
and \U$2137 ( \2480 , \438 , RI986f700_57);
and \U$2138 ( \2481 , RI986f9d0_63, \436 );
nor \U$2139 ( \2482 , \2480 , \2481 );
and \U$2140 ( \2483 , \2482 , \444 );
not \U$2141 ( \2484 , \2482 );
and \U$2142 ( \2485 , \2484 , \443 );
nor \U$2143 ( \2486 , \2483 , \2485 );
xor \U$2144 ( \2487 , \2479 , \2486 );
not \U$2145 ( \2488 , \454 );
and \U$2146 ( \2489 , \465 , RI986e620_21);
and \U$2147 ( \2490 , RI986f7f0_59, \463 );
nor \U$2148 ( \2491 , \2489 , \2490 );
not \U$2149 ( \2492 , \2491 );
or \U$2150 ( \2493 , \2488 , \2492 );
or \U$2151 ( \2494 , \2491 , \454 );
nand \U$2152 ( \2495 , \2493 , \2494 );
and \U$2153 ( \2496 , \2487 , \2495 );
and \U$2154 ( \2497 , \2479 , \2486 );
nor \U$2155 ( \2498 , \2496 , \2497 );
or \U$2156 ( \2499 , \2472 , \2498 );
not \U$2157 ( \2500 , \2472 );
not \U$2158 ( \2501 , \2498 );
or \U$2159 ( \2502 , \2500 , \2501 );
not \U$2160 ( \2503 , \1301 );
and \U$2161 ( \2504 , \1293 , RI986f340_49);
and \U$2162 ( \2505 , RI986f520_53, \1291 );
nor \U$2163 ( \2506 , \2504 , \2505 );
not \U$2164 ( \2507 , \2506 );
or \U$2165 ( \2508 , \2503 , \2507 );
or \U$2166 ( \2509 , \2506 , \1128 );
nand \U$2167 ( \2510 , \2508 , \2509 );
and \U$2168 ( \2511 , \1329 , RI986f610_55);
and \U$2169 ( \2512 , RI986df90_7, \1327 );
nor \U$2170 ( \2513 , \2511 , \2512 );
and \U$2171 ( \2514 , \2513 , \1336 );
not \U$2172 ( \2515 , \2513 );
and \U$2173 ( \2516 , \2515 , \1337 );
nor \U$2174 ( \2517 , \2514 , \2516 );
xor \U$2175 ( \2518 , \2510 , \2517 );
and \U$2176 ( \2519 , \1311 , RI986dea0_5);
and \U$2177 ( \2520 , RI986ddb0_3, \1309 );
nor \U$2178 ( \2521 , \2519 , \2520 );
and \U$2179 ( \2522 , \2521 , \1458 );
not \U$2180 ( \2523 , \2521 );
and \U$2181 ( \2524 , \2523 , \1318 );
nor \U$2182 ( \2525 , \2522 , \2524 );
and \U$2183 ( \2526 , \2518 , \2525 );
and \U$2184 ( \2527 , \2510 , \2517 );
or \U$2185 ( \2528 , \2526 , \2527 );
nand \U$2186 ( \2529 , \2502 , \2528 );
nand \U$2187 ( \2530 , \2499 , \2529 );
nand \U$2188 ( \2531 , RI986ebc0_33, RI9871fc8_144);
and \U$2189 ( \2532 , \416 , RI986ecb0_35);
and \U$2190 ( \2533 , RI986f070_43, \414 );
nor \U$2191 ( \2534 , \2532 , \2533 );
and \U$2192 ( \2535 , \2534 , \421 );
not \U$2193 ( \2536 , \2534 );
and \U$2194 ( \2537 , \2536 , \422 );
nor \U$2195 ( \2538 , \2535 , \2537 );
nand \U$2196 ( \2539 , \2531 , \2538 );
and \U$2197 ( \2540 , \416 , RI986f070_43);
and \U$2198 ( \2541 , RI986ef80_41, \414 );
nor \U$2199 ( \2542 , \2540 , \2541 );
and \U$2200 ( \2543 , \2542 , \422 );
not \U$2201 ( \2544 , \2542 );
and \U$2202 ( \2545 , \2544 , \421 );
nor \U$2203 ( \2546 , \2543 , \2545 );
xor \U$2204 ( \2547 , \2539 , \2546 );
not \U$2205 ( \2548 , \386 );
and \U$2206 ( \2549 , \395 , RI986f160_45);
and \U$2207 ( \2550 , RI986e530_19, \393 );
nor \U$2208 ( \2551 , \2549 , \2550 );
not \U$2209 ( \2552 , \2551 );
or \U$2210 ( \2553 , \2548 , \2552 );
or \U$2211 ( \2554 , \2551 , \487 );
nand \U$2212 ( \2555 , \2553 , \2554 );
not \U$2213 ( \2556 , \365 );
and \U$2214 ( \2557 , \376 , RI986e440_17);
and \U$2215 ( \2558 , RI986e710_23, \374 );
nor \U$2216 ( \2559 , \2557 , \2558 );
not \U$2217 ( \2560 , \2559 );
or \U$2218 ( \2561 , \2556 , \2560 );
or \U$2219 ( \2562 , \2559 , \367 );
nand \U$2220 ( \2563 , \2561 , \2562 );
xor \U$2221 ( \2564 , \2555 , \2563 );
not \U$2222 ( \2565 , \361 );
and \U$2223 ( \2566 , \354 , RI986ef80_41);
and \U$2224 ( \2567 , RI986f250_47, \352 );
nor \U$2225 ( \2568 , \2566 , \2567 );
not \U$2226 ( \2569 , \2568 );
or \U$2227 ( \2570 , \2565 , \2569 );
or \U$2228 ( \2571 , \2568 , \345 );
nand \U$2229 ( \2572 , \2570 , \2571 );
and \U$2230 ( \2573 , \2564 , \2572 );
and \U$2231 ( \2574 , \2555 , \2563 );
or \U$2232 ( \2575 , \2573 , \2574 );
and \U$2233 ( \2576 , \2547 , \2575 );
and \U$2234 ( \2577 , \2539 , \2546 );
or \U$2235 ( \2578 , \2576 , \2577 );
and \U$2236 ( \2579 , \2530 , \2578 );
not \U$2237 ( \2580 , \2530 );
not \U$2238 ( \2581 , \2578 );
and \U$2239 ( \2582 , \2580 , \2581 );
not \U$2240 ( \2583 , \2232 );
not \U$2241 ( \2584 , \2251 );
or \U$2242 ( \2585 , \2583 , \2584 );
or \U$2243 ( \2586 , \2232 , \2251 );
nand \U$2244 ( \2587 , \2585 , \2586 );
not \U$2245 ( \2588 , \2587 );
not \U$2246 ( \2589 , \2240 );
and \U$2247 ( \2590 , \2588 , \2589 );
and \U$2248 ( \2591 , \2587 , \2240 );
nor \U$2249 ( \2592 , \2590 , \2591 );
nand \U$2250 ( \2593 , RI986ecb0_35, RI9871fc8_144);
xor \U$2251 ( \2594 , \2592 , \2593 );
not \U$2252 ( \2595 , \2193 );
not \U$2253 ( \2596 , \2213 );
or \U$2254 ( \2597 , \2595 , \2596 );
or \U$2255 ( \2598 , \2193 , \2213 );
nand \U$2256 ( \2599 , \2597 , \2598 );
not \U$2257 ( \2600 , \2599 );
not \U$2258 ( \2601 , \2201 );
and \U$2259 ( \2602 , \2600 , \2601 );
and \U$2260 ( \2603 , \2599 , \2201 );
nor \U$2261 ( \2604 , \2602 , \2603 );
and \U$2262 ( \2605 , \2594 , \2604 );
and \U$2263 ( \2606 , \2592 , \2593 );
or \U$2264 ( \2607 , \2605 , \2606 );
nor \U$2265 ( \2608 , \2582 , \2607 );
nor \U$2266 ( \2609 , \2579 , \2608 );
not \U$2267 ( \2610 , \2609 );
xor \U$2268 ( \2611 , \2411 , \2417 );
xor \U$2269 ( \2612 , \2611 , \2424 );
not \U$2270 ( \2613 , \2612 );
and \U$2271 ( \2614 , \2610 , \2613 );
and \U$2272 ( \2615 , \2609 , \2612 );
xor \U$2273 ( \2616 , \2215 , \2066 );
xor \U$2274 ( \2617 , \2616 , \2222 );
xor \U$2275 ( \2618 , \2253 , \2283 );
xor \U$2276 ( \2619 , \2618 , \2312 );
xor \U$2277 ( \2620 , \2617 , \2619 );
xor \U$2278 ( \2621 , \2344 , \2370 );
xor \U$2279 ( \2622 , \2621 , \2400 );
and \U$2280 ( \2623 , \2620 , \2622 );
and \U$2281 ( \2624 , \2617 , \2619 );
nor \U$2282 ( \2625 , \2623 , \2624 );
nor \U$2283 ( \2626 , \2615 , \2625 );
nor \U$2284 ( \2627 , \2614 , \2626 );
and \U$2285 ( \2628 , \2438 , \2627 );
and \U$2286 ( \2629 , \2405 , \2437 );
or \U$2287 ( \2630 , \2628 , \2629 );
not \U$2288 ( \2631 , \2630 );
xor \U$2289 ( \2632 , \2225 , \2315 );
and \U$2290 ( \2633 , \2632 , \2403 );
and \U$2291 ( \2634 , \2225 , \2315 );
or \U$2292 ( \2635 , \2633 , \2634 );
xor \U$2293 ( \2636 , \2065 , \2098 );
and \U$2294 ( \2637 , \2636 , \2183 );
and \U$2295 ( \2638 , \2065 , \2098 );
nor \U$2296 ( \2639 , \2637 , \2638 );
xor \U$2297 ( \2640 , \2635 , \2639 );
or \U$2298 ( \2641 , \2107 , \2128 );
not \U$2299 ( \2642 , \2128 );
not \U$2300 ( \2643 , \2107 );
or \U$2301 ( \2644 , \2642 , \2643 );
nand \U$2302 ( \2645 , \2644 , \2115 );
nand \U$2303 ( \2646 , \2641 , \2645 );
or \U$2304 ( \2647 , \2061 , \2031 );
not \U$2305 ( \2648 , \2031 );
not \U$2306 ( \2649 , \2061 );
or \U$2307 ( \2650 , \2648 , \2649 );
nand \U$2308 ( \2651 , \2650 , \2049 );
nand \U$2309 ( \2652 , \2647 , \2651 );
xor \U$2310 ( \2653 , \2646 , \2652 );
xor \U$2311 ( \2654 , \2166 , \2173 );
and \U$2312 ( \2655 , \2654 , \2181 );
and \U$2313 ( \2656 , \2166 , \2173 );
nor \U$2314 ( \2657 , \2655 , \2656 );
xor \U$2315 ( \2658 , \2653 , \2657 );
and \U$2316 ( \2659 , \354 , RI986e440_17);
and \U$2317 ( \2660 , RI986e710_23, \352 );
nor \U$2318 ( \2661 , \2659 , \2660 );
not \U$2319 ( \2662 , \2661 );
not \U$2320 ( \2663 , \361 );
and \U$2321 ( \2664 , \2662 , \2663 );
and \U$2322 ( \2665 , \2661 , \361 );
nor \U$2323 ( \2666 , \2664 , \2665 );
nand \U$2324 ( \2667 , RI986f250_47, RI9871fc8_144);
xor \U$2325 ( \2668 , \2666 , \2667 );
and \U$2326 ( \2669 , \416 , RI986f160_45);
and \U$2327 ( \2670 , RI986e530_19, \414 );
nor \U$2328 ( \2671 , \2669 , \2670 );
and \U$2329 ( \2672 , \2671 , \421 );
not \U$2330 ( \2673 , \2671 );
and \U$2331 ( \2674 , \2673 , \422 );
nor \U$2332 ( \2675 , \2672 , \2674 );
xor \U$2333 ( \2676 , \2668 , \2675 );
xor \U$2334 ( \2677 , \2139 , \2147 );
and \U$2335 ( \2678 , \2677 , \2156 );
and \U$2336 ( \2679 , \2139 , \2147 );
or \U$2337 ( \2680 , \2678 , \2679 );
or \U$2338 ( \2681 , \2676 , \2680 );
nand \U$2339 ( \2682 , \2680 , \2676 );
nand \U$2340 ( \2683 , \2681 , \2682 );
and \U$2341 ( \2684 , \776 , RI986f610_55);
and \U$2342 ( \2685 , RI986df90_7, \774 );
nor \U$2343 ( \2686 , \2684 , \2685 );
and \U$2344 ( \2687 , \2686 , \474 );
not \U$2345 ( \2688 , \2686 );
and \U$2346 ( \2689 , \2688 , \451 );
nor \U$2347 ( \2690 , \2687 , \2689 );
not \U$2348 ( \2691 , \1301 );
and \U$2349 ( \2692 , \1293 , RI986dea0_5);
and \U$2350 ( \2693 , RI986ddb0_3, \1291 );
nor \U$2351 ( \2694 , \2692 , \2693 );
not \U$2352 ( \2695 , \2694 );
or \U$2353 ( \2696 , \2691 , \2695 );
or \U$2354 ( \2697 , \2694 , \1128 );
nand \U$2355 ( \2698 , \2696 , \2697 );
xor \U$2356 ( \2699 , \2690 , \2698 );
and \U$2357 ( \2700 , \438 , RI986f340_49);
and \U$2358 ( \2701 , RI986f520_53, \436 );
nor \U$2359 ( \2702 , \2700 , \2701 );
and \U$2360 ( \2703 , \2702 , \444 );
not \U$2361 ( \2704 , \2702 );
and \U$2362 ( \2705 , \2704 , \443 );
nor \U$2363 ( \2706 , \2703 , \2705 );
xor \U$2364 ( \2707 , \2699 , \2706 );
and \U$2365 ( \2708 , \1329 , RI986dcc0_1);
and \U$2366 ( \2709 , RI986e170_11, \1327 );
nor \U$2367 ( \2710 , \2708 , \2709 );
and \U$2368 ( \2711 , \2710 , \1337 );
not \U$2369 ( \2712 , \2710 );
and \U$2370 ( \2713 , \2712 , \1336 );
nor \U$2371 ( \2714 , \2711 , \2713 );
not \U$2372 ( \2715 , \2714 );
nand \U$2373 ( \2716 , RI986e350_15, \2042 );
not \U$2374 ( \2717 , \2716 );
not \U$2375 ( \2718 , \2034 );
and \U$2376 ( \2719 , \2717 , \2718 );
and \U$2377 ( \2720 , \2716 , \1462 );
nor \U$2378 ( \2721 , \2719 , \2720 );
and \U$2379 ( \2722 , \1311 , RI986e080_9);
and \U$2380 ( \2723 , RI986e260_13, \1309 );
nor \U$2381 ( \2724 , \2722 , \2723 );
and \U$2382 ( \2725 , \2724 , \1315 );
not \U$2383 ( \2726 , \2724 );
and \U$2384 ( \2727 , \2726 , \1458 );
nor \U$2385 ( \2728 , \2725 , \2727 );
xor \U$2386 ( \2729 , \2721 , \2728 );
not \U$2387 ( \2730 , \2729 );
or \U$2388 ( \2731 , \2715 , \2730 );
or \U$2389 ( \2732 , \2729 , \2714 );
nand \U$2390 ( \2733 , \2731 , \2732 );
xor \U$2391 ( \2734 , \2707 , \2733 );
and \U$2392 ( \2735 , \395 , RI986e620_21);
and \U$2393 ( \2736 , RI986f7f0_59, \393 );
nor \U$2394 ( \2737 , \2735 , \2736 );
not \U$2395 ( \2738 , \2737 );
not \U$2396 ( \2739 , \386 );
and \U$2397 ( \2740 , \2738 , \2739 );
and \U$2398 ( \2741 , \2737 , \386 );
nor \U$2399 ( \2742 , \2740 , \2741 );
not \U$2400 ( \2743 , \2742 );
and \U$2401 ( \2744 , \465 , RI986f8e0_61);
and \U$2402 ( \2745 , RI986f430_51, \463 );
nor \U$2403 ( \2746 , \2744 , \2745 );
not \U$2404 ( \2747 , \2746 );
not \U$2405 ( \2748 , \456 );
and \U$2406 ( \2749 , \2747 , \2748 );
and \U$2407 ( \2750 , \2746 , \456 );
nor \U$2408 ( \2751 , \2749 , \2750 );
and \U$2409 ( \2752 , \376 , RI986f700_57);
and \U$2410 ( \2753 , RI986f9d0_63, \374 );
nor \U$2411 ( \2754 , \2752 , \2753 );
not \U$2412 ( \2755 , \2754 );
not \U$2413 ( \2756 , \365 );
and \U$2414 ( \2757 , \2755 , \2756 );
and \U$2415 ( \2758 , \2754 , \365 );
nor \U$2416 ( \2759 , \2757 , \2758 );
xor \U$2417 ( \2760 , \2751 , \2759 );
not \U$2418 ( \2761 , \2760 );
or \U$2419 ( \2762 , \2743 , \2761 );
or \U$2420 ( \2763 , \2760 , \2742 );
nand \U$2421 ( \2764 , \2762 , \2763 );
xor \U$2422 ( \2765 , \2734 , \2764 );
xor \U$2423 ( \2766 , \2683 , \2765 );
xor \U$2424 ( \2767 , \2658 , \2766 );
and \U$2425 ( \2768 , \2640 , \2767 );
and \U$2426 ( \2769 , \2635 , \2639 );
or \U$2427 ( \2770 , \2768 , \2769 );
xor \U$2428 ( \2771 , \2646 , \2652 );
and \U$2429 ( \2772 , \2771 , \2657 );
and \U$2430 ( \2773 , \2646 , \2652 );
or \U$2431 ( \2774 , \2772 , \2773 );
xor \U$2432 ( \2775 , \2682 , \2774 );
xor \U$2433 ( \2776 , \2707 , \2733 );
and \U$2434 ( \2777 , \2776 , \2764 );
and \U$2435 ( \2778 , \2707 , \2733 );
or \U$2436 ( \2779 , \2777 , \2778 );
xor \U$2437 ( \2780 , \2775 , \2779 );
xor \U$2438 ( \2781 , \2770 , \2780 );
not \U$2439 ( \2782 , \2751 );
not \U$2440 ( \2783 , \2742 );
and \U$2441 ( \2784 , \2782 , \2783 );
and \U$2442 ( \2785 , \2751 , \2742 );
nor \U$2443 ( \2786 , \2785 , \2759 );
nor \U$2444 ( \2787 , \2784 , \2786 );
not \U$2445 ( \2788 , \2714 );
not \U$2446 ( \2789 , \2728 );
and \U$2447 ( \2790 , \2788 , \2789 );
and \U$2448 ( \2791 , \2728 , \2714 );
nor \U$2449 ( \2792 , \2791 , \2721 );
nor \U$2450 ( \2793 , \2790 , \2792 );
xor \U$2451 ( \2794 , \2787 , \2793 );
xor \U$2452 ( \2795 , \2690 , \2698 );
and \U$2453 ( \2796 , \2795 , \2706 );
and \U$2454 ( \2797 , \2690 , \2698 );
nor \U$2455 ( \2798 , \2796 , \2797 );
xor \U$2456 ( \2799 , \2794 , \2798 );
xor \U$2457 ( \2800 , \1460 , \1462 );
xor \U$2458 ( \2801 , \2800 , \1470 );
not \U$2459 ( \2802 , \2801 );
not \U$2460 ( \2803 , \1517 );
xor \U$2461 ( \2804 , \1509 , \1528 );
not \U$2462 ( \2805 , \2804 );
or \U$2463 ( \2806 , \2803 , \2805 );
or \U$2464 ( \2807 , \2804 , \1517 );
nand \U$2465 ( \2808 , \2806 , \2807 );
not \U$2466 ( \2809 , \2808 );
and \U$2467 ( \2810 , \2802 , \2809 );
and \U$2468 ( \2811 , \2801 , \2808 );
nor \U$2469 ( \2812 , \2810 , \2811 );
xor \U$2470 ( \2813 , \1553 , \1554 );
xor \U$2471 ( \2814 , \2813 , \1563 );
xor \U$2472 ( \2815 , \2666 , \2667 );
and \U$2473 ( \2816 , \2815 , \2675 );
and \U$2474 ( \2817 , \2666 , \2667 );
or \U$2475 ( \2818 , \2816 , \2817 );
xor \U$2476 ( \2819 , \1481 , \1489 );
xor \U$2477 ( \2820 , \2819 , \1498 );
xor \U$2478 ( \2821 , \2818 , \2820 );
xor \U$2479 ( \2822 , \2814 , \2821 );
xor \U$2480 ( \2823 , \2812 , \2822 );
xor \U$2481 ( \2824 , \2799 , \2823 );
not \U$2482 ( \2825 , \2824 );
xor \U$2483 ( \2826 , \2427 , \2431 );
and \U$2484 ( \2827 , \2826 , \2436 );
and \U$2485 ( \2828 , \2427 , \2431 );
or \U$2486 ( \2829 , \2827 , \2828 );
not \U$2487 ( \2830 , \2829 );
xor \U$2488 ( \2831 , \2646 , \2652 );
xor \U$2489 ( \2832 , \2831 , \2657 );
and \U$2490 ( \2833 , \2683 , \2832 );
xor \U$2491 ( \2834 , \2646 , \2652 );
xor \U$2492 ( \2835 , \2834 , \2657 );
and \U$2493 ( \2836 , \2765 , \2835 );
and \U$2494 ( \2837 , \2683 , \2765 );
or \U$2495 ( \2838 , \2833 , \2836 , \2837 );
not \U$2496 ( \2839 , \2838 );
or \U$2497 ( \2840 , \2830 , \2839 );
or \U$2498 ( \2841 , \2838 , \2829 );
nand \U$2499 ( \2842 , \2840 , \2841 );
not \U$2500 ( \2843 , \2842 );
or \U$2501 ( \2844 , \2825 , \2843 );
or \U$2502 ( \2845 , \2842 , \2824 );
nand \U$2503 ( \2846 , \2844 , \2845 );
xor \U$2504 ( \2847 , \2781 , \2846 );
nand \U$2505 ( \2848 , \2631 , \2847 );
not \U$2506 ( \2849 , \2824 );
not \U$2507 ( \2850 , \2829 );
and \U$2508 ( \2851 , \2849 , \2850 );
and \U$2509 ( \2852 , \2824 , \2829 );
not \U$2510 ( \2853 , \2838 );
nor \U$2511 ( \2854 , \2852 , \2853 );
nor \U$2512 ( \2855 , \2851 , \2854 );
xor \U$2513 ( \2856 , \2787 , \2793 );
and \U$2514 ( \2857 , \2856 , \2798 );
and \U$2515 ( \2858 , \2787 , \2793 );
or \U$2516 ( \2859 , \2857 , \2858 );
not \U$2517 ( \2860 , \2801 );
nand \U$2518 ( \2861 , \2860 , \2808 );
xor \U$2519 ( \2862 , \2859 , \2861 );
xor \U$2520 ( \2863 , \1553 , \1554 );
xor \U$2521 ( \2864 , \2863 , \1563 );
and \U$2522 ( \2865 , \2818 , \2864 );
xor \U$2523 ( \2866 , \1553 , \1554 );
xor \U$2524 ( \2867 , \2866 , \1563 );
and \U$2525 ( \2868 , \2820 , \2867 );
and \U$2526 ( \2869 , \2818 , \2820 );
or \U$2527 ( \2870 , \2865 , \2868 , \2869 );
xor \U$2528 ( \2871 , \2862 , \2870 );
xor \U$2529 ( \2872 , \2855 , \2871 );
xor \U$2530 ( \2873 , \2787 , \2793 );
xor \U$2531 ( \2874 , \2873 , \2798 );
and \U$2532 ( \2875 , \2812 , \2874 );
xor \U$2533 ( \2876 , \2787 , \2793 );
xor \U$2534 ( \2877 , \2876 , \2798 );
and \U$2535 ( \2878 , \2822 , \2877 );
and \U$2536 ( \2879 , \2812 , \2822 );
or \U$2537 ( \2880 , \2875 , \2878 , \2879 );
xor \U$2538 ( \2881 , \2682 , \2774 );
and \U$2539 ( \2882 , \2881 , \2779 );
and \U$2540 ( \2883 , \2682 , \2774 );
nor \U$2541 ( \2884 , \2882 , \2883 );
xor \U$2542 ( \2885 , \2880 , \2884 );
xor \U$2543 ( \2886 , \1473 , \1501 );
xor \U$2544 ( \2887 , \2886 , \1530 );
not \U$2545 ( \2888 , \1450 );
not \U$2546 ( \2889 , \1447 );
and \U$2547 ( \2890 , \2888 , \2889 );
and \U$2548 ( \2891 , \1450 , \1447 );
nor \U$2549 ( \2892 , \2890 , \2891 );
xor \U$2550 ( \2893 , \2887 , \2892 );
xnor \U$2551 ( \2894 , \1566 , \1546 );
not \U$2552 ( \2895 , \2894 );
not \U$2553 ( \2896 , \1572 );
and \U$2554 ( \2897 , \2895 , \2896 );
and \U$2555 ( \2898 , \2894 , \1572 );
nor \U$2556 ( \2899 , \2897 , \2898 );
xor \U$2557 ( \2900 , \2893 , \2899 );
xor \U$2558 ( \2901 , \2885 , \2900 );
xor \U$2559 ( \2902 , \2872 , \2901 );
not \U$2560 ( \2903 , \2902 );
xor \U$2561 ( \2904 , \2770 , \2780 );
and \U$2562 ( \2905 , \2904 , \2846 );
and \U$2563 ( \2906 , \2770 , \2780 );
or \U$2564 ( \2907 , \2905 , \2906 );
not \U$2565 ( \2908 , \2907 );
and \U$2566 ( \2909 , \2903 , \2908 );
and \U$2567 ( \2910 , \2902 , \2907 );
nor \U$2568 ( \2911 , \2909 , \2910 );
xor \U$2569 ( \2912 , \2848 , \2911 );
not \U$2570 ( \2913 , \2630 );
not \U$2571 ( \2914 , \2847 );
or \U$2572 ( \2915 , \2913 , \2914 );
or \U$2573 ( \2916 , \2847 , \2630 );
nand \U$2574 ( \2917 , \2915 , \2916 );
xor \U$2575 ( \2918 , \2405 , \2437 );
xor \U$2576 ( \2919 , \2918 , \2627 );
xor \U$2577 ( \2920 , \2635 , \2639 );
xor \U$2578 ( \2921 , \2920 , \2767 );
not \U$2579 ( \2922 , \2921 );
or \U$2580 ( \2923 , \2919 , \2922 );
not \U$2581 ( \2924 , \2922 );
not \U$2582 ( \2925 , \2919 );
or \U$2583 ( \2926 , \2924 , \2925 );
and \U$2584 ( \2927 , \2274 , RI986e170_11);
and \U$2585 ( \2928 , RI986e080_9, \2272 );
nor \U$2586 ( \2929 , \2927 , \2928 );
and \U$2587 ( \2930 , \2929 , \2031 );
not \U$2588 ( \2931 , \2929 );
and \U$2589 ( \2932 , \2931 , \2030 );
nor \U$2590 ( \2933 , \2930 , \2932 );
nand \U$2591 ( \2934 , RI9872388_152, RI98727c0_161);
and \U$2592 ( \2935 , \2934 , RI98725e0_157);
xor \U$2593 ( \2936 , \2933 , \2935 );
and \U$2594 ( \2937 , \2464 , RI986e260_13);
and \U$2595 ( \2938 , RI986e350_15, \2462 );
nor \U$2596 ( \2939 , \2937 , \2938 );
and \U$2597 ( \2940 , \2939 , \2263 );
not \U$2598 ( \2941 , \2939 );
and \U$2599 ( \2942 , \2941 , \2468 );
nor \U$2600 ( \2943 , \2940 , \2942 );
and \U$2601 ( \2944 , \2936 , \2943 );
and \U$2602 ( \2945 , \2933 , \2935 );
or \U$2603 ( \2946 , \2944 , \2945 );
and \U$2604 ( \2947 , \2042 , RI986ddb0_3);
and \U$2605 ( \2948 , RI986dcc0_1, \2040 );
nor \U$2606 ( \2949 , \2947 , \2948 );
not \U$2607 ( \2950 , \2949 );
not \U$2608 ( \2951 , \1462 );
and \U$2609 ( \2952 , \2950 , \2951 );
and \U$2610 ( \2953 , \2949 , \1462 );
nor \U$2611 ( \2954 , \2952 , \2953 );
and \U$2612 ( \2955 , \1329 , RI986f520_53);
and \U$2613 ( \2956 , RI986f610_55, \1327 );
nor \U$2614 ( \2957 , \2955 , \2956 );
and \U$2615 ( \2958 , \2957 , \1337 );
not \U$2616 ( \2959 , \2957 );
and \U$2617 ( \2960 , \2959 , \1336 );
nor \U$2618 ( \2961 , \2958 , \2960 );
xor \U$2619 ( \2962 , \2954 , \2961 );
and \U$2620 ( \2963 , \1311 , RI986df90_7);
and \U$2621 ( \2964 , RI986dea0_5, \1309 );
nor \U$2622 ( \2965 , \2963 , \2964 );
and \U$2623 ( \2966 , \2965 , \1318 );
not \U$2624 ( \2967 , \2965 );
and \U$2625 ( \2968 , \2967 , \1458 );
nor \U$2626 ( \2969 , \2966 , \2968 );
and \U$2627 ( \2970 , \2962 , \2969 );
and \U$2628 ( \2971 , \2954 , \2961 );
or \U$2629 ( \2972 , \2970 , \2971 );
xor \U$2630 ( \2973 , \2946 , \2972 );
and \U$2631 ( \2974 , \1293 , RI986f430_51);
and \U$2632 ( \2975 , RI986f340_49, \1291 );
nor \U$2633 ( \2976 , \2974 , \2975 );
not \U$2634 ( \2977 , \2976 );
not \U$2635 ( \2978 , \1301 );
and \U$2636 ( \2979 , \2977 , \2978 );
and \U$2637 ( \2980 , \2976 , \1301 );
nor \U$2638 ( \2981 , \2979 , \2980 );
and \U$2639 ( \2982 , \776 , RI986f9d0_63);
and \U$2640 ( \2983 , RI986f8e0_61, \774 );
nor \U$2641 ( \2984 , \2982 , \2983 );
and \U$2642 ( \2985 , \2984 , \451 );
not \U$2643 ( \2986 , \2984 );
and \U$2644 ( \2987 , \2986 , \474 );
nor \U$2645 ( \2988 , \2985 , \2987 );
xor \U$2646 ( \2989 , \2981 , \2988 );
and \U$2647 ( \2990 , \438 , RI986f7f0_59);
and \U$2648 ( \2991 , RI986f700_57, \436 );
nor \U$2649 ( \2992 , \2990 , \2991 );
and \U$2650 ( \2993 , \2992 , \443 );
not \U$2651 ( \2994 , \2992 );
and \U$2652 ( \2995 , \2994 , \444 );
nor \U$2653 ( \2996 , \2993 , \2995 );
and \U$2654 ( \2997 , \2989 , \2996 );
and \U$2655 ( \2998 , \2981 , \2988 );
or \U$2656 ( \2999 , \2997 , \2998 );
and \U$2657 ( \3000 , \2973 , \2999 );
and \U$2658 ( \3001 , \2946 , \2972 );
nor \U$2659 ( \3002 , \3000 , \3001 );
and \U$2660 ( \3003 , \416 , RI986ebc0_33);
and \U$2661 ( \3004 , RI986ecb0_35, \414 );
nor \U$2662 ( \3005 , \3003 , \3004 );
and \U$2663 ( \3006 , \3005 , \421 );
not \U$2664 ( \3007 , \3005 );
and \U$2665 ( \3008 , \3007 , \422 );
nor \U$2666 ( \3009 , \3006 , \3008 );
nand \U$2667 ( \3010 , RI986eda0_37, RI9871fc8_144);
or \U$2668 ( \3011 , \3009 , \3010 );
not \U$2669 ( \3012 , \3010 );
not \U$2670 ( \3013 , \3009 );
or \U$2671 ( \3014 , \3012 , \3013 );
not \U$2672 ( \3015 , \361 );
and \U$2673 ( \3016 , \354 , RI986f070_43);
and \U$2674 ( \3017 , RI986ef80_41, \352 );
nor \U$2675 ( \3018 , \3016 , \3017 );
not \U$2676 ( \3019 , \3018 );
or \U$2677 ( \3020 , \3015 , \3019 );
or \U$2678 ( \3021 , \3018 , \345 );
nand \U$2679 ( \3022 , \3020 , \3021 );
nand \U$2680 ( \3023 , \3014 , \3022 );
nand \U$2681 ( \3024 , \3011 , \3023 );
or \U$2682 ( \3025 , \2538 , \2531 );
nand \U$2683 ( \3026 , \3025 , \2539 );
xor \U$2684 ( \3027 , \3024 , \3026 );
and \U$2685 ( \3028 , \465 , RI986e710_23);
and \U$2686 ( \3029 , RI986e620_21, \463 );
nor \U$2687 ( \3030 , \3028 , \3029 );
not \U$2688 ( \3031 , \3030 );
not \U$2689 ( \3032 , \454 );
and \U$2690 ( \3033 , \3031 , \3032 );
and \U$2691 ( \3034 , \3030 , \454 );
nor \U$2692 ( \3035 , \3033 , \3034 );
and \U$2693 ( \3036 , \376 , RI986e530_19);
and \U$2694 ( \3037 , RI986e440_17, \374 );
nor \U$2695 ( \3038 , \3036 , \3037 );
not \U$2696 ( \3039 , \3038 );
not \U$2697 ( \3040 , \367 );
and \U$2698 ( \3041 , \3039 , \3040 );
and \U$2699 ( \3042 , \3038 , \365 );
nor \U$2700 ( \3043 , \3041 , \3042 );
xor \U$2701 ( \3044 , \3035 , \3043 );
and \U$2702 ( \3045 , \395 , RI986f250_47);
and \U$2703 ( \3046 , RI986f160_45, \393 );
nor \U$2704 ( \3047 , \3045 , \3046 );
not \U$2705 ( \3048 , \3047 );
not \U$2706 ( \3049 , \386 );
and \U$2707 ( \3050 , \3048 , \3049 );
and \U$2708 ( \3051 , \3047 , \386 );
nor \U$2709 ( \3052 , \3050 , \3051 );
and \U$2710 ( \3053 , \3044 , \3052 );
and \U$2711 ( \3054 , \3035 , \3043 );
nor \U$2712 ( \3055 , \3053 , \3054 );
and \U$2713 ( \3056 , \3027 , \3055 );
and \U$2714 ( \3057 , \3024 , \3026 );
or \U$2715 ( \3058 , \3056 , \3057 );
xor \U$2716 ( \3059 , \3002 , \3058 );
xor \U$2717 ( \3060 , \2479 , \2486 );
xor \U$2718 ( \3061 , \3060 , \2495 );
xor \U$2719 ( \3062 , \2510 , \2517 );
xor \U$2720 ( \3063 , \3062 , \2525 );
and \U$2721 ( \3064 , \3061 , \3063 );
xor \U$2722 ( \3065 , \2555 , \2563 );
xor \U$2723 ( \3066 , \3065 , \2572 );
xor \U$2724 ( \3067 , \2510 , \2517 );
xor \U$2725 ( \3068 , \3067 , \2525 );
and \U$2726 ( \3069 , \3066 , \3068 );
and \U$2727 ( \3070 , \3061 , \3066 );
or \U$2728 ( \3071 , \3064 , \3069 , \3070 );
and \U$2729 ( \3072 , \3059 , \3071 );
and \U$2730 ( \3073 , \3002 , \3058 );
or \U$2731 ( \3074 , \3072 , \3073 );
and \U$2732 ( \3075 , \2281 , \2468 );
not \U$2733 ( \3076 , \2281 );
and \U$2734 ( \3077 , \3076 , \2263 );
nor \U$2735 ( \3078 , \3075 , \3077 );
not \U$2736 ( \3079 , \3078 );
not \U$2737 ( \3080 , \2261 );
and \U$2738 ( \3081 , \3079 , \3080 );
and \U$2739 ( \3082 , \3078 , \2261 );
nor \U$2740 ( \3083 , \3081 , \3082 );
not \U$2741 ( \3084 , \2299 );
not \U$2742 ( \3085 , \2310 );
or \U$2743 ( \3086 , \3084 , \3085 );
or \U$2744 ( \3087 , \2299 , \2310 );
nand \U$2745 ( \3088 , \3086 , \3087 );
not \U$2746 ( \3089 , \3088 );
not \U$2747 ( \3090 , \2292 );
and \U$2748 ( \3091 , \3089 , \3090 );
and \U$2749 ( \3092 , \3088 , \2292 );
nor \U$2750 ( \3093 , \3091 , \3092 );
or \U$2751 ( \3094 , \3083 , \3093 );
and \U$2752 ( \3095 , \3083 , \3093 );
xor \U$2753 ( \3096 , \2592 , \2593 );
xor \U$2754 ( \3097 , \3096 , \2604 );
nor \U$2755 ( \3098 , \3095 , \3097 );
not \U$2756 ( \3099 , \3098 );
nand \U$2757 ( \3100 , \3094 , \3099 );
xor \U$2758 ( \3101 , \3074 , \3100 );
xor \U$2759 ( \3102 , \2617 , \2619 );
xor \U$2760 ( \3103 , \3102 , \2622 );
and \U$2761 ( \3104 , \3101 , \3103 );
and \U$2762 ( \3105 , \3074 , \3100 );
or \U$2763 ( \3106 , \3104 , \3105 );
not \U$2764 ( \3107 , \2184 );
not \U$2765 ( \3108 , \2404 );
or \U$2766 ( \3109 , \3107 , \3108 );
or \U$2767 ( \3110 , \2404 , \2184 );
nand \U$2768 ( \3111 , \3109 , \3110 );
xor \U$2769 ( \3112 , \3106 , \3111 );
not \U$2770 ( \3113 , \2612 );
xor \U$2771 ( \3114 , \2609 , \2625 );
not \U$2772 ( \3115 , \3114 );
or \U$2773 ( \3116 , \3113 , \3115 );
or \U$2774 ( \3117 , \3114 , \2612 );
nand \U$2775 ( \3118 , \3116 , \3117 );
and \U$2776 ( \3119 , \3112 , \3118 );
and \U$2777 ( \3120 , \3106 , \3111 );
or \U$2778 ( \3121 , \3119 , \3120 );
nand \U$2779 ( \3122 , \2926 , \3121 );
nand \U$2780 ( \3123 , \2923 , \3122 );
and \U$2781 ( \3124 , \2917 , \3123 );
xor \U$2782 ( \3125 , \3123 , \2917 );
xor \U$2783 ( \3126 , \3106 , \3111 );
xor \U$2784 ( \3127 , \3126 , \3118 );
not \U$2785 ( \3128 , \3127 );
not \U$2786 ( \3129 , \3097 );
xor \U$2787 ( \3130 , \3083 , \3093 );
not \U$2788 ( \3131 , \3130 );
and \U$2789 ( \3132 , \3129 , \3131 );
and \U$2790 ( \3133 , \3097 , \3130 );
nor \U$2791 ( \3134 , \3132 , \3133 );
not \U$2792 ( \3135 , \2528 );
not \U$2793 ( \3136 , \2498 );
or \U$2794 ( \3137 , \3135 , \3136 );
or \U$2795 ( \3138 , \2498 , \2528 );
nand \U$2796 ( \3139 , \3137 , \3138 );
not \U$2797 ( \3140 , \3139 );
not \U$2798 ( \3141 , \2472 );
and \U$2799 ( \3142 , \3140 , \3141 );
and \U$2800 ( \3143 , \3139 , \2472 );
nor \U$2801 ( \3144 , \3142 , \3143 );
or \U$2802 ( \3145 , \3134 , \3144 );
not \U$2803 ( \3146 , \3144 );
not \U$2804 ( \3147 , \3134 );
or \U$2805 ( \3148 , \3146 , \3147 );
xor \U$2806 ( \3149 , \3002 , \3058 );
xor \U$2807 ( \3150 , \3149 , \3071 );
nand \U$2808 ( \3151 , \3148 , \3150 );
nand \U$2809 ( \3152 , \3145 , \3151 );
not \U$2810 ( \3153 , \2607 );
xor \U$2811 ( \3154 , \2578 , \2530 );
not \U$2812 ( \3155 , \3154 );
or \U$2813 ( \3156 , \3153 , \3155 );
or \U$2814 ( \3157 , \3154 , \2607 );
nand \U$2815 ( \3158 , \3156 , \3157 );
xor \U$2816 ( \3159 , \3152 , \3158 );
xor \U$2817 ( \3160 , \2539 , \2546 );
xor \U$2818 ( \3161 , \3160 , \2575 );
not \U$2819 ( \3162 , \3161 );
not \U$2820 ( \3163 , \3009 );
not \U$2821 ( \3164 , \3022 );
or \U$2822 ( \3165 , \3163 , \3164 );
or \U$2823 ( \3166 , \3009 , \3022 );
nand \U$2824 ( \3167 , \3165 , \3166 );
not \U$2825 ( \3168 , \3167 );
not \U$2826 ( \3169 , \3010 );
and \U$2827 ( \3170 , \3168 , \3169 );
and \U$2828 ( \3171 , \3167 , \3010 );
nor \U$2829 ( \3172 , \3170 , \3171 );
and \U$2830 ( \3173 , \416 , RI986eda0_37);
and \U$2831 ( \3174 , RI986ebc0_33, \414 );
nor \U$2832 ( \3175 , \3173 , \3174 );
and \U$2833 ( \3176 , \3175 , \421 );
not \U$2834 ( \3177 , \3175 );
and \U$2835 ( \3178 , \3177 , \422 );
nor \U$2836 ( \3179 , \3176 , \3178 );
not \U$2837 ( \3180 , \3179 );
nand \U$2838 ( \3181 , RI986ee90_39, RI9871fc8_144);
not \U$2839 ( \3182 , \3181 );
and \U$2840 ( \3183 , \3180 , \3182 );
and \U$2841 ( \3184 , \3179 , \3181 );
and \U$2842 ( \3185 , \354 , RI986ecb0_35);
and \U$2843 ( \3186 , RI986f070_43, \352 );
nor \U$2844 ( \3187 , \3185 , \3186 );
not \U$2845 ( \3188 , \3187 );
not \U$2846 ( \3189 , \361 );
and \U$2847 ( \3190 , \3188 , \3189 );
and \U$2848 ( \3191 , \3187 , \345 );
nor \U$2849 ( \3192 , \3190 , \3191 );
nor \U$2850 ( \3193 , \3184 , \3192 );
nor \U$2851 ( \3194 , \3183 , \3193 );
or \U$2852 ( \3195 , \3172 , \3194 );
not \U$2853 ( \3196 , \3194 );
not \U$2854 ( \3197 , \3172 );
or \U$2855 ( \3198 , \3196 , \3197 );
not \U$2856 ( \3199 , \365 );
and \U$2857 ( \3200 , \376 , RI986f160_45);
and \U$2858 ( \3201 , RI986e530_19, \374 );
nor \U$2859 ( \3202 , \3200 , \3201 );
not \U$2860 ( \3203 , \3202 );
or \U$2861 ( \3204 , \3199 , \3203 );
or \U$2862 ( \3205 , \3202 , \367 );
nand \U$2863 ( \3206 , \3204 , \3205 );
not \U$2864 ( \3207 , \456 );
and \U$2865 ( \3208 , \465 , RI986e440_17);
and \U$2866 ( \3209 , RI986e710_23, \463 );
nor \U$2867 ( \3210 , \3208 , \3209 );
not \U$2868 ( \3211 , \3210 );
or \U$2869 ( \3212 , \3207 , \3211 );
or \U$2870 ( \3213 , \3210 , \454 );
nand \U$2871 ( \3214 , \3212 , \3213 );
xor \U$2872 ( \3215 , \3206 , \3214 );
not \U$2873 ( \3216 , \487 );
and \U$2874 ( \3217 , \395 , RI986ef80_41);
and \U$2875 ( \3218 , RI986f250_47, \393 );
nor \U$2876 ( \3219 , \3217 , \3218 );
not \U$2877 ( \3220 , \3219 );
or \U$2878 ( \3221 , \3216 , \3220 );
or \U$2879 ( \3222 , \3219 , \386 );
nand \U$2880 ( \3223 , \3221 , \3222 );
and \U$2881 ( \3224 , \3215 , \3223 );
and \U$2882 ( \3225 , \3206 , \3214 );
or \U$2883 ( \3226 , \3224 , \3225 );
nand \U$2884 ( \3227 , \3198 , \3226 );
nand \U$2885 ( \3228 , \3195 , \3227 );
and \U$2886 ( \3229 , \2274 , RI986dcc0_1);
and \U$2887 ( \3230 , RI986e170_11, \2272 );
nor \U$2888 ( \3231 , \3229 , \3230 );
and \U$2889 ( \3232 , \3231 , \2031 );
not \U$2890 ( \3233 , \3231 );
and \U$2891 ( \3234 , \3233 , \2030 );
nor \U$2892 ( \3235 , \3232 , \3234 );
not \U$2893 ( \3236 , \3235 );
and \U$2894 ( \3237 , \2464 , RI986e080_9);
and \U$2895 ( \3238 , RI986e260_13, \2462 );
nor \U$2896 ( \3239 , \3237 , \3238 );
and \U$2897 ( \3240 , \3239 , \2263 );
not \U$2898 ( \3241 , \3239 );
and \U$2899 ( \3242 , \3241 , \2468 );
nor \U$2900 ( \3243 , \3240 , \3242 );
not \U$2901 ( \3244 , \3243 );
and \U$2902 ( \3245 , \3236 , \3244 );
and \U$2903 ( \3246 , \3243 , \3235 );
and \U$2904 ( \3247 , RI98725e0_157, RI98727c0_161);
not \U$2905 ( \3248 , RI98727c0_161);
nor \U$2906 ( \3249 , \3248 , RI9872388_152);
not \U$2907 ( \3250 , RI9872388_152);
nor \U$2908 ( \3251 , \3250 , RI98727c0_161);
or \U$2909 ( \3252 , \3249 , \3251 );
nor \U$2910 ( \3253 , RI98725e0_157, RI98727c0_161);
nor \U$2911 ( \3254 , \3247 , \3252 , \3253 );
nand \U$2912 ( \3255 , RI986e350_15, \3254 );
not \U$2913 ( \3256 , \3255 );
not \U$2914 ( \3257 , \2935 );
and \U$2915 ( \3258 , \3256 , \3257 );
and \U$2916 ( \3259 , \3255 , \2935 );
nor \U$2917 ( \3260 , \3258 , \3259 );
nor \U$2918 ( \3261 , \3246 , \3260 );
nor \U$2919 ( \3262 , \3245 , \3261 );
and \U$2920 ( \3263 , \438 , RI986e620_21);
and \U$2921 ( \3264 , RI986f7f0_59, \436 );
nor \U$2922 ( \3265 , \3263 , \3264 );
and \U$2923 ( \3266 , \3265 , \443 );
not \U$2924 ( \3267 , \3265 );
and \U$2925 ( \3268 , \3267 , \444 );
nor \U$2926 ( \3269 , \3266 , \3268 );
not \U$2927 ( \3270 , \3269 );
and \U$2928 ( \3271 , \1293 , RI986f8e0_61);
and \U$2929 ( \3272 , RI986f430_51, \1291 );
nor \U$2930 ( \3273 , \3271 , \3272 );
not \U$2931 ( \3274 , \3273 );
not \U$2932 ( \3275 , \1301 );
and \U$2933 ( \3276 , \3274 , \3275 );
and \U$2934 ( \3277 , \3273 , \1301 );
nor \U$2935 ( \3278 , \3276 , \3277 );
not \U$2936 ( \3279 , \3278 );
and \U$2937 ( \3280 , \3270 , \3279 );
and \U$2938 ( \3281 , \3278 , \3269 );
and \U$2939 ( \3282 , \776 , RI986f700_57);
and \U$2940 ( \3283 , RI986f9d0_63, \774 );
nor \U$2941 ( \3284 , \3282 , \3283 );
and \U$2942 ( \3285 , \3284 , \451 );
not \U$2943 ( \3286 , \3284 );
and \U$2944 ( \3287 , \3286 , \474 );
nor \U$2945 ( \3288 , \3285 , \3287 );
nor \U$2946 ( \3289 , \3281 , \3288 );
nor \U$2947 ( \3290 , \3280 , \3289 );
or \U$2948 ( \3291 , \3262 , \3290 );
not \U$2949 ( \3292 , \3262 );
not \U$2950 ( \3293 , \3290 );
or \U$2951 ( \3294 , \3292 , \3293 );
and \U$2952 ( \3295 , \1311 , RI986f610_55);
and \U$2953 ( \3296 , RI986df90_7, \1309 );
nor \U$2954 ( \3297 , \3295 , \3296 );
and \U$2955 ( \3298 , \3297 , \1458 );
not \U$2956 ( \3299 , \3297 );
and \U$2957 ( \3300 , \3299 , \1318 );
nor \U$2958 ( \3301 , \3298 , \3300 );
and \U$2959 ( \3302 , \1329 , RI986f340_49);
and \U$2960 ( \3303 , RI986f520_53, \1327 );
nor \U$2961 ( \3304 , \3302 , \3303 );
and \U$2962 ( \3305 , \3304 , \1336 );
not \U$2963 ( \3306 , \3304 );
and \U$2964 ( \3307 , \3306 , \1337 );
nor \U$2965 ( \3308 , \3305 , \3307 );
xor \U$2966 ( \3309 , \3301 , \3308 );
not \U$2967 ( \3310 , \1462 );
and \U$2968 ( \3311 , \2042 , RI986dea0_5);
and \U$2969 ( \3312 , RI986ddb0_3, \2040 );
nor \U$2970 ( \3313 , \3311 , \3312 );
not \U$2971 ( \3314 , \3313 );
or \U$2972 ( \3315 , \3310 , \3314 );
or \U$2973 ( \3316 , \3313 , \2034 );
nand \U$2974 ( \3317 , \3315 , \3316 );
and \U$2975 ( \3318 , \3309 , \3317 );
and \U$2976 ( \3319 , \3301 , \3308 );
or \U$2977 ( \3320 , \3318 , \3319 );
nand \U$2978 ( \3321 , \3294 , \3320 );
nand \U$2979 ( \3322 , \3291 , \3321 );
xor \U$2980 ( \3323 , \3228 , \3322 );
xor \U$2981 ( \3324 , \3035 , \3043 );
xor \U$2982 ( \3325 , \3324 , \3052 );
xor \U$2983 ( \3326 , \2954 , \2961 );
xor \U$2984 ( \3327 , \3326 , \2969 );
xor \U$2985 ( \3328 , \3325 , \3327 );
xor \U$2986 ( \3329 , \2981 , \2988 );
xor \U$2987 ( \3330 , \3329 , \2996 );
and \U$2988 ( \3331 , \3328 , \3330 );
and \U$2989 ( \3332 , \3325 , \3327 );
nor \U$2990 ( \3333 , \3331 , \3332 );
and \U$2991 ( \3334 , \3323 , \3333 );
and \U$2992 ( \3335 , \3228 , \3322 );
or \U$2993 ( \3336 , \3334 , \3335 );
not \U$2994 ( \3337 , \3336 );
or \U$2995 ( \3338 , \3162 , \3337 );
or \U$2996 ( \3339 , \3336 , \3161 );
not \U$2997 ( \3340 , \2446 );
xor \U$2998 ( \3341 , \2470 , \2454 );
not \U$2999 ( \3342 , \3341 );
or \U$3000 ( \3343 , \3340 , \3342 );
or \U$3001 ( \3344 , \3341 , \2446 );
nand \U$3002 ( \3345 , \3343 , \3344 );
xor \U$3003 ( \3346 , \3024 , \3026 );
xor \U$3004 ( \3347 , \3346 , \3055 );
and \U$3005 ( \3348 , \3345 , \3347 );
xor \U$3006 ( \3349 , \2510 , \2517 );
xor \U$3007 ( \3350 , \3349 , \2525 );
xor \U$3008 ( \3351 , \3061 , \3066 );
xor \U$3009 ( \3352 , \3350 , \3351 );
xor \U$3010 ( \3353 , \3024 , \3026 );
xor \U$3011 ( \3354 , \3353 , \3055 );
and \U$3012 ( \3355 , \3352 , \3354 );
and \U$3013 ( \3356 , \3345 , \3352 );
or \U$3014 ( \3357 , \3348 , \3355 , \3356 );
nand \U$3015 ( \3358 , \3339 , \3357 );
nand \U$3016 ( \3359 , \3338 , \3358 );
xor \U$3017 ( \3360 , \3159 , \3359 );
xor \U$3018 ( \3361 , \3074 , \3100 );
xor \U$3019 ( \3362 , \3361 , \3103 );
and \U$3020 ( \3363 , \3360 , \3362 );
not \U$3021 ( \3364 , \3360 );
not \U$3022 ( \3365 , \3362 );
and \U$3023 ( \3366 , \3364 , \3365 );
xnor \U$3024 ( \3367 , \3357 , \3336 );
not \U$3025 ( \3368 , \3367 );
not \U$3026 ( \3369 , \3161 );
and \U$3027 ( \3370 , \3368 , \3369 );
and \U$3028 ( \3371 , \3367 , \3161 );
nor \U$3029 ( \3372 , \3370 , \3371 );
and \U$3030 ( \3373 , \1311 , RI986f520_53);
and \U$3031 ( \3374 , RI986f610_55, \1309 );
nor \U$3032 ( \3375 , \3373 , \3374 );
and \U$3033 ( \3376 , \3375 , \1315 );
not \U$3034 ( \3377 , \3375 );
and \U$3035 ( \3378 , \3377 , \1458 );
nor \U$3036 ( \3379 , \3376 , \3378 );
not \U$3037 ( \3380 , \3379 );
and \U$3038 ( \3381 , \2274 , RI986ddb0_3);
and \U$3039 ( \3382 , RI986dcc0_1, \2272 );
nor \U$3040 ( \3383 , \3381 , \3382 );
and \U$3041 ( \3384 , \3383 , \2031 );
not \U$3042 ( \3385 , \3383 );
and \U$3043 ( \3386 , \3385 , \2030 );
nor \U$3044 ( \3387 , \3384 , \3386 );
not \U$3045 ( \3388 , \3387 );
and \U$3046 ( \3389 , \3380 , \3388 );
and \U$3047 ( \3390 , \3387 , \3379 );
and \U$3048 ( \3391 , \2042 , RI986df90_7);
and \U$3049 ( \3392 , RI986dea0_5, \2040 );
nor \U$3050 ( \3393 , \3391 , \3392 );
not \U$3051 ( \3394 , \3393 );
not \U$3052 ( \3395 , \2034 );
and \U$3053 ( \3396 , \3394 , \3395 );
and \U$3054 ( \3397 , \3393 , \1462 );
nor \U$3055 ( \3398 , \3396 , \3397 );
nor \U$3056 ( \3399 , \3390 , \3398 );
nor \U$3057 ( \3400 , \3389 , \3399 );
and \U$3058 ( \3401 , \3254 , RI986e260_13);
and \U$3059 ( \3402 , RI986e350_15, \3252 );
nor \U$3060 ( \3403 , \3401 , \3402 );
not \U$3061 ( \3404 , \3403 );
not \U$3062 ( \3405 , \2935 );
not \U$3063 ( \3406 , \3405 );
not \U$3064 ( \3407 , \3406 );
and \U$3065 ( \3408 , \3404 , \3407 );
and \U$3066 ( \3409 , \3403 , \2935 );
nor \U$3067 ( \3410 , \3408 , \3409 );
nand \U$3068 ( \3411 , RI9872478_154, RI9872400_153);
and \U$3069 ( \3412 , \3411 , RI9872388_152);
xor \U$3070 ( \3413 , \3410 , \3412 );
and \U$3071 ( \3414 , \2464 , RI986e170_11);
and \U$3072 ( \3415 , RI986e080_9, \2462 );
nor \U$3073 ( \3416 , \3414 , \3415 );
and \U$3074 ( \3417 , \3416 , \2263 );
not \U$3075 ( \3418 , \3416 );
and \U$3076 ( \3419 , \3418 , \2468 );
nor \U$3077 ( \3420 , \3417 , \3419 );
and \U$3078 ( \3421 , \3413 , \3420 );
and \U$3079 ( \3422 , \3410 , \3412 );
or \U$3080 ( \3423 , \3421 , \3422 );
xor \U$3081 ( \3424 , \3400 , \3423 );
and \U$3082 ( \3425 , \1293 , RI986f9d0_63);
and \U$3083 ( \3426 , RI986f8e0_61, \1291 );
nor \U$3084 ( \3427 , \3425 , \3426 );
not \U$3085 ( \3428 , \3427 );
not \U$3086 ( \3429 , \1301 );
and \U$3087 ( \3430 , \3428 , \3429 );
and \U$3088 ( \3431 , \3427 , \1128 );
nor \U$3089 ( \3432 , \3430 , \3431 );
and \U$3090 ( \3433 , \776 , RI986f7f0_59);
and \U$3091 ( \3434 , RI986f700_57, \774 );
nor \U$3092 ( \3435 , \3433 , \3434 );
and \U$3093 ( \3436 , \3435 , \451 );
not \U$3094 ( \3437 , \3435 );
and \U$3095 ( \3438 , \3437 , \474 );
nor \U$3096 ( \3439 , \3436 , \3438 );
xor \U$3097 ( \3440 , \3432 , \3439 );
and \U$3098 ( \3441 , \1329 , RI986f430_51);
and \U$3099 ( \3442 , RI986f340_49, \1327 );
nor \U$3100 ( \3443 , \3441 , \3442 );
and \U$3101 ( \3444 , \3443 , \1337 );
not \U$3102 ( \3445 , \3443 );
and \U$3103 ( \3446 , \3445 , \1336 );
nor \U$3104 ( \3447 , \3444 , \3446 );
and \U$3105 ( \3448 , \3440 , \3447 );
and \U$3106 ( \3449 , \3432 , \3439 );
or \U$3107 ( \3450 , \3448 , \3449 );
and \U$3108 ( \3451 , \3424 , \3450 );
and \U$3109 ( \3452 , \3400 , \3423 );
or \U$3110 ( \3453 , \3451 , \3452 );
and \U$3111 ( \3454 , \465 , RI986e530_19);
and \U$3112 ( \3455 , RI986e440_17, \463 );
nor \U$3113 ( \3456 , \3454 , \3455 );
not \U$3114 ( \3457 , \3456 );
not \U$3115 ( \3458 , \454 );
and \U$3116 ( \3459 , \3457 , \3458 );
and \U$3117 ( \3460 , \3456 , \454 );
nor \U$3118 ( \3461 , \3459 , \3460 );
and \U$3119 ( \3462 , \438 , RI986e710_23);
and \U$3120 ( \3463 , RI986e620_21, \436 );
nor \U$3121 ( \3464 , \3462 , \3463 );
and \U$3122 ( \3465 , \3464 , \443 );
not \U$3123 ( \3466 , \3464 );
and \U$3124 ( \3467 , \3466 , \444 );
nor \U$3125 ( \3468 , \3465 , \3467 );
xor \U$3126 ( \3469 , \3461 , \3468 );
and \U$3127 ( \3470 , \376 , RI986f250_47);
and \U$3128 ( \3471 , RI986f160_45, \374 );
nor \U$3129 ( \3472 , \3470 , \3471 );
not \U$3130 ( \3473 , \3472 );
not \U$3131 ( \3474 , \367 );
and \U$3132 ( \3475 , \3473 , \3474 );
and \U$3133 ( \3476 , \3472 , \367 );
nor \U$3134 ( \3477 , \3475 , \3476 );
and \U$3135 ( \3478 , \3469 , \3477 );
and \U$3136 ( \3479 , \3461 , \3468 );
nor \U$3137 ( \3480 , \3478 , \3479 );
not \U$3138 ( \3481 , \487 );
and \U$3139 ( \3482 , \395 , RI986f070_43);
and \U$3140 ( \3483 , RI986ef80_41, \393 );
nor \U$3141 ( \3484 , \3482 , \3483 );
not \U$3142 ( \3485 , \3484 );
or \U$3143 ( \3486 , \3481 , \3485 );
or \U$3144 ( \3487 , \3484 , \386 );
nand \U$3145 ( \3488 , \3486 , \3487 );
not \U$3146 ( \3489 , \345 );
and \U$3147 ( \3490 , \354 , RI986ebc0_33);
and \U$3148 ( \3491 , RI986ecb0_35, \352 );
nor \U$3149 ( \3492 , \3490 , \3491 );
not \U$3150 ( \3493 , \3492 );
or \U$3151 ( \3494 , \3489 , \3493 );
or \U$3152 ( \3495 , \3492 , \361 );
nand \U$3153 ( \3496 , \3494 , \3495 );
xor \U$3154 ( \3497 , \3488 , \3496 );
and \U$3155 ( \3498 , \416 , RI986ee90_39);
and \U$3156 ( \3499 , RI986eda0_37, \414 );
nor \U$3157 ( \3500 , \3498 , \3499 );
and \U$3158 ( \3501 , \3500 , \422 );
not \U$3159 ( \3502 , \3500 );
and \U$3160 ( \3503 , \3502 , \421 );
nor \U$3161 ( \3504 , \3501 , \3503 );
and \U$3162 ( \3505 , \3497 , \3504 );
and \U$3163 ( \3506 , \3488 , \3496 );
or \U$3164 ( \3507 , \3505 , \3506 );
nor \U$3165 ( \3508 , \3480 , \3507 );
xor \U$3166 ( \3509 , \3453 , \3508 );
not \U$3167 ( \3510 , \3181 );
xor \U$3168 ( \3511 , \3192 , \3179 );
not \U$3169 ( \3512 , \3511 );
or \U$3170 ( \3513 , \3510 , \3512 );
or \U$3171 ( \3514 , \3511 , \3181 );
nand \U$3172 ( \3515 , \3513 , \3514 );
xor \U$3173 ( \3516 , \3206 , \3214 );
xor \U$3174 ( \3517 , \3516 , \3223 );
and \U$3175 ( \3518 , \3515 , \3517 );
not \U$3176 ( \3519 , \3269 );
xor \U$3177 ( \3520 , \3288 , \3278 );
not \U$3178 ( \3521 , \3520 );
or \U$3179 ( \3522 , \3519 , \3521 );
or \U$3180 ( \3523 , \3520 , \3269 );
nand \U$3181 ( \3524 , \3522 , \3523 );
xor \U$3182 ( \3525 , \3206 , \3214 );
xor \U$3183 ( \3526 , \3525 , \3223 );
and \U$3184 ( \3527 , \3524 , \3526 );
and \U$3185 ( \3528 , \3515 , \3524 );
or \U$3186 ( \3529 , \3518 , \3527 , \3528 );
not \U$3187 ( \3530 , \3529 );
and \U$3188 ( \3531 , \3509 , \3530 );
and \U$3189 ( \3532 , \3453 , \3508 );
or \U$3190 ( \3533 , \3531 , \3532 );
not \U$3191 ( \3534 , \3533 );
xor \U$3192 ( \3535 , \2946 , \2972 );
xor \U$3193 ( \3536 , \3535 , \2999 );
not \U$3194 ( \3537 , \3536 );
and \U$3195 ( \3538 , \3534 , \3537 );
and \U$3196 ( \3539 , \3533 , \3536 );
not \U$3197 ( \3540 , \3226 );
not \U$3198 ( \3541 , \3194 );
or \U$3199 ( \3542 , \3540 , \3541 );
or \U$3200 ( \3543 , \3194 , \3226 );
nand \U$3201 ( \3544 , \3542 , \3543 );
not \U$3202 ( \3545 , \3544 );
not \U$3203 ( \3546 , \3172 );
and \U$3204 ( \3547 , \3545 , \3546 );
and \U$3205 ( \3548 , \3544 , \3172 );
nor \U$3206 ( \3549 , \3547 , \3548 );
xor \U$3207 ( \3550 , \2933 , \2935 );
xor \U$3208 ( \3551 , \3550 , \2943 );
xor \U$3209 ( \3552 , \3549 , \3551 );
xor \U$3210 ( \3553 , \3325 , \3327 );
xor \U$3211 ( \3554 , \3553 , \3330 );
and \U$3212 ( \3555 , \3552 , \3554 );
and \U$3213 ( \3556 , \3549 , \3551 );
or \U$3214 ( \3557 , \3555 , \3556 );
nor \U$3215 ( \3558 , \3539 , \3557 );
nor \U$3216 ( \3559 , \3538 , \3558 );
xor \U$3217 ( \3560 , \3372 , \3559 );
not \U$3218 ( \3561 , \3144 );
not \U$3219 ( \3562 , \3150 );
or \U$3220 ( \3563 , \3561 , \3562 );
or \U$3221 ( \3564 , \3150 , \3144 );
nand \U$3222 ( \3565 , \3563 , \3564 );
not \U$3223 ( \3566 , \3565 );
not \U$3224 ( \3567 , \3134 );
and \U$3225 ( \3568 , \3566 , \3567 );
and \U$3226 ( \3569 , \3565 , \3134 );
nor \U$3227 ( \3570 , \3568 , \3569 );
and \U$3228 ( \3571 , \3560 , \3570 );
and \U$3229 ( \3572 , \3372 , \3559 );
or \U$3230 ( \3573 , \3571 , \3572 );
nor \U$3231 ( \3574 , \3366 , \3573 );
nor \U$3232 ( \3575 , \3363 , \3574 );
not \U$3233 ( \3576 , \3575 );
xor \U$3234 ( \3577 , \3152 , \3158 );
and \U$3235 ( \3578 , \3577 , \3359 );
and \U$3236 ( \3579 , \3152 , \3158 );
or \U$3237 ( \3580 , \3578 , \3579 );
not \U$3238 ( \3581 , \3580 );
and \U$3239 ( \3582 , \3576 , \3581 );
and \U$3240 ( \3583 , \3575 , \3580 );
nor \U$3241 ( \3584 , \3582 , \3583 );
not \U$3242 ( \3585 , \3584 );
or \U$3243 ( \3586 , \3128 , \3585 );
or \U$3244 ( \3587 , \3584 , \3127 );
nand \U$3245 ( \3588 , \3586 , \3587 );
not \U$3246 ( \3589 , \3362 );
not \U$3247 ( \3590 , \3573 );
not \U$3248 ( \3591 , \3360 );
and \U$3249 ( \3592 , \3590 , \3591 );
and \U$3250 ( \3593 , \3573 , \3360 );
nor \U$3251 ( \3594 , \3592 , \3593 );
not \U$3252 ( \3595 , \3594 );
or \U$3253 ( \3596 , \3589 , \3595 );
or \U$3254 ( \3597 , \3594 , \3362 );
nand \U$3255 ( \3598 , \3596 , \3597 );
not \U$3256 ( \3599 , \3598 );
xor \U$3257 ( \3600 , \3372 , \3559 );
xor \U$3258 ( \3601 , \3600 , \3570 );
not \U$3259 ( \3602 , \3601 );
xor \U$3260 ( \3603 , \3228 , \3322 );
xor \U$3261 ( \3604 , \3603 , \3333 );
not \U$3262 ( \3605 , \3536 );
xor \U$3263 ( \3606 , \3533 , \3557 );
not \U$3264 ( \3607 , \3606 );
or \U$3265 ( \3608 , \3605 , \3607 );
or \U$3266 ( \3609 , \3606 , \3536 );
nand \U$3267 ( \3610 , \3608 , \3609 );
and \U$3268 ( \3611 , \3604 , \3610 );
and \U$3269 ( \3612 , \3602 , \3611 );
not \U$3270 ( \3613 , \3602 );
not \U$3271 ( \3614 , \3611 );
and \U$3272 ( \3615 , \3613 , \3614 );
not \U$3273 ( \3616 , \3320 );
not \U$3274 ( \3617 , \3262 );
or \U$3275 ( \3618 , \3616 , \3617 );
or \U$3276 ( \3619 , \3262 , \3320 );
nand \U$3277 ( \3620 , \3618 , \3619 );
not \U$3278 ( \3621 , \3620 );
not \U$3279 ( \3622 , \3290 );
and \U$3280 ( \3623 , \3621 , \3622 );
and \U$3281 ( \3624 , \3620 , \3290 );
nor \U$3282 ( \3625 , \3623 , \3624 );
xor \U$3283 ( \3626 , \3453 , \3508 );
xor \U$3284 ( \3627 , \3626 , \3530 );
and \U$3285 ( \3628 , \3625 , \3627 );
xor \U$3286 ( \3629 , \3549 , \3551 );
xor \U$3287 ( \3630 , \3629 , \3554 );
xor \U$3288 ( \3631 , \3453 , \3508 );
xor \U$3289 ( \3632 , \3631 , \3530 );
and \U$3290 ( \3633 , \3630 , \3632 );
and \U$3291 ( \3634 , \3625 , \3630 );
or \U$3292 ( \3635 , \3628 , \3633 , \3634 );
not \U$3293 ( \3636 , \3635 );
xor \U$3294 ( \3637 , \3024 , \3026 );
xor \U$3295 ( \3638 , \3637 , \3055 );
xor \U$3296 ( \3639 , \3345 , \3352 );
xor \U$3297 ( \3640 , \3638 , \3639 );
and \U$3298 ( \3641 , \3636 , \3640 );
and \U$3299 ( \3642 , \2274 , RI986dea0_5);
and \U$3300 ( \3643 , RI986ddb0_3, \2272 );
nor \U$3301 ( \3644 , \3642 , \3643 );
and \U$3302 ( \3645 , \3644 , \2030 );
not \U$3303 ( \3646 , \3644 );
and \U$3304 ( \3647 , \3646 , \2031 );
nor \U$3305 ( \3648 , \3645 , \3647 );
and \U$3306 ( \3649 , \1311 , RI986f340_49);
and \U$3307 ( \3650 , RI986f520_53, \1309 );
nor \U$3308 ( \3651 , \3649 , \3650 );
and \U$3309 ( \3652 , \3651 , \1458 );
not \U$3310 ( \3653 , \3651 );
and \U$3311 ( \3654 , \3653 , \1315 );
nor \U$3312 ( \3655 , \3652 , \3654 );
xor \U$3313 ( \3656 , \3648 , \3655 );
not \U$3314 ( \3657 , \1462 );
and \U$3315 ( \3658 , \2042 , RI986f610_55);
and \U$3316 ( \3659 , RI986df90_7, \2040 );
nor \U$3317 ( \3660 , \3658 , \3659 );
not \U$3318 ( \3661 , \3660 );
or \U$3319 ( \3662 , \3657 , \3661 );
or \U$3320 ( \3663 , \3660 , \1462 );
nand \U$3321 ( \3664 , \3662 , \3663 );
and \U$3322 ( \3665 , \3656 , \3664 );
and \U$3323 ( \3666 , \3648 , \3655 );
or \U$3324 ( \3667 , \3665 , \3666 );
and \U$3325 ( \3668 , \2464 , RI986dcc0_1);
and \U$3326 ( \3669 , RI986e170_11, \2462 );
nor \U$3327 ( \3670 , \3668 , \3669 );
and \U$3328 ( \3671 , \3670 , \2468 );
not \U$3329 ( \3672 , \3670 );
and \U$3330 ( \3673 , \3672 , \2263 );
nor \U$3331 ( \3674 , \3671 , \3673 );
not \U$3332 ( \3675 , \3412 );
and \U$3333 ( \3676 , RI9872388_152, RI9872400_153);
not \U$3334 ( \3677 , RI9872478_154);
and \U$3335 ( \3678 , RI9872400_153, \3677 );
not \U$3336 ( \3679 , RI9872400_153);
and \U$3337 ( \3680 , \3679 , RI9872478_154);
or \U$3338 ( \3681 , \3678 , \3680 );
nor \U$3339 ( \3682 , RI9872388_152, RI9872400_153);
nor \U$3340 ( \3683 , \3676 , \3681 , \3682 );
nand \U$3341 ( \3684 , RI986e350_15, \3683 );
not \U$3342 ( \3685 , \3684 );
or \U$3343 ( \3686 , \3675 , \3685 );
or \U$3344 ( \3687 , \3684 , \3412 );
nand \U$3345 ( \3688 , \3686 , \3687 );
xor \U$3346 ( \3689 , \3674 , \3688 );
not \U$3347 ( \3690 , \3406 );
and \U$3348 ( \3691 , \3254 , RI986e080_9);
and \U$3349 ( \3692 , RI986e260_13, \3252 );
nor \U$3350 ( \3693 , \3691 , \3692 );
not \U$3351 ( \3694 , \3693 );
or \U$3352 ( \3695 , \3690 , \3694 );
or \U$3353 ( \3696 , \3693 , \3406 );
nand \U$3354 ( \3697 , \3695 , \3696 );
and \U$3355 ( \3698 , \3689 , \3697 );
and \U$3356 ( \3699 , \3674 , \3688 );
or \U$3357 ( \3700 , \3698 , \3699 );
xor \U$3358 ( \3701 , \3667 , \3700 );
and \U$3359 ( \3702 , \776 , RI986e620_21);
and \U$3360 ( \3703 , RI986f7f0_59, \774 );
nor \U$3361 ( \3704 , \3702 , \3703 );
and \U$3362 ( \3705 , \3704 , \474 );
not \U$3363 ( \3706 , \3704 );
and \U$3364 ( \3707 , \3706 , \451 );
nor \U$3365 ( \3708 , \3705 , \3707 );
not \U$3366 ( \3709 , \1301 );
and \U$3367 ( \3710 , \1293 , RI986f700_57);
and \U$3368 ( \3711 , RI986f9d0_63, \1291 );
nor \U$3369 ( \3712 , \3710 , \3711 );
not \U$3370 ( \3713 , \3712 );
or \U$3371 ( \3714 , \3709 , \3713 );
or \U$3372 ( \3715 , \3712 , \1301 );
nand \U$3373 ( \3716 , \3714 , \3715 );
xor \U$3374 ( \3717 , \3708 , \3716 );
and \U$3375 ( \3718 , \1329 , RI986f8e0_61);
and \U$3376 ( \3719 , RI986f430_51, \1327 );
nor \U$3377 ( \3720 , \3718 , \3719 );
and \U$3378 ( \3721 , \3720 , \1336 );
not \U$3379 ( \3722 , \3720 );
and \U$3380 ( \3723 , \3722 , \1337 );
nor \U$3381 ( \3724 , \3721 , \3723 );
and \U$3382 ( \3725 , \3717 , \3724 );
and \U$3383 ( \3726 , \3708 , \3716 );
or \U$3384 ( \3727 , \3725 , \3726 );
and \U$3385 ( \3728 , \3701 , \3727 );
and \U$3386 ( \3729 , \3667 , \3700 );
or \U$3387 ( \3730 , \3728 , \3729 );
not \U$3388 ( \3731 , \361 );
and \U$3389 ( \3732 , \354 , RI986eda0_37);
and \U$3390 ( \3733 , RI986ebc0_33, \352 );
nor \U$3391 ( \3734 , \3732 , \3733 );
not \U$3392 ( \3735 , \3734 );
or \U$3393 ( \3736 , \3731 , \3735 );
or \U$3394 ( \3737 , \3734 , \361 );
nand \U$3395 ( \3738 , \3736 , \3737 );
not \U$3396 ( \3739 , \386 );
and \U$3397 ( \3740 , \395 , RI986ecb0_35);
and \U$3398 ( \3741 , RI986f070_43, \393 );
nor \U$3399 ( \3742 , \3740 , \3741 );
not \U$3400 ( \3743 , \3742 );
or \U$3401 ( \3744 , \3739 , \3743 );
or \U$3402 ( \3745 , \3742 , \487 );
nand \U$3403 ( \3746 , \3744 , \3745 );
xor \U$3404 ( \3747 , \3738 , \3746 );
and \U$3405 ( \3748 , \416 , RI986e800_25);
and \U$3406 ( \3749 , RI986ee90_39, \414 );
nor \U$3407 ( \3750 , \3748 , \3749 );
and \U$3408 ( \3751 , \3750 , \422 );
not \U$3409 ( \3752 , \3750 );
and \U$3410 ( \3753 , \3752 , \421 );
nor \U$3411 ( \3754 , \3751 , \3753 );
and \U$3412 ( \3755 , \3747 , \3754 );
and \U$3413 ( \3756 , \3738 , \3746 );
or \U$3414 ( \3757 , \3755 , \3756 );
nand \U$3415 ( \3758 , RI986e8f0_27, RI9871fc8_144);
not \U$3416 ( \3759 , \3758 );
xor \U$3417 ( \3760 , \3757 , \3759 );
not \U$3418 ( \3761 , \367 );
and \U$3419 ( \3762 , \376 , RI986ef80_41);
and \U$3420 ( \3763 , RI986f250_47, \374 );
nor \U$3421 ( \3764 , \3762 , \3763 );
not \U$3422 ( \3765 , \3764 );
or \U$3423 ( \3766 , \3761 , \3765 );
or \U$3424 ( \3767 , \3764 , \365 );
nand \U$3425 ( \3768 , \3766 , \3767 );
and \U$3426 ( \3769 , \438 , RI986e440_17);
and \U$3427 ( \3770 , RI986e710_23, \436 );
nor \U$3428 ( \3771 , \3769 , \3770 );
and \U$3429 ( \3772 , \3771 , \444 );
not \U$3430 ( \3773 , \3771 );
and \U$3431 ( \3774 , \3773 , \443 );
nor \U$3432 ( \3775 , \3772 , \3774 );
xor \U$3433 ( \3776 , \3768 , \3775 );
not \U$3434 ( \3777 , \456 );
and \U$3435 ( \3778 , \465 , RI986f160_45);
and \U$3436 ( \3779 , RI986e530_19, \463 );
nor \U$3437 ( \3780 , \3778 , \3779 );
not \U$3438 ( \3781 , \3780 );
or \U$3439 ( \3782 , \3777 , \3781 );
or \U$3440 ( \3783 , \3780 , \454 );
nand \U$3441 ( \3784 , \3782 , \3783 );
and \U$3442 ( \3785 , \3776 , \3784 );
and \U$3443 ( \3786 , \3768 , \3775 );
or \U$3444 ( \3787 , \3785 , \3786 );
and \U$3445 ( \3788 , \3760 , \3787 );
and \U$3446 ( \3789 , \3757 , \3759 );
or \U$3447 ( \3790 , \3788 , \3789 );
xor \U$3448 ( \3791 , \3730 , \3790 );
xor \U$3449 ( \3792 , \3461 , \3468 );
xor \U$3450 ( \3793 , \3792 , \3477 );
nand \U$3451 ( \3794 , RI986e800_25, RI9871fc8_144);
or \U$3452 ( \3795 , \3793 , \3794 );
not \U$3453 ( \3796 , \3794 );
not \U$3454 ( \3797 , \3793 );
or \U$3455 ( \3798 , \3796 , \3797 );
xor \U$3456 ( \3799 , \3488 , \3496 );
xor \U$3457 ( \3800 , \3799 , \3504 );
nand \U$3458 ( \3801 , \3798 , \3800 );
nand \U$3459 ( \3802 , \3795 , \3801 );
and \U$3460 ( \3803 , \3791 , \3802 );
and \U$3461 ( \3804 , \3730 , \3790 );
or \U$3462 ( \3805 , \3803 , \3804 );
not \U$3463 ( \3806 , \3235 );
xor \U$3464 ( \3807 , \3260 , \3243 );
not \U$3465 ( \3808 , \3807 );
or \U$3466 ( \3809 , \3806 , \3808 );
or \U$3467 ( \3810 , \3807 , \3235 );
nand \U$3468 ( \3811 , \3809 , \3810 );
xor \U$3469 ( \3812 , \3301 , \3308 );
xor \U$3470 ( \3813 , \3812 , \3317 );
and \U$3471 ( \3814 , \3811 , \3813 );
xor \U$3472 ( \3815 , \3410 , \3412 );
xor \U$3473 ( \3816 , \3815 , \3420 );
xor \U$3474 ( \3817 , \3432 , \3439 );
xor \U$3475 ( \3818 , \3817 , \3447 );
or \U$3476 ( \3819 , \3816 , \3818 );
not \U$3477 ( \3820 , \3818 );
not \U$3478 ( \3821 , \3816 );
or \U$3479 ( \3822 , \3820 , \3821 );
not \U$3480 ( \3823 , \3379 );
xor \U$3481 ( \3824 , \3398 , \3387 );
not \U$3482 ( \3825 , \3824 );
or \U$3483 ( \3826 , \3823 , \3825 );
or \U$3484 ( \3827 , \3824 , \3379 );
nand \U$3485 ( \3828 , \3826 , \3827 );
nand \U$3486 ( \3829 , \3822 , \3828 );
nand \U$3487 ( \3830 , \3819 , \3829 );
xor \U$3488 ( \3831 , \3301 , \3308 );
xor \U$3489 ( \3832 , \3831 , \3317 );
and \U$3490 ( \3833 , \3830 , \3832 );
and \U$3491 ( \3834 , \3811 , \3830 );
or \U$3492 ( \3835 , \3814 , \3833 , \3834 );
xor \U$3493 ( \3836 , \3805 , \3835 );
xor \U$3494 ( \3837 , \3400 , \3423 );
xor \U$3495 ( \3838 , \3837 , \3450 );
and \U$3496 ( \3839 , \3480 , \3507 );
nor \U$3497 ( \3840 , \3839 , \3508 );
or \U$3498 ( \3841 , \3838 , \3840 );
not \U$3499 ( \3842 , \3840 );
not \U$3500 ( \3843 , \3838 );
or \U$3501 ( \3844 , \3842 , \3843 );
xor \U$3502 ( \3845 , \3206 , \3214 );
xor \U$3503 ( \3846 , \3845 , \3223 );
xor \U$3504 ( \3847 , \3515 , \3524 );
xor \U$3505 ( \3848 , \3846 , \3847 );
nand \U$3506 ( \3849 , \3844 , \3848 );
nand \U$3507 ( \3850 , \3841 , \3849 );
and \U$3508 ( \3851 , \3836 , \3850 );
and \U$3509 ( \3852 , \3805 , \3835 );
or \U$3510 ( \3853 , \3851 , \3852 );
not \U$3511 ( \3854 , \3640 );
nand \U$3512 ( \3855 , \3854 , \3635 );
and \U$3513 ( \3856 , \3853 , \3855 );
nor \U$3514 ( \3857 , \3641 , \3856 );
nor \U$3515 ( \3858 , \3615 , \3857 );
nor \U$3516 ( \3859 , \3612 , \3858 );
nor \U$3517 ( \3860 , \3599 , \3859 );
and \U$3518 ( \3861 , \3588 , \3860 );
xor \U$3519 ( \3862 , \3860 , \3588 );
not \U$3520 ( \3863 , \3640 );
not \U$3521 ( \3864 , \3635 );
not \U$3522 ( \3865 , \3853 );
and \U$3523 ( \3866 , \3864 , \3865 );
and \U$3524 ( \3867 , \3635 , \3853 );
nor \U$3525 ( \3868 , \3866 , \3867 );
not \U$3526 ( \3869 , \3868 );
or \U$3527 ( \3870 , \3863 , \3869 );
or \U$3528 ( \3871 , \3868 , \3640 );
nand \U$3529 ( \3872 , \3870 , \3871 );
xor \U$3530 ( \3873 , \3604 , \3610 );
and \U$3531 ( \3874 , \3872 , \3873 );
not \U$3532 ( \3875 , \3872 );
not \U$3533 ( \3876 , \3873 );
and \U$3534 ( \3877 , \3875 , \3876 );
xor \U$3535 ( \3878 , \3453 , \3508 );
xor \U$3536 ( \3879 , \3878 , \3530 );
xor \U$3537 ( \3880 , \3625 , \3630 );
xor \U$3538 ( \3881 , \3879 , \3880 );
not \U$3539 ( \3882 , \3881 );
and \U$3540 ( \3883 , \1293 , RI986f7f0_59);
and \U$3541 ( \3884 , RI986f700_57, \1291 );
nor \U$3542 ( \3885 , \3883 , \3884 );
not \U$3543 ( \3886 , \3885 );
not \U$3544 ( \3887 , \1128 );
and \U$3545 ( \3888 , \3886 , \3887 );
and \U$3546 ( \3889 , \3885 , \1128 );
nor \U$3547 ( \3890 , \3888 , \3889 );
and \U$3548 ( \3891 , \1329 , RI986f9d0_63);
and \U$3549 ( \3892 , RI986f8e0_61, \1327 );
nor \U$3550 ( \3893 , \3891 , \3892 );
and \U$3551 ( \3894 , \3893 , \1337 );
not \U$3552 ( \3895 , \3893 );
and \U$3553 ( \3896 , \3895 , \1336 );
nor \U$3554 ( \3897 , \3894 , \3896 );
or \U$3555 ( \3898 , \3890 , \3897 );
not \U$3556 ( \3899 , \3897 );
not \U$3557 ( \3900 , \3890 );
or \U$3558 ( \3901 , \3899 , \3900 );
and \U$3559 ( \3902 , \1311 , RI986f430_51);
and \U$3560 ( \3903 , RI986f340_49, \1309 );
nor \U$3561 ( \3904 , \3902 , \3903 );
and \U$3562 ( \3905 , \3904 , \1458 );
not \U$3563 ( \3906 , \3904 );
and \U$3564 ( \3907 , \3906 , \1315 );
nor \U$3565 ( \3908 , \3905 , \3907 );
nand \U$3566 ( \3909 , \3901 , \3908 );
nand \U$3567 ( \3910 , \3898 , \3909 );
and \U$3568 ( \3911 , \3683 , RI986e260_13);
and \U$3569 ( \3912 , RI986e350_15, \3681 );
nor \U$3570 ( \3913 , \3911 , \3912 );
not \U$3571 ( \3914 , \3913 );
not \U$3572 ( \3915 , \3412 );
and \U$3573 ( \3916 , \3914 , \3915 );
not \U$3574 ( \3917 , \3412 );
not \U$3575 ( \3918 , \3917 );
and \U$3576 ( \3919 , \3913 , \3918 );
nor \U$3577 ( \3920 , \3916 , \3919 );
and \U$3578 ( \3921 , RI98724f0_155, RI9872568_156);
nor \U$3579 ( \3922 , \3921 , \3677 );
buf \U$3580 ( \3923 , \3922 );
or \U$3581 ( \3924 , \3920 , \3923 );
and \U$3582 ( \3925 , \3920 , \3922 );
and \U$3583 ( \3926 , \3254 , RI986e170_11);
and \U$3584 ( \3927 , RI986e080_9, \3252 );
nor \U$3585 ( \3928 , \3926 , \3927 );
not \U$3586 ( \3929 , \3928 );
not \U$3587 ( \3930 , \3406 );
and \U$3588 ( \3931 , \3929 , \3930 );
and \U$3589 ( \3932 , \3928 , \2935 );
nor \U$3590 ( \3933 , \3931 , \3932 );
nor \U$3591 ( \3934 , \3925 , \3933 );
not \U$3592 ( \3935 , \3934 );
nand \U$3593 ( \3936 , \3924 , \3935 );
xor \U$3594 ( \3937 , \3910 , \3936 );
and \U$3595 ( \3938 , \2042 , RI986f520_53);
and \U$3596 ( \3939 , RI986f610_55, \2040 );
nor \U$3597 ( \3940 , \3938 , \3939 );
not \U$3598 ( \3941 , \3940 );
not \U$3599 ( \3942 , \1462 );
and \U$3600 ( \3943 , \3941 , \3942 );
and \U$3601 ( \3944 , \3940 , \1462 );
nor \U$3602 ( \3945 , \3943 , \3944 );
and \U$3603 ( \3946 , \2274 , RI986df90_7);
and \U$3604 ( \3947 , RI986dea0_5, \2272 );
nor \U$3605 ( \3948 , \3946 , \3947 );
and \U$3606 ( \3949 , \3948 , \2031 );
not \U$3607 ( \3950 , \3948 );
and \U$3608 ( \3951 , \3950 , \2030 );
nor \U$3609 ( \3952 , \3949 , \3951 );
or \U$3610 ( \3953 , \3945 , \3952 );
not \U$3611 ( \3954 , \3952 );
not \U$3612 ( \3955 , \3945 );
or \U$3613 ( \3956 , \3954 , \3955 );
and \U$3614 ( \3957 , \2464 , RI986ddb0_3);
and \U$3615 ( \3958 , RI986dcc0_1, \2462 );
nor \U$3616 ( \3959 , \3957 , \3958 );
and \U$3617 ( \3960 , \3959 , \2468 );
not \U$3618 ( \3961 , \3959 );
and \U$3619 ( \3962 , \3961 , \2263 );
nor \U$3620 ( \3963 , \3960 , \3962 );
nand \U$3621 ( \3964 , \3956 , \3963 );
nand \U$3622 ( \3965 , \3953 , \3964 );
and \U$3623 ( \3966 , \3937 , \3965 );
and \U$3624 ( \3967 , \3910 , \3936 );
or \U$3625 ( \3968 , \3966 , \3967 );
not \U$3626 ( \3969 , \487 );
and \U$3627 ( \3970 , \395 , RI986ebc0_33);
and \U$3628 ( \3971 , RI986ecb0_35, \393 );
nor \U$3629 ( \3972 , \3970 , \3971 );
not \U$3630 ( \3973 , \3972 );
or \U$3631 ( \3974 , \3969 , \3973 );
or \U$3632 ( \3975 , \3972 , \487 );
nand \U$3633 ( \3976 , \3974 , \3975 );
not \U$3634 ( \3977 , \367 );
and \U$3635 ( \3978 , \376 , RI986f070_43);
and \U$3636 ( \3979 , RI986ef80_41, \374 );
nor \U$3637 ( \3980 , \3978 , \3979 );
not \U$3638 ( \3981 , \3980 );
or \U$3639 ( \3982 , \3977 , \3981 );
or \U$3640 ( \3983 , \3980 , \367 );
nand \U$3641 ( \3984 , \3982 , \3983 );
xor \U$3642 ( \3985 , \3976 , \3984 );
not \U$3643 ( \3986 , \345 );
and \U$3644 ( \3987 , \354 , RI986ee90_39);
and \U$3645 ( \3988 , RI986eda0_37, \352 );
nor \U$3646 ( \3989 , \3987 , \3988 );
not \U$3647 ( \3990 , \3989 );
or \U$3648 ( \3991 , \3986 , \3990 );
or \U$3649 ( \3992 , \3989 , \345 );
nand \U$3650 ( \3993 , \3991 , \3992 );
and \U$3651 ( \3994 , \3985 , \3993 );
and \U$3652 ( \3995 , \3976 , \3984 );
or \U$3653 ( \3996 , \3994 , \3995 );
not \U$3654 ( \3997 , RI986e9e0_29);
nor \U$3655 ( \3998 , \3997 , \407 );
and \U$3656 ( \3999 , \416 , RI986e8f0_27);
and \U$3657 ( \4000 , RI986e800_25, \414 );
nor \U$3658 ( \4001 , \3999 , \4000 );
and \U$3659 ( \4002 , \4001 , \422 );
not \U$3660 ( \4003 , \4001 );
and \U$3661 ( \4004 , \4003 , \421 );
nor \U$3662 ( \4005 , \4002 , \4004 );
and \U$3663 ( \4006 , \3998 , \4005 );
xor \U$3664 ( \4007 , \3996 , \4006 );
and \U$3665 ( \4008 , \776 , RI986e710_23);
and \U$3666 ( \4009 , RI986e620_21, \774 );
nor \U$3667 ( \4010 , \4008 , \4009 );
and \U$3668 ( \4011 , \4010 , \474 );
not \U$3669 ( \4012 , \4010 );
and \U$3670 ( \4013 , \4012 , \451 );
nor \U$3671 ( \4014 , \4011 , \4013 );
and \U$3672 ( \4015 , \438 , RI986e530_19);
and \U$3673 ( \4016 , RI986e440_17, \436 );
nor \U$3674 ( \4017 , \4015 , \4016 );
and \U$3675 ( \4018 , \4017 , \444 );
not \U$3676 ( \4019 , \4017 );
and \U$3677 ( \4020 , \4019 , \443 );
nor \U$3678 ( \4021 , \4018 , \4020 );
xor \U$3679 ( \4022 , \4014 , \4021 );
not \U$3680 ( \4023 , \456 );
and \U$3681 ( \4024 , \465 , RI986f250_47);
and \U$3682 ( \4025 , RI986f160_45, \463 );
nor \U$3683 ( \4026 , \4024 , \4025 );
not \U$3684 ( \4027 , \4026 );
or \U$3685 ( \4028 , \4023 , \4027 );
or \U$3686 ( \4029 , \4026 , \454 );
nand \U$3687 ( \4030 , \4028 , \4029 );
and \U$3688 ( \4031 , \4022 , \4030 );
and \U$3689 ( \4032 , \4014 , \4021 );
or \U$3690 ( \4033 , \4031 , \4032 );
and \U$3691 ( \4034 , \4007 , \4033 );
and \U$3692 ( \4035 , \3996 , \4006 );
or \U$3693 ( \4036 , \4034 , \4035 );
xor \U$3694 ( \4037 , \3968 , \4036 );
xor \U$3695 ( \4038 , \3768 , \3775 );
xor \U$3696 ( \4039 , \4038 , \3784 );
xor \U$3697 ( \4040 , \4039 , \3758 );
xor \U$3698 ( \4041 , \3738 , \3746 );
xor \U$3699 ( \4042 , \4041 , \3754 );
and \U$3700 ( \4043 , \4040 , \4042 );
and \U$3701 ( \4044 , \4039 , \3758 );
or \U$3702 ( \4045 , \4043 , \4044 );
and \U$3703 ( \4046 , \4037 , \4045 );
and \U$3704 ( \4047 , \3968 , \4036 );
or \U$3705 ( \4048 , \4046 , \4047 );
xor \U$3706 ( \4049 , \3667 , \3700 );
xor \U$3707 ( \4050 , \4049 , \3727 );
xor \U$3708 ( \4051 , \3757 , \3759 );
xor \U$3709 ( \4052 , \4051 , \3787 );
and \U$3710 ( \4053 , \4050 , \4052 );
and \U$3711 ( \4054 , \4048 , \4053 );
not \U$3712 ( \4055 , \4048 );
not \U$3713 ( \4056 , \4053 );
and \U$3714 ( \4057 , \4055 , \4056 );
not \U$3715 ( \4058 , \3828 );
not \U$3716 ( \4059 , \3816 );
or \U$3717 ( \4060 , \4058 , \4059 );
or \U$3718 ( \4061 , \3816 , \3828 );
nand \U$3719 ( \4062 , \4060 , \4061 );
not \U$3720 ( \4063 , \4062 );
not \U$3721 ( \4064 , \3818 );
and \U$3722 ( \4065 , \4063 , \4064 );
and \U$3723 ( \4066 , \4062 , \3818 );
nor \U$3724 ( \4067 , \4065 , \4066 );
not \U$3725 ( \4068 , \4067 );
not \U$3726 ( \4069 , \3794 );
not \U$3727 ( \4070 , \3800 );
or \U$3728 ( \4071 , \4069 , \4070 );
or \U$3729 ( \4072 , \3800 , \3794 );
nand \U$3730 ( \4073 , \4071 , \4072 );
not \U$3731 ( \4074 , \4073 );
not \U$3732 ( \4075 , \3793 );
and \U$3733 ( \4076 , \4074 , \4075 );
and \U$3734 ( \4077 , \4073 , \3793 );
nor \U$3735 ( \4078 , \4076 , \4077 );
not \U$3736 ( \4079 , \4078 );
and \U$3737 ( \4080 , \4068 , \4079 );
and \U$3738 ( \4081 , \4067 , \4078 );
xor \U$3739 ( \4082 , \3674 , \3688 );
xor \U$3740 ( \4083 , \4082 , \3697 );
xor \U$3741 ( \4084 , \3708 , \3716 );
xor \U$3742 ( \4085 , \4084 , \3724 );
and \U$3743 ( \4086 , \4083 , \4085 );
xor \U$3744 ( \4087 , \3648 , \3655 );
xor \U$3745 ( \4088 , \4087 , \3664 );
xor \U$3746 ( \4089 , \3708 , \3716 );
xor \U$3747 ( \4090 , \4089 , \3724 );
and \U$3748 ( \4091 , \4088 , \4090 );
and \U$3749 ( \4092 , \4083 , \4088 );
or \U$3750 ( \4093 , \4086 , \4091 , \4092 );
not \U$3751 ( \4094 , \4093 );
nor \U$3752 ( \4095 , \4081 , \4094 );
nor \U$3753 ( \4096 , \4080 , \4095 );
nor \U$3754 ( \4097 , \4057 , \4096 );
nor \U$3755 ( \4098 , \4054 , \4097 );
not \U$3756 ( \4099 , \4098 );
and \U$3757 ( \4100 , \3882 , \4099 );
and \U$3758 ( \4101 , \3881 , \4098 );
xor \U$3759 ( \4102 , \3301 , \3308 );
xor \U$3760 ( \4103 , \4102 , \3317 );
xor \U$3761 ( \4104 , \3811 , \3830 );
xor \U$3762 ( \4105 , \4103 , \4104 );
xor \U$3763 ( \4106 , \3730 , \3790 );
xor \U$3764 ( \4107 , \4106 , \3802 );
and \U$3765 ( \4108 , \4105 , \4107 );
not \U$3766 ( \4109 , \4105 );
not \U$3767 ( \4110 , \4107 );
and \U$3768 ( \4111 , \4109 , \4110 );
not \U$3769 ( \4112 , \3838 );
not \U$3770 ( \4113 , \3848 );
or \U$3771 ( \4114 , \4112 , \4113 );
or \U$3772 ( \4115 , \3848 , \3838 );
nand \U$3773 ( \4116 , \4114 , \4115 );
not \U$3774 ( \4117 , \4116 );
not \U$3775 ( \4118 , \3840 );
and \U$3776 ( \4119 , \4117 , \4118 );
and \U$3777 ( \4120 , \4116 , \3840 );
nor \U$3778 ( \4121 , \4119 , \4120 );
nor \U$3779 ( \4122 , \4111 , \4121 );
nor \U$3780 ( \4123 , \4108 , \4122 );
nor \U$3781 ( \4124 , \4101 , \4123 );
nor \U$3782 ( \4125 , \4100 , \4124 );
nor \U$3783 ( \4126 , \3877 , \4125 );
nor \U$3784 ( \4127 , \3874 , \4126 );
not \U$3785 ( \4128 , \4127 );
not \U$3786 ( \4129 , \3601 );
not \U$3787 ( \4130 , \3611 );
not \U$3788 ( \4131 , \3857 );
or \U$3789 ( \4132 , \4130 , \4131 );
or \U$3790 ( \4133 , \3857 , \3611 );
nand \U$3791 ( \4134 , \4132 , \4133 );
not \U$3792 ( \4135 , \4134 );
or \U$3793 ( \4136 , \4129 , \4135 );
or \U$3794 ( \4137 , \4134 , \3601 );
nand \U$3795 ( \4138 , \4136 , \4137 );
nand \U$3796 ( \4139 , \4128 , \4138 );
not \U$3797 ( \4140 , \3598 );
not \U$3798 ( \4141 , \3859 );
and \U$3799 ( \4142 , \4140 , \4141 );
and \U$3800 ( \4143 , \3598 , \3859 );
nor \U$3801 ( \4144 , \4142 , \4143 );
xor \U$3802 ( \4145 , \4139 , \4144 );
xor \U$3803 ( \4146 , \3805 , \3835 );
xor \U$3804 ( \4147 , \4146 , \3850 );
not \U$3805 ( \4148 , \4147 );
not \U$3806 ( \4149 , \3881 );
xor \U$3807 ( \4150 , \4098 , \4123 );
not \U$3808 ( \4151 , \4150 );
or \U$3809 ( \4152 , \4149 , \4151 );
or \U$3810 ( \4153 , \4150 , \3881 );
nand \U$3811 ( \4154 , \4152 , \4153 );
not \U$3812 ( \4155 , \4154 );
or \U$3813 ( \4156 , \4148 , \4155 );
or \U$3814 ( \4157 , \4154 , \4147 );
xor \U$3815 ( \4158 , \4050 , \4052 );
xor \U$3816 ( \4159 , \3968 , \4036 );
xor \U$3817 ( \4160 , \4159 , \4045 );
and \U$3818 ( \4161 , \4158 , \4160 );
not \U$3819 ( \4162 , \4078 );
not \U$3820 ( \4163 , \4093 );
not \U$3821 ( \4164 , \4067 );
or \U$3822 ( \4165 , \4163 , \4164 );
or \U$3823 ( \4166 , \4067 , \4093 );
nand \U$3824 ( \4167 , \4165 , \4166 );
not \U$3825 ( \4168 , \4167 );
or \U$3826 ( \4169 , \4162 , \4168 );
or \U$3827 ( \4170 , \4167 , \4078 );
nand \U$3828 ( \4171 , \4169 , \4170 );
xor \U$3829 ( \4172 , \3968 , \4036 );
xor \U$3830 ( \4173 , \4172 , \4045 );
and \U$3831 ( \4174 , \4171 , \4173 );
and \U$3832 ( \4175 , \4158 , \4171 );
or \U$3833 ( \4176 , \4161 , \4174 , \4175 );
and \U$3834 ( \4177 , \3254 , RI986dcc0_1);
and \U$3835 ( \4178 , RI986e170_11, \3252 );
nor \U$3836 ( \4179 , \4177 , \4178 );
not \U$3837 ( \4180 , \4179 );
not \U$3838 ( \4181 , \2935 );
and \U$3839 ( \4182 , \4180 , \4181 );
and \U$3840 ( \4183 , \4179 , \3406 );
nor \U$3841 ( \4184 , \4182 , \4183 );
not \U$3842 ( \4185 , \4184 );
and \U$3843 ( \4186 , \3683 , RI986e080_9);
and \U$3844 ( \4187 , RI986e260_13, \3681 );
nor \U$3845 ( \4188 , \4186 , \4187 );
not \U$3846 ( \4189 , \4188 );
not \U$3847 ( \4190 , \3918 );
and \U$3848 ( \4191 , \4189 , \4190 );
and \U$3849 ( \4192 , \4188 , \3412 );
nor \U$3850 ( \4193 , \4191 , \4192 );
not \U$3851 ( \4194 , \4193 );
and \U$3852 ( \4195 , \4185 , \4194 );
and \U$3853 ( \4196 , \4193 , \4184 );
and \U$3854 ( \4197 , RI9872478_154, RI98724f0_155);
not \U$3855 ( \4198 , RI9872568_156);
and \U$3856 ( \4199 , \4198 , RI98724f0_155);
nor \U$3857 ( \4200 , \4198 , RI98724f0_155);
or \U$3858 ( \4201 , \4199 , \4200 );
nor \U$3859 ( \4202 , RI9872478_154, RI98724f0_155);
nor \U$3860 ( \4203 , \4197 , \4201 , \4202 );
nand \U$3861 ( \4204 , RI986e350_15, \4203 );
and \U$3862 ( \4205 , \4204 , \3922 );
not \U$3863 ( \4206 , \4204 );
not \U$3864 ( \4207 , \3922 );
and \U$3865 ( \4208 , \4206 , \4207 );
nor \U$3866 ( \4209 , \4205 , \4208 );
nor \U$3867 ( \4210 , \4196 , \4209 );
nor \U$3868 ( \4211 , \4195 , \4210 );
and \U$3869 ( \4212 , \2042 , RI986f340_49);
and \U$3870 ( \4213 , RI986f520_53, \2040 );
nor \U$3871 ( \4214 , \4212 , \4213 );
not \U$3872 ( \4215 , \4214 );
not \U$3873 ( \4216 , \2034 );
and \U$3874 ( \4217 , \4215 , \4216 );
and \U$3875 ( \4218 , \4214 , \1462 );
nor \U$3876 ( \4219 , \4217 , \4218 );
not \U$3877 ( \4220 , \4219 );
and \U$3878 ( \4221 , \2464 , RI986dea0_5);
and \U$3879 ( \4222 , RI986ddb0_3, \2462 );
nor \U$3880 ( \4223 , \4221 , \4222 );
and \U$3881 ( \4224 , \4223 , \2263 );
not \U$3882 ( \4225 , \4223 );
and \U$3883 ( \4226 , \4225 , \2468 );
nor \U$3884 ( \4227 , \4224 , \4226 );
not \U$3885 ( \4228 , \4227 );
and \U$3886 ( \4229 , \4220 , \4228 );
and \U$3887 ( \4230 , \4227 , \4219 );
and \U$3888 ( \4231 , \2274 , RI986f610_55);
and \U$3889 ( \4232 , RI986df90_7, \2272 );
nor \U$3890 ( \4233 , \4231 , \4232 );
and \U$3891 ( \4234 , \4233 , \2031 );
not \U$3892 ( \4235 , \4233 );
and \U$3893 ( \4236 , \4235 , \2030 );
nor \U$3894 ( \4237 , \4234 , \4236 );
nor \U$3895 ( \4238 , \4230 , \4237 );
nor \U$3896 ( \4239 , \4229 , \4238 );
or \U$3897 ( \4240 , \4211 , \4239 );
not \U$3898 ( \4241 , \4211 );
not \U$3899 ( \4242 , \4239 );
or \U$3900 ( \4243 , \4241 , \4242 );
and \U$3901 ( \4244 , \1311 , RI986f8e0_61);
and \U$3902 ( \4245 , RI986f430_51, \1309 );
nor \U$3903 ( \4246 , \4244 , \4245 );
and \U$3904 ( \4247 , \4246 , \1458 );
not \U$3905 ( \4248 , \4246 );
and \U$3906 ( \4249 , \4248 , \1318 );
nor \U$3907 ( \4250 , \4247 , \4249 );
not \U$3908 ( \4251 , \1128 );
and \U$3909 ( \4252 , \1293 , RI986e620_21);
and \U$3910 ( \4253 , RI986f7f0_59, \1291 );
nor \U$3911 ( \4254 , \4252 , \4253 );
not \U$3912 ( \4255 , \4254 );
or \U$3913 ( \4256 , \4251 , \4255 );
or \U$3914 ( \4257 , \4254 , \1301 );
nand \U$3915 ( \4258 , \4256 , \4257 );
xor \U$3916 ( \4259 , \4250 , \4258 );
and \U$3917 ( \4260 , \1329 , RI986f700_57);
and \U$3918 ( \4261 , RI986f9d0_63, \1327 );
nor \U$3919 ( \4262 , \4260 , \4261 );
and \U$3920 ( \4263 , \4262 , \1336 );
not \U$3921 ( \4264 , \4262 );
and \U$3922 ( \4265 , \4264 , \1337 );
nor \U$3923 ( \4266 , \4263 , \4265 );
and \U$3924 ( \4267 , \4259 , \4266 );
and \U$3925 ( \4268 , \4250 , \4258 );
or \U$3926 ( \4269 , \4267 , \4268 );
nand \U$3927 ( \4270 , \4243 , \4269 );
nand \U$3928 ( \4271 , \4240 , \4270 );
not \U$3929 ( \4272 , \365 );
and \U$3930 ( \4273 , \376 , RI986ecb0_35);
and \U$3931 ( \4274 , RI986f070_43, \374 );
nor \U$3932 ( \4275 , \4273 , \4274 );
not \U$3933 ( \4276 , \4275 );
or \U$3934 ( \4277 , \4272 , \4276 );
or \U$3935 ( \4278 , \4275 , \365 );
nand \U$3936 ( \4279 , \4277 , \4278 );
not \U$3937 ( \4280 , \487 );
and \U$3938 ( \4281 , \395 , RI986eda0_37);
and \U$3939 ( \4282 , RI986ebc0_33, \393 );
nor \U$3940 ( \4283 , \4281 , \4282 );
not \U$3941 ( \4284 , \4283 );
or \U$3942 ( \4285 , \4280 , \4284 );
or \U$3943 ( \4286 , \4283 , \487 );
nand \U$3944 ( \4287 , \4285 , \4286 );
xor \U$3945 ( \4288 , \4279 , \4287 );
not \U$3946 ( \4289 , \361 );
and \U$3947 ( \4290 , \354 , RI986e800_25);
and \U$3948 ( \4291 , RI986ee90_39, \352 );
nor \U$3949 ( \4292 , \4290 , \4291 );
not \U$3950 ( \4293 , \4292 );
or \U$3951 ( \4294 , \4289 , \4293 );
or \U$3952 ( \4295 , \4292 , \361 );
nand \U$3953 ( \4296 , \4294 , \4295 );
and \U$3954 ( \4297 , \4288 , \4296 );
and \U$3955 ( \4298 , \4279 , \4287 );
or \U$3956 ( \4299 , \4297 , \4298 );
nand \U$3957 ( \4300 , RI986ead0_31, RI9871fc8_144);
and \U$3958 ( \4301 , \416 , RI986e9e0_29);
and \U$3959 ( \4302 , RI986e8f0_27, \414 );
nor \U$3960 ( \4303 , \4301 , \4302 );
and \U$3961 ( \4304 , \4303 , \421 );
not \U$3962 ( \4305 , \4303 );
and \U$3963 ( \4306 , \4305 , \422 );
nor \U$3964 ( \4307 , \4304 , \4306 );
nand \U$3965 ( \4308 , \4300 , \4307 );
xor \U$3966 ( \4309 , \4299 , \4308 );
and \U$3967 ( \4310 , \776 , RI986e440_17);
and \U$3968 ( \4311 , RI986e710_23, \774 );
nor \U$3969 ( \4312 , \4310 , \4311 );
and \U$3970 ( \4313 , \4312 , \474 );
not \U$3971 ( \4314 , \4312 );
and \U$3972 ( \4315 , \4314 , \451 );
nor \U$3973 ( \4316 , \4313 , \4315 );
and \U$3974 ( \4317 , \438 , RI986f160_45);
and \U$3975 ( \4318 , RI986e530_19, \436 );
nor \U$3976 ( \4319 , \4317 , \4318 );
and \U$3977 ( \4320 , \4319 , \444 );
not \U$3978 ( \4321 , \4319 );
and \U$3979 ( \4322 , \4321 , \443 );
nor \U$3980 ( \4323 , \4320 , \4322 );
xor \U$3981 ( \4324 , \4316 , \4323 );
not \U$3982 ( \4325 , \454 );
and \U$3983 ( \4326 , \465 , RI986ef80_41);
and \U$3984 ( \4327 , RI986f250_47, \463 );
nor \U$3985 ( \4328 , \4326 , \4327 );
not \U$3986 ( \4329 , \4328 );
or \U$3987 ( \4330 , \4325 , \4329 );
or \U$3988 ( \4331 , \4328 , \456 );
nand \U$3989 ( \4332 , \4330 , \4331 );
and \U$3990 ( \4333 , \4324 , \4332 );
and \U$3991 ( \4334 , \4316 , \4323 );
or \U$3992 ( \4335 , \4333 , \4334 );
and \U$3993 ( \4336 , \4309 , \4335 );
and \U$3994 ( \4337 , \4299 , \4308 );
or \U$3995 ( \4338 , \4336 , \4337 );
xor \U$3996 ( \4339 , \4271 , \4338 );
xor \U$3997 ( \4340 , \3998 , \4005 );
not \U$3998 ( \4341 , \4340 );
xor \U$3999 ( \4342 , \3976 , \3984 );
xor \U$4000 ( \4343 , \4342 , \3993 );
not \U$4001 ( \4344 , \4343 );
or \U$4002 ( \4345 , \4341 , \4344 );
or \U$4003 ( \4346 , \4343 , \4340 );
xor \U$4004 ( \4347 , \4014 , \4021 );
xor \U$4005 ( \4348 , \4347 , \4030 );
nand \U$4006 ( \4349 , \4346 , \4348 );
nand \U$4007 ( \4350 , \4345 , \4349 );
and \U$4008 ( \4351 , \4339 , \4350 );
and \U$4009 ( \4352 , \4271 , \4338 );
or \U$4010 ( \4353 , \4351 , \4352 );
xor \U$4011 ( \4354 , \3910 , \3936 );
xor \U$4012 ( \4355 , \4354 , \3965 );
xor \U$4013 ( \4356 , \3996 , \4006 );
xor \U$4014 ( \4357 , \4356 , \4033 );
and \U$4015 ( \4358 , \4355 , \4357 );
xor \U$4016 ( \4359 , \4353 , \4358 );
and \U$4017 ( \4360 , \3920 , \3922 );
not \U$4018 ( \4361 , \3920 );
and \U$4019 ( \4362 , \4361 , \4207 );
nor \U$4020 ( \4363 , \4360 , \4362 );
not \U$4021 ( \4364 , \4363 );
not \U$4022 ( \4365 , \3933 );
and \U$4023 ( \4366 , \4364 , \4365 );
and \U$4024 ( \4367 , \4363 , \3933 );
nor \U$4025 ( \4368 , \4366 , \4367 );
not \U$4026 ( \4369 , \3897 );
not \U$4027 ( \4370 , \3908 );
or \U$4028 ( \4371 , \4369 , \4370 );
or \U$4029 ( \4372 , \3897 , \3908 );
nand \U$4030 ( \4373 , \4371 , \4372 );
not \U$4031 ( \4374 , \4373 );
not \U$4032 ( \4375 , \3890 );
and \U$4033 ( \4376 , \4374 , \4375 );
and \U$4034 ( \4377 , \4373 , \3890 );
nor \U$4035 ( \4378 , \4376 , \4377 );
xor \U$4036 ( \4379 , \4368 , \4378 );
not \U$4037 ( \4380 , \3952 );
not \U$4038 ( \4381 , \3963 );
or \U$4039 ( \4382 , \4380 , \4381 );
or \U$4040 ( \4383 , \3952 , \3963 );
nand \U$4041 ( \4384 , \4382 , \4383 );
not \U$4042 ( \4385 , \4384 );
not \U$4043 ( \4386 , \3945 );
and \U$4044 ( \4387 , \4385 , \4386 );
and \U$4045 ( \4388 , \4384 , \3945 );
nor \U$4046 ( \4389 , \4387 , \4388 );
and \U$4047 ( \4390 , \4379 , \4389 );
and \U$4048 ( \4391 , \4368 , \4378 );
nor \U$4049 ( \4392 , \4390 , \4391 );
xor \U$4050 ( \4393 , \4039 , \3758 );
xor \U$4051 ( \4394 , \4393 , \4042 );
and \U$4052 ( \4395 , \4392 , \4394 );
xor \U$4053 ( \4396 , \3708 , \3716 );
xor \U$4054 ( \4397 , \4396 , \3724 );
xor \U$4055 ( \4398 , \4083 , \4088 );
xor \U$4056 ( \4399 , \4397 , \4398 );
xor \U$4057 ( \4400 , \4039 , \3758 );
xor \U$4058 ( \4401 , \4400 , \4042 );
and \U$4059 ( \4402 , \4399 , \4401 );
and \U$4060 ( \4403 , \4392 , \4399 );
or \U$4061 ( \4404 , \4395 , \4402 , \4403 );
and \U$4062 ( \4405 , \4359 , \4404 );
and \U$4063 ( \4406 , \4353 , \4358 );
or \U$4064 ( \4407 , \4405 , \4406 );
xor \U$4065 ( \4408 , \4176 , \4407 );
not \U$4066 ( \4409 , \4121 );
xor \U$4067 ( \4410 , \4107 , \4105 );
not \U$4068 ( \4411 , \4410 );
or \U$4069 ( \4412 , \4409 , \4411 );
or \U$4070 ( \4413 , \4410 , \4121 );
nand \U$4071 ( \4414 , \4412 , \4413 );
and \U$4072 ( \4415 , \4408 , \4414 );
and \U$4073 ( \4416 , \4176 , \4407 );
or \U$4074 ( \4417 , \4415 , \4416 );
nand \U$4075 ( \4418 , \4157 , \4417 );
nand \U$4076 ( \4419 , \4156 , \4418 );
not \U$4077 ( \4420 , \3873 );
not \U$4078 ( \4421 , \4125 );
not \U$4079 ( \4422 , \3872 );
and \U$4080 ( \4423 , \4421 , \4422 );
and \U$4081 ( \4424 , \4125 , \3872 );
nor \U$4082 ( \4425 , \4423 , \4424 );
not \U$4083 ( \4426 , \4425 );
or \U$4084 ( \4427 , \4420 , \4426 );
or \U$4085 ( \4428 , \4425 , \3873 );
nand \U$4086 ( \4429 , \4427 , \4428 );
and \U$4087 ( \4430 , \4419 , \4429 );
not \U$4088 ( \4431 , \4127 );
not \U$4089 ( \4432 , \4138 );
or \U$4090 ( \4433 , \4431 , \4432 );
or \U$4091 ( \4434 , \4138 , \4127 );
nand \U$4092 ( \4435 , \4433 , \4434 );
and \U$4093 ( \4436 , \4430 , \4435 );
xor \U$4094 ( \4437 , \4430 , \4435 );
xor \U$4095 ( \4438 , \4299 , \4308 );
xor \U$4096 ( \4439 , \4438 , \4335 );
not \U$4097 ( \4440 , \4439 );
not \U$4098 ( \4441 , \4269 );
not \U$4099 ( \4442 , \4211 );
or \U$4100 ( \4443 , \4441 , \4442 );
or \U$4101 ( \4444 , \4211 , \4269 );
nand \U$4102 ( \4445 , \4443 , \4444 );
not \U$4103 ( \4446 , \4445 );
not \U$4104 ( \4447 , \4239 );
and \U$4105 ( \4448 , \4446 , \4447 );
and \U$4106 ( \4449 , \4445 , \4239 );
nor \U$4107 ( \4450 , \4448 , \4449 );
not \U$4108 ( \4451 , \4450 );
and \U$4109 ( \4452 , \4440 , \4451 );
and \U$4110 ( \4453 , \4439 , \4450 );
nor \U$4111 ( \4454 , \4452 , \4453 );
not \U$4112 ( \4455 , \1462 );
and \U$4113 ( \4456 , \2042 , RI986f430_51);
and \U$4114 ( \4457 , RI986f340_49, \2040 );
nor \U$4115 ( \4458 , \4456 , \4457 );
not \U$4116 ( \4459 , \4458 );
or \U$4117 ( \4460 , \4455 , \4459 );
or \U$4118 ( \4461 , \4458 , \1462 );
nand \U$4119 ( \4462 , \4460 , \4461 );
and \U$4120 ( \4463 , \1329 , RI986f7f0_59);
and \U$4121 ( \4464 , RI986f700_57, \1327 );
nor \U$4122 ( \4465 , \4463 , \4464 );
and \U$4123 ( \4466 , \4465 , \1336 );
not \U$4124 ( \4467 , \4465 );
and \U$4125 ( \4468 , \4467 , \1337 );
nor \U$4126 ( \4469 , \4466 , \4468 );
xor \U$4127 ( \4470 , \4462 , \4469 );
and \U$4128 ( \4471 , \1311 , RI986f9d0_63);
and \U$4129 ( \4472 , RI986f8e0_61, \1309 );
nor \U$4130 ( \4473 , \4471 , \4472 );
and \U$4131 ( \4474 , \4473 , \1458 );
not \U$4132 ( \4475 , \4473 );
and \U$4133 ( \4476 , \4475 , \1318 );
nor \U$4134 ( \4477 , \4474 , \4476 );
and \U$4135 ( \4478 , \4470 , \4477 );
and \U$4136 ( \4479 , \4462 , \4469 );
or \U$4137 ( \4480 , \4478 , \4479 );
not \U$4138 ( \4481 , \2935 );
and \U$4139 ( \4482 , \3254 , RI986ddb0_3);
and \U$4140 ( \4483 , RI986dcc0_1, \3252 );
nor \U$4141 ( \4484 , \4482 , \4483 );
not \U$4142 ( \4485 , \4484 );
or \U$4143 ( \4486 , \4481 , \4485 );
or \U$4144 ( \4487 , \4484 , \2935 );
nand \U$4145 ( \4488 , \4486 , \4487 );
and \U$4146 ( \4489 , \2274 , RI986f520_53);
and \U$4147 ( \4490 , RI986f610_55, \2272 );
nor \U$4148 ( \4491 , \4489 , \4490 );
and \U$4149 ( \4492 , \4491 , \2030 );
not \U$4150 ( \4493 , \4491 );
and \U$4151 ( \4494 , \4493 , \2031 );
nor \U$4152 ( \4495 , \4492 , \4494 );
xor \U$4153 ( \4496 , \4488 , \4495 );
and \U$4154 ( \4497 , \2464 , RI986df90_7);
and \U$4155 ( \4498 , RI986dea0_5, \2462 );
nor \U$4156 ( \4499 , \4497 , \4498 );
and \U$4157 ( \4500 , \4499 , \2468 );
not \U$4158 ( \4501 , \4499 );
and \U$4159 ( \4502 , \4501 , \2263 );
nor \U$4160 ( \4503 , \4500 , \4502 );
and \U$4161 ( \4504 , \4496 , \4503 );
and \U$4162 ( \4505 , \4488 , \4495 );
or \U$4163 ( \4506 , \4504 , \4505 );
and \U$4164 ( \4507 , \4480 , \4506 );
not \U$4165 ( \4508 , \4506 );
not \U$4166 ( \4509 , \4480 );
and \U$4167 ( \4510 , \4508 , \4509 );
and \U$4168 ( \4511 , \4203 , RI986e260_13);
and \U$4169 ( \4512 , RI986e350_15, \4201 );
nor \U$4170 ( \4513 , \4511 , \4512 );
and \U$4171 ( \4514 , \4513 , \3922 );
not \U$4172 ( \4515 , \4513 );
and \U$4173 ( \4516 , \4515 , \4207 );
nor \U$4174 ( \4517 , \4514 , \4516 );
nand \U$4175 ( \4518 , RI98728b0_163, RI9872838_162);
and \U$4176 ( \4519 , \4518 , RI9872568_156);
not \U$4177 ( \4520 , \4519 );
not \U$4178 ( \4521 , \4520 );
xor \U$4179 ( \4522 , \4517 , \4521 );
and \U$4180 ( \4523 , \3683 , RI986e170_11);
and \U$4181 ( \4524 , RI986e080_9, \3681 );
nor \U$4182 ( \4525 , \4523 , \4524 );
not \U$4183 ( \4526 , \4525 );
not \U$4184 ( \4527 , \3412 );
and \U$4185 ( \4528 , \4526 , \4527 );
and \U$4186 ( \4529 , \4525 , \3918 );
nor \U$4187 ( \4530 , \4528 , \4529 );
and \U$4188 ( \4531 , \4522 , \4530 );
and \U$4189 ( \4532 , \4517 , \4521 );
or \U$4190 ( \4533 , \4531 , \4532 );
nor \U$4191 ( \4534 , \4510 , \4533 );
nor \U$4192 ( \4535 , \4507 , \4534 );
and \U$4193 ( \4536 , \395 , RI986ee90_39);
and \U$4194 ( \4537 , RI986eda0_37, \393 );
nor \U$4195 ( \4538 , \4536 , \4537 );
not \U$4196 ( \4539 , \4538 );
not \U$4197 ( \4540 , \487 );
and \U$4198 ( \4541 , \4539 , \4540 );
and \U$4199 ( \4542 , \4538 , \386 );
nor \U$4200 ( \4543 , \4541 , \4542 );
and \U$4201 ( \4544 , \465 , RI986f070_43);
and \U$4202 ( \4545 , RI986ef80_41, \463 );
nor \U$4203 ( \4546 , \4544 , \4545 );
not \U$4204 ( \4547 , \4546 );
not \U$4205 ( \4548 , \456 );
and \U$4206 ( \4549 , \4547 , \4548 );
and \U$4207 ( \4550 , \4546 , \454 );
nor \U$4208 ( \4551 , \4549 , \4550 );
xor \U$4209 ( \4552 , \4543 , \4551 );
and \U$4210 ( \4553 , \376 , RI986ebc0_33);
and \U$4211 ( \4554 , RI986ecb0_35, \374 );
nor \U$4212 ( \4555 , \4553 , \4554 );
not \U$4213 ( \4556 , \4555 );
not \U$4214 ( \4557 , \365 );
and \U$4215 ( \4558 , \4556 , \4557 );
and \U$4216 ( \4559 , \4555 , \365 );
nor \U$4217 ( \4560 , \4558 , \4559 );
and \U$4218 ( \4561 , \4552 , \4560 );
and \U$4219 ( \4562 , \4543 , \4551 );
or \U$4220 ( \4563 , \4561 , \4562 );
and \U$4221 ( \4564 , \416 , RI986ead0_31);
and \U$4222 ( \4565 , RI986e9e0_29, \414 );
nor \U$4223 ( \4566 , \4564 , \4565 );
and \U$4224 ( \4567 , \4566 , \421 );
not \U$4225 ( \4568 , \4566 );
and \U$4226 ( \4569 , \4568 , \422 );
nor \U$4227 ( \4570 , \4567 , \4569 );
nand \U$4228 ( \4571 , RI98715f0_123, RI9871fc8_144);
xor \U$4229 ( \4572 , \4570 , \4571 );
and \U$4230 ( \4573 , \354 , RI986e8f0_27);
and \U$4231 ( \4574 , RI986e800_25, \352 );
nor \U$4232 ( \4575 , \4573 , \4574 );
not \U$4233 ( \4576 , \4575 );
not \U$4234 ( \4577 , \361 );
and \U$4235 ( \4578 , \4576 , \4577 );
and \U$4236 ( \4579 , \4575 , \345 );
nor \U$4237 ( \4580 , \4578 , \4579 );
and \U$4238 ( \4581 , \4572 , \4580 );
and \U$4239 ( \4582 , \4570 , \4571 );
or \U$4240 ( \4583 , \4581 , \4582 );
xor \U$4241 ( \4584 , \4563 , \4583 );
and \U$4242 ( \4585 , \438 , RI986f250_47);
and \U$4243 ( \4586 , RI986f160_45, \436 );
nor \U$4244 ( \4587 , \4585 , \4586 );
and \U$4245 ( \4588 , \4587 , \443 );
not \U$4246 ( \4589 , \4587 );
and \U$4247 ( \4590 , \4589 , \444 );
nor \U$4248 ( \4591 , \4588 , \4590 );
and \U$4249 ( \4592 , \776 , RI986e530_19);
and \U$4250 ( \4593 , RI986e440_17, \774 );
nor \U$4251 ( \4594 , \4592 , \4593 );
and \U$4252 ( \4595 , \4594 , \451 );
not \U$4253 ( \4596 , \4594 );
and \U$4254 ( \4597 , \4596 , \474 );
nor \U$4255 ( \4598 , \4595 , \4597 );
xor \U$4256 ( \4599 , \4591 , \4598 );
and \U$4257 ( \4600 , \1293 , RI986e710_23);
and \U$4258 ( \4601 , RI986e620_21, \1291 );
nor \U$4259 ( \4602 , \4600 , \4601 );
not \U$4260 ( \4603 , \4602 );
not \U$4261 ( \4604 , \1128 );
and \U$4262 ( \4605 , \4603 , \4604 );
and \U$4263 ( \4606 , \4602 , \1128 );
nor \U$4264 ( \4607 , \4605 , \4606 );
and \U$4265 ( \4608 , \4599 , \4607 );
and \U$4266 ( \4609 , \4591 , \4598 );
or \U$4267 ( \4610 , \4608 , \4609 );
and \U$4268 ( \4611 , \4584 , \4610 );
and \U$4269 ( \4612 , \4563 , \4583 );
or \U$4270 ( \4613 , \4611 , \4612 );
xor \U$4271 ( \4614 , \4535 , \4613 );
xor \U$4272 ( \4615 , \4316 , \4323 );
xor \U$4273 ( \4616 , \4615 , \4332 );
xor \U$4274 ( \4617 , \4279 , \4287 );
xor \U$4275 ( \4618 , \4617 , \4296 );
xor \U$4276 ( \4619 , \4616 , \4618 );
or \U$4277 ( \4620 , \4307 , \4300 );
nand \U$4278 ( \4621 , \4620 , \4308 );
and \U$4279 ( \4622 , \4619 , \4621 );
and \U$4280 ( \4623 , \4616 , \4618 );
nor \U$4281 ( \4624 , \4622 , \4623 );
xor \U$4282 ( \4625 , \4614 , \4624 );
and \U$4283 ( \4626 , \4454 , \4625 );
not \U$4284 ( \4627 , \4184 );
xor \U$4285 ( \4628 , \4209 , \4193 );
not \U$4286 ( \4629 , \4628 );
or \U$4287 ( \4630 , \4627 , \4629 );
or \U$4288 ( \4631 , \4628 , \4184 );
nand \U$4289 ( \4632 , \4630 , \4631 );
xor \U$4290 ( \4633 , \4250 , \4258 );
xor \U$4291 ( \4634 , \4633 , \4266 );
xor \U$4292 ( \4635 , \4632 , \4634 );
not \U$4293 ( \4636 , \4219 );
xor \U$4294 ( \4637 , \4237 , \4227 );
not \U$4295 ( \4638 , \4637 );
or \U$4296 ( \4639 , \4636 , \4638 );
or \U$4297 ( \4640 , \4637 , \4219 );
nand \U$4298 ( \4641 , \4639 , \4640 );
and \U$4299 ( \4642 , \4635 , \4641 );
and \U$4300 ( \4643 , \4632 , \4634 );
or \U$4301 ( \4644 , \4642 , \4643 );
not \U$4302 ( \4645 , \4644 );
xor \U$4303 ( \4646 , \4368 , \4378 );
xor \U$4304 ( \4647 , \4646 , \4389 );
not \U$4305 ( \4648 , \4647 );
or \U$4306 ( \4649 , \4645 , \4648 );
or \U$4307 ( \4650 , \4647 , \4644 );
nand \U$4308 ( \4651 , \4649 , \4650 );
not \U$4309 ( \4652 , \4651 );
xnor \U$4310 ( \4653 , \4343 , \4348 );
not \U$4311 ( \4654 , \4653 );
not \U$4312 ( \4655 , \4340 );
and \U$4313 ( \4656 , \4654 , \4655 );
and \U$4314 ( \4657 , \4653 , \4340 );
nor \U$4315 ( \4658 , \4656 , \4657 );
not \U$4316 ( \4659 , \4658 );
and \U$4317 ( \4660 , \4652 , \4659 );
and \U$4318 ( \4661 , \4651 , \4658 );
nor \U$4319 ( \4662 , \4660 , \4661 );
xor \U$4320 ( \4663 , \4535 , \4613 );
xor \U$4321 ( \4664 , \4663 , \4624 );
and \U$4322 ( \4665 , \4662 , \4664 );
and \U$4323 ( \4666 , \4454 , \4662 );
or \U$4324 ( \4667 , \4626 , \4665 , \4666 );
and \U$4325 ( \4668 , \2274 , RI986f340_49);
and \U$4326 ( \4669 , RI986f520_53, \2272 );
nor \U$4327 ( \4670 , \4668 , \4669 );
and \U$4328 ( \4671 , \4670 , \2030 );
not \U$4329 ( \4672 , \4670 );
and \U$4330 ( \4673 , \4672 , \2031 );
nor \U$4331 ( \4674 , \4671 , \4673 );
and \U$4332 ( \4675 , \2464 , RI986f610_55);
and \U$4333 ( \4676 , RI986df90_7, \2462 );
nor \U$4334 ( \4677 , \4675 , \4676 );
and \U$4335 ( \4678 , \4677 , \2468 );
not \U$4336 ( \4679 , \4677 );
and \U$4337 ( \4680 , \4679 , \2263 );
nor \U$4338 ( \4681 , \4678 , \4680 );
xor \U$4339 ( \4682 , \4674 , \4681 );
not \U$4340 ( \4683 , \2935 );
and \U$4341 ( \4684 , \3254 , RI986dea0_5);
and \U$4342 ( \4685 , RI986ddb0_3, \3252 );
nor \U$4343 ( \4686 , \4684 , \4685 );
not \U$4344 ( \4687 , \4686 );
or \U$4345 ( \4688 , \4683 , \4687 );
or \U$4346 ( \4689 , \4686 , \3406 );
nand \U$4347 ( \4690 , \4688 , \4689 );
and \U$4348 ( \4691 , \4682 , \4690 );
and \U$4349 ( \4692 , \4674 , \4681 );
or \U$4350 ( \4693 , \4691 , \4692 );
not \U$4351 ( \4694 , \3412 );
and \U$4352 ( \4695 , \3683 , RI986dcc0_1);
and \U$4353 ( \4696 , RI986e170_11, \3681 );
nor \U$4354 ( \4697 , \4695 , \4696 );
not \U$4355 ( \4698 , \4697 );
or \U$4356 ( \4699 , \4694 , \4698 );
or \U$4357 ( \4700 , \4697 , \3918 );
nand \U$4358 ( \4701 , \4699 , \4700 );
not \U$4359 ( \4702 , \4519 );
and \U$4360 ( \4703 , RI9872568_156, RI9872838_162);
not \U$4361 ( \4704 , RI9872838_162);
nor \U$4362 ( \4705 , \4704 , RI98728b0_163);
not \U$4363 ( \4706 , RI98728b0_163);
nor \U$4364 ( \4707 , \4706 , RI9872838_162);
or \U$4365 ( \4708 , \4705 , \4707 );
nor \U$4366 ( \4709 , RI9872568_156, RI9872838_162);
nor \U$4367 ( \4710 , \4703 , \4708 , \4709 );
nand \U$4368 ( \4711 , RI986e350_15, \4710 );
not \U$4369 ( \4712 , \4711 );
or \U$4370 ( \4713 , \4702 , \4712 );
or \U$4371 ( \4714 , \4711 , \4519 );
nand \U$4372 ( \4715 , \4713 , \4714 );
xor \U$4373 ( \4716 , \4701 , \4715 );
and \U$4374 ( \4717 , \4203 , RI986e080_9);
and \U$4375 ( \4718 , RI986e260_13, \4201 );
nor \U$4376 ( \4719 , \4717 , \4718 );
and \U$4377 ( \4720 , \4719 , \4207 );
not \U$4378 ( \4721 , \4719 );
and \U$4379 ( \4722 , \4721 , \3923 );
nor \U$4380 ( \4723 , \4720 , \4722 );
and \U$4381 ( \4724 , \4716 , \4723 );
and \U$4382 ( \4725 , \4701 , \4715 );
or \U$4383 ( \4726 , \4724 , \4725 );
xor \U$4384 ( \4727 , \4693 , \4726 );
and \U$4385 ( \4728 , \1329 , RI986e620_21);
and \U$4386 ( \4729 , RI986f7f0_59, \1327 );
nor \U$4387 ( \4730 , \4728 , \4729 );
and \U$4388 ( \4731 , \4730 , \1336 );
not \U$4389 ( \4732 , \4730 );
and \U$4390 ( \4733 , \4732 , \1337 );
nor \U$4391 ( \4734 , \4731 , \4733 );
and \U$4392 ( \4735 , \1311 , RI986f700_57);
and \U$4393 ( \4736 , RI986f9d0_63, \1309 );
nor \U$4394 ( \4737 , \4735 , \4736 );
and \U$4395 ( \4738 , \4737 , \1319 );
not \U$4396 ( \4739 , \4737 );
and \U$4397 ( \4740 , \4739 , \1318 );
nor \U$4398 ( \4741 , \4738 , \4740 );
xor \U$4399 ( \4742 , \4734 , \4741 );
not \U$4400 ( \4743 , \2034 );
and \U$4401 ( \4744 , \2042 , RI986f8e0_61);
and \U$4402 ( \4745 , RI986f430_51, \2040 );
nor \U$4403 ( \4746 , \4744 , \4745 );
not \U$4404 ( \4747 , \4746 );
or \U$4405 ( \4748 , \4743 , \4747 );
or \U$4406 ( \4749 , \4746 , \1462 );
nand \U$4407 ( \4750 , \4748 , \4749 );
and \U$4408 ( \4751 , \4742 , \4750 );
and \U$4409 ( \4752 , \4734 , \4741 );
or \U$4410 ( \4753 , \4751 , \4752 );
and \U$4411 ( \4754 , \4727 , \4753 );
and \U$4412 ( \4755 , \4693 , \4726 );
or \U$4413 ( \4756 , \4754 , \4755 );
and \U$4414 ( \4757 , \376 , RI986eda0_37);
and \U$4415 ( \4758 , RI986ebc0_33, \374 );
nor \U$4416 ( \4759 , \4757 , \4758 );
not \U$4417 ( \4760 , \4759 );
not \U$4418 ( \4761 , \365 );
and \U$4419 ( \4762 , \4760 , \4761 );
and \U$4420 ( \4763 , \4759 , \365 );
nor \U$4421 ( \4764 , \4762 , \4763 );
and \U$4422 ( \4765 , \395 , RI986e800_25);
and \U$4423 ( \4766 , RI986ee90_39, \393 );
nor \U$4424 ( \4767 , \4765 , \4766 );
not \U$4425 ( \4768 , \4767 );
not \U$4426 ( \4769 , \487 );
and \U$4427 ( \4770 , \4768 , \4769 );
and \U$4428 ( \4771 , \4767 , \386 );
nor \U$4429 ( \4772 , \4770 , \4771 );
or \U$4430 ( \4773 , \4764 , \4772 );
not \U$4431 ( \4774 , \4772 );
not \U$4432 ( \4775 , \4764 );
or \U$4433 ( \4776 , \4774 , \4775 );
not \U$4434 ( \4777 , \456 );
and \U$4435 ( \4778 , \465 , RI986ecb0_35);
and \U$4436 ( \4779 , RI986f070_43, \463 );
nor \U$4437 ( \4780 , \4778 , \4779 );
not \U$4438 ( \4781 , \4780 );
or \U$4439 ( \4782 , \4777 , \4781 );
or \U$4440 ( \4783 , \4780 , \454 );
nand \U$4441 ( \4784 , \4782 , \4783 );
nand \U$4442 ( \4785 , \4776 , \4784 );
nand \U$4443 ( \4786 , \4773 , \4785 );
and \U$4444 ( \4787 , \416 , RI98715f0_123);
and \U$4445 ( \4788 , RI986ead0_31, \414 );
nor \U$4446 ( \4789 , \4787 , \4788 );
and \U$4447 ( \4790 , \4789 , \421 );
not \U$4448 ( \4791 , \4789 );
and \U$4449 ( \4792 , \4791 , \422 );
nor \U$4450 ( \4793 , \4790 , \4792 );
nand \U$4451 ( \4794 , RI9871500_121, RI9871fc8_144);
or \U$4452 ( \4795 , \4793 , \4794 );
not \U$4453 ( \4796 , \4794 );
not \U$4454 ( \4797 , \4793 );
or \U$4455 ( \4798 , \4796 , \4797 );
not \U$4456 ( \4799 , \361 );
and \U$4457 ( \4800 , \354 , RI986e9e0_29);
and \U$4458 ( \4801 , RI986e8f0_27, \352 );
nor \U$4459 ( \4802 , \4800 , \4801 );
not \U$4460 ( \4803 , \4802 );
or \U$4461 ( \4804 , \4799 , \4803 );
or \U$4462 ( \4805 , \4802 , \345 );
nand \U$4463 ( \4806 , \4804 , \4805 );
nand \U$4464 ( \4807 , \4798 , \4806 );
nand \U$4465 ( \4808 , \4795 , \4807 );
xor \U$4466 ( \4809 , \4786 , \4808 );
and \U$4467 ( \4810 , \776 , RI986f160_45);
and \U$4468 ( \4811 , RI986e530_19, \774 );
nor \U$4469 ( \4812 , \4810 , \4811 );
and \U$4470 ( \4813 , \4812 , \474 );
not \U$4471 ( \4814 , \4812 );
and \U$4472 ( \4815 , \4814 , \451 );
nor \U$4473 ( \4816 , \4813 , \4815 );
and \U$4474 ( \4817 , \438 , RI986ef80_41);
and \U$4475 ( \4818 , RI986f250_47, \436 );
nor \U$4476 ( \4819 , \4817 , \4818 );
and \U$4477 ( \4820 , \4819 , \444 );
not \U$4478 ( \4821 , \4819 );
and \U$4479 ( \4822 , \4821 , \443 );
nor \U$4480 ( \4823 , \4820 , \4822 );
xor \U$4481 ( \4824 , \4816 , \4823 );
not \U$4482 ( \4825 , \1301 );
and \U$4483 ( \4826 , \1293 , RI986e440_17);
and \U$4484 ( \4827 , RI986e710_23, \1291 );
nor \U$4485 ( \4828 , \4826 , \4827 );
not \U$4486 ( \4829 , \4828 );
or \U$4487 ( \4830 , \4825 , \4829 );
or \U$4488 ( \4831 , \4828 , \1301 );
nand \U$4489 ( \4832 , \4830 , \4831 );
and \U$4490 ( \4833 , \4824 , \4832 );
and \U$4491 ( \4834 , \4816 , \4823 );
or \U$4492 ( \4835 , \4833 , \4834 );
and \U$4493 ( \4836 , \4809 , \4835 );
and \U$4494 ( \4837 , \4786 , \4808 );
or \U$4495 ( \4838 , \4836 , \4837 );
and \U$4496 ( \4839 , \4756 , \4838 );
not \U$4497 ( \4840 , \4756 );
not \U$4498 ( \4841 , \4838 );
and \U$4499 ( \4842 , \4840 , \4841 );
xor \U$4500 ( \4843 , \4543 , \4551 );
xor \U$4501 ( \4844 , \4843 , \4560 );
not \U$4502 ( \4845 , \4844 );
xor \U$4503 ( \4846 , \4591 , \4598 );
xor \U$4504 ( \4847 , \4846 , \4607 );
not \U$4505 ( \4848 , \4847 );
and \U$4506 ( \4849 , \4845 , \4848 );
and \U$4507 ( \4850 , \4847 , \4844 );
xor \U$4508 ( \4851 , \4570 , \4571 );
xor \U$4509 ( \4852 , \4851 , \4580 );
nor \U$4510 ( \4853 , \4850 , \4852 );
nor \U$4511 ( \4854 , \4849 , \4853 );
nor \U$4512 ( \4855 , \4842 , \4854 );
nor \U$4513 ( \4856 , \4839 , \4855 );
xor \U$4514 ( \4857 , \4563 , \4583 );
xor \U$4515 ( \4858 , \4857 , \4610 );
not \U$4516 ( \4859 , \4858 );
not \U$4517 ( \4860 , \4533 );
xor \U$4518 ( \4861 , \4506 , \4480 );
not \U$4519 ( \4862 , \4861 );
or \U$4520 ( \4863 , \4860 , \4862 );
or \U$4521 ( \4864 , \4861 , \4533 );
nand \U$4522 ( \4865 , \4863 , \4864 );
nand \U$4523 ( \4866 , \4859 , \4865 );
xor \U$4524 ( \4867 , \4856 , \4866 );
xor \U$4525 ( \4868 , \4632 , \4634 );
xor \U$4526 ( \4869 , \4868 , \4641 );
xor \U$4527 ( \4870 , \4616 , \4618 );
xor \U$4528 ( \4871 , \4870 , \4621 );
and \U$4529 ( \4872 , \4869 , \4871 );
not \U$4530 ( \4873 , \4869 );
not \U$4531 ( \4874 , \4871 );
and \U$4532 ( \4875 , \4873 , \4874 );
xor \U$4533 ( \4876 , \4488 , \4495 );
xor \U$4534 ( \4877 , \4876 , \4503 );
xor \U$4535 ( \4878 , \4462 , \4469 );
xor \U$4536 ( \4879 , \4878 , \4477 );
and \U$4537 ( \4880 , \4877 , \4879 );
not \U$4538 ( \4881 , \4879 );
not \U$4539 ( \4882 , \4877 );
and \U$4540 ( \4883 , \4881 , \4882 );
xor \U$4541 ( \4884 , \4517 , \4521 );
xor \U$4542 ( \4885 , \4884 , \4530 );
nor \U$4543 ( \4886 , \4883 , \4885 );
nor \U$4544 ( \4887 , \4880 , \4886 );
nor \U$4545 ( \4888 , \4875 , \4887 );
nor \U$4546 ( \4889 , \4872 , \4888 );
and \U$4547 ( \4890 , \4867 , \4889 );
and \U$4548 ( \4891 , \4856 , \4866 );
or \U$4549 ( \4892 , \4890 , \4891 );
or \U$4550 ( \4893 , \4667 , \4892 );
not \U$4551 ( \4894 , \4892 );
not \U$4552 ( \4895 , \4667 );
or \U$4553 ( \4896 , \4894 , \4895 );
xor \U$4554 ( \4897 , \4271 , \4338 );
xor \U$4555 ( \4898 , \4897 , \4350 );
xor \U$4556 ( \4899 , \4355 , \4357 );
xor \U$4557 ( \4900 , \4039 , \3758 );
xor \U$4558 ( \4901 , \4900 , \4042 );
xor \U$4559 ( \4902 , \4392 , \4399 );
xor \U$4560 ( \4903 , \4901 , \4902 );
xor \U$4561 ( \4904 , \4899 , \4903 );
xor \U$4562 ( \4905 , \4898 , \4904 );
nand \U$4563 ( \4906 , \4896 , \4905 );
nand \U$4564 ( \4907 , \4893 , \4906 );
xor \U$4565 ( \4908 , \4353 , \4358 );
xor \U$4566 ( \4909 , \4908 , \4404 );
xor \U$4567 ( \4910 , \4907 , \4909 );
xor \U$4568 ( \4911 , \4271 , \4338 );
xor \U$4569 ( \4912 , \4911 , \4350 );
and \U$4570 ( \4913 , \4899 , \4912 );
xor \U$4571 ( \4914 , \4271 , \4338 );
xor \U$4572 ( \4915 , \4914 , \4350 );
and \U$4573 ( \4916 , \4903 , \4915 );
and \U$4574 ( \4917 , \4899 , \4903 );
or \U$4575 ( \4918 , \4913 , \4916 , \4917 );
xor \U$4576 ( \4919 , \4535 , \4613 );
and \U$4577 ( \4920 , \4919 , \4624 );
and \U$4578 ( \4921 , \4535 , \4613 );
or \U$4579 ( \4922 , \4920 , \4921 );
not \U$4580 ( \4923 , \4450 );
nand \U$4581 ( \4924 , \4923 , \4439 );
or \U$4582 ( \4925 , \4922 , \4924 );
not \U$4583 ( \4926 , \4924 );
not \U$4584 ( \4927 , \4922 );
or \U$4585 ( \4928 , \4926 , \4927 );
or \U$4586 ( \4929 , \4658 , \4647 );
not \U$4587 ( \4930 , \4658 );
not \U$4588 ( \4931 , \4647 );
or \U$4589 ( \4932 , \4930 , \4931 );
nand \U$4590 ( \4933 , \4932 , \4644 );
nand \U$4591 ( \4934 , \4929 , \4933 );
nand \U$4592 ( \4935 , \4928 , \4934 );
nand \U$4593 ( \4936 , \4925 , \4935 );
xor \U$4594 ( \4937 , \4918 , \4936 );
xor \U$4595 ( \4938 , \3968 , \4036 );
xor \U$4596 ( \4939 , \4938 , \4045 );
xor \U$4597 ( \4940 , \4158 , \4171 );
xor \U$4598 ( \4941 , \4939 , \4940 );
xor \U$4599 ( \4942 , \4937 , \4941 );
and \U$4600 ( \4943 , \4910 , \4942 );
and \U$4601 ( \4944 , \4907 , \4909 );
or \U$4602 ( \4945 , \4943 , \4944 );
xor \U$4603 ( \4946 , \4176 , \4407 );
xor \U$4604 ( \4947 , \4946 , \4414 );
not \U$4605 ( \4948 , \4053 );
not \U$4606 ( \4949 , \4096 );
not \U$4607 ( \4950 , \4048 );
and \U$4608 ( \4951 , \4949 , \4950 );
and \U$4609 ( \4952 , \4096 , \4048 );
nor \U$4610 ( \4953 , \4951 , \4952 );
not \U$4611 ( \4954 , \4953 );
or \U$4612 ( \4955 , \4948 , \4954 );
or \U$4613 ( \4956 , \4953 , \4053 );
nand \U$4614 ( \4957 , \4955 , \4956 );
xor \U$4615 ( \4958 , \4918 , \4936 );
and \U$4616 ( \4959 , \4958 , \4941 );
and \U$4617 ( \4960 , \4918 , \4936 );
or \U$4618 ( \4961 , \4959 , \4960 );
xor \U$4619 ( \4962 , \4957 , \4961 );
xor \U$4620 ( \4963 , \4947 , \4962 );
xor \U$4621 ( \4964 , \4945 , \4963 );
xor \U$4622 ( \4965 , \4907 , \4909 );
xor \U$4623 ( \4966 , \4965 , \4942 );
not \U$4624 ( \4967 , \4966 );
xnor \U$4625 ( \4968 , \4892 , \4667 );
not \U$4626 ( \4969 , \4968 );
not \U$4627 ( \4970 , \4905 );
and \U$4628 ( \4971 , \4969 , \4970 );
and \U$4629 ( \4972 , \4968 , \4905 );
nor \U$4630 ( \4973 , \4971 , \4972 );
not \U$4631 ( \4974 , \4922 );
not \U$4632 ( \4975 , \4934 );
or \U$4633 ( \4976 , \4974 , \4975 );
or \U$4634 ( \4977 , \4934 , \4922 );
nand \U$4635 ( \4978 , \4976 , \4977 );
not \U$4636 ( \4979 , \4978 );
not \U$4637 ( \4980 , \4924 );
and \U$4638 ( \4981 , \4979 , \4980 );
and \U$4639 ( \4982 , \4978 , \4924 );
nor \U$4640 ( \4983 , \4981 , \4982 );
xor \U$4641 ( \4984 , \4973 , \4983 );
not \U$4642 ( \4985 , \4865 );
not \U$4643 ( \4986 , \4858 );
or \U$4644 ( \4987 , \4985 , \4986 );
or \U$4645 ( \4988 , \4858 , \4865 );
nand \U$4646 ( \4989 , \4987 , \4988 );
not \U$4647 ( \4990 , \4854 );
xor \U$4648 ( \4991 , \4756 , \4838 );
not \U$4649 ( \4992 , \4991 );
or \U$4650 ( \4993 , \4990 , \4992 );
or \U$4651 ( \4994 , \4991 , \4854 );
nand \U$4652 ( \4995 , \4993 , \4994 );
xor \U$4653 ( \4996 , \4989 , \4995 );
not \U$4654 ( \4997 , \4871 );
not \U$4655 ( \4998 , \4869 );
not \U$4656 ( \4999 , \4887 );
and \U$4657 ( \5000 , \4998 , \4999 );
and \U$4658 ( \5001 , \4869 , \4887 );
nor \U$4659 ( \5002 , \5000 , \5001 );
not \U$4660 ( \5003 , \5002 );
or \U$4661 ( \5004 , \4997 , \5003 );
or \U$4662 ( \5005 , \5002 , \4871 );
nand \U$4663 ( \5006 , \5004 , \5005 );
and \U$4664 ( \5007 , \4996 , \5006 );
and \U$4665 ( \5008 , \4989 , \4995 );
nor \U$4666 ( \5009 , \5007 , \5008 );
xor \U$4667 ( \5010 , \4693 , \4726 );
xor \U$4668 ( \5011 , \5010 , \4753 );
xor \U$4669 ( \5012 , \4786 , \4808 );
xor \U$4670 ( \5013 , \5012 , \4835 );
and \U$4671 ( \5014 , \5011 , \5013 );
and \U$4672 ( \5015 , \2274 , RI986f430_51);
and \U$4673 ( \5016 , RI986f340_49, \2272 );
nor \U$4674 ( \5017 , \5015 , \5016 );
and \U$4675 ( \5018 , \5017 , \2030 );
not \U$4676 ( \5019 , \5017 );
and \U$4677 ( \5020 , \5019 , \2031 );
nor \U$4678 ( \5021 , \5018 , \5020 );
and \U$4679 ( \5022 , \1311 , RI986f7f0_59);
and \U$4680 ( \5023 , RI986f700_57, \1309 );
nor \U$4681 ( \5024 , \5022 , \5023 );
and \U$4682 ( \5025 , \5024 , \1458 );
not \U$4683 ( \5026 , \5024 );
and \U$4684 ( \5027 , \5026 , \1315 );
nor \U$4685 ( \5028 , \5025 , \5027 );
xor \U$4686 ( \5029 , \5021 , \5028 );
not \U$4687 ( \5030 , \2034 );
and \U$4688 ( \5031 , \2042 , RI986f9d0_63);
and \U$4689 ( \5032 , RI986f8e0_61, \2040 );
nor \U$4690 ( \5033 , \5031 , \5032 );
not \U$4691 ( \5034 , \5033 );
or \U$4692 ( \5035 , \5030 , \5034 );
or \U$4693 ( \5036 , \5033 , \2034 );
nand \U$4694 ( \5037 , \5035 , \5036 );
and \U$4695 ( \5038 , \5029 , \5037 );
and \U$4696 ( \5039 , \5021 , \5028 );
or \U$4697 ( \5040 , \5038 , \5039 );
not \U$4698 ( \5041 , \4519 );
and \U$4699 ( \5042 , \4710 , RI986e260_13);
and \U$4700 ( \5043 , RI986e350_15, \4708 );
nor \U$4701 ( \5044 , \5042 , \5043 );
not \U$4702 ( \5045 , \5044 );
or \U$4703 ( \5046 , \5041 , \5045 );
or \U$4704 ( \5047 , \5044 , \4521 );
nand \U$4705 ( \5048 , \5046 , \5047 );
not \U$4706 ( \5049 , RI98729a0_165);
not \U$4707 ( \5050 , RI9872928_164);
or \U$4708 ( \5051 , \5049 , \5050 );
nand \U$4709 ( \5052 , \5051 , RI98728b0_163);
xor \U$4710 ( \5053 , \5048 , \5052 );
and \U$4711 ( \5054 , \4203 , RI986e170_11);
and \U$4712 ( \5055 , RI986e080_9, \4201 );
nor \U$4713 ( \5056 , \5054 , \5055 );
and \U$4714 ( \5057 , \5056 , \4207 );
not \U$4715 ( \5058 , \5056 );
and \U$4716 ( \5059 , \5058 , \3922 );
nor \U$4717 ( \5060 , \5057 , \5059 );
and \U$4718 ( \5061 , \5053 , \5060 );
and \U$4719 ( \5062 , \5048 , \5052 );
or \U$4720 ( \5063 , \5061 , \5062 );
xor \U$4721 ( \5064 , \5040 , \5063 );
not \U$4722 ( \5065 , \3918 );
and \U$4723 ( \5066 , \3683 , RI986ddb0_3);
and \U$4724 ( \5067 , RI986dcc0_1, \3681 );
nor \U$4725 ( \5068 , \5066 , \5067 );
not \U$4726 ( \5069 , \5068 );
or \U$4727 ( \5070 , \5065 , \5069 );
or \U$4728 ( \5071 , \5068 , \3412 );
nand \U$4729 ( \5072 , \5070 , \5071 );
and \U$4730 ( \5073 , \2464 , RI986f520_53);
and \U$4731 ( \5074 , RI986f610_55, \2462 );
nor \U$4732 ( \5075 , \5073 , \5074 );
and \U$4733 ( \5076 , \5075 , \2468 );
not \U$4734 ( \5077 , \5075 );
and \U$4735 ( \5078 , \5077 , \2263 );
nor \U$4736 ( \5079 , \5076 , \5078 );
xor \U$4737 ( \5080 , \5072 , \5079 );
not \U$4738 ( \5081 , \3406 );
and \U$4739 ( \5082 , \3254 , RI986df90_7);
and \U$4740 ( \5083 , RI986dea0_5, \3252 );
nor \U$4741 ( \5084 , \5082 , \5083 );
not \U$4742 ( \5085 , \5084 );
or \U$4743 ( \5086 , \5081 , \5085 );
or \U$4744 ( \5087 , \5084 , \2935 );
nand \U$4745 ( \5088 , \5086 , \5087 );
and \U$4746 ( \5089 , \5080 , \5088 );
and \U$4747 ( \5090 , \5072 , \5079 );
or \U$4748 ( \5091 , \5089 , \5090 );
and \U$4749 ( \5092 , \5064 , \5091 );
and \U$4750 ( \5093 , \5040 , \5063 );
or \U$4751 ( \5094 , \5092 , \5093 );
not \U$4752 ( \5095 , \4793 );
not \U$4753 ( \5096 , \4806 );
or \U$4754 ( \5097 , \5095 , \5096 );
or \U$4755 ( \5098 , \4793 , \4806 );
nand \U$4756 ( \5099 , \5097 , \5098 );
not \U$4757 ( \5100 , \5099 );
not \U$4758 ( \5101 , \4794 );
and \U$4759 ( \5102 , \5100 , \5101 );
and \U$4760 ( \5103 , \5099 , \4794 );
nor \U$4761 ( \5104 , \5102 , \5103 );
not \U$4762 ( \5105 , \4764 );
not \U$4763 ( \5106 , \4784 );
or \U$4764 ( \5107 , \5105 , \5106 );
or \U$4765 ( \5108 , \4764 , \4784 );
nand \U$4766 ( \5109 , \5107 , \5108 );
not \U$4767 ( \5110 , \5109 );
not \U$4768 ( \5111 , \4772 );
and \U$4769 ( \5112 , \5110 , \5111 );
and \U$4770 ( \5113 , \5109 , \4772 );
nor \U$4771 ( \5114 , \5112 , \5113 );
nand \U$4772 ( \5115 , \5104 , \5114 );
xor \U$4773 ( \5116 , \5094 , \5115 );
and \U$4774 ( \5117 , \438 , RI986f070_43);
and \U$4775 ( \5118 , RI986ef80_41, \436 );
nor \U$4776 ( \5119 , \5117 , \5118 );
and \U$4777 ( \5120 , \5119 , \444 );
not \U$4778 ( \5121 , \5119 );
and \U$4779 ( \5122 , \5121 , \443 );
nor \U$4780 ( \5123 , \5120 , \5122 );
not \U$4781 ( \5124 , \456 );
and \U$4782 ( \5125 , \465 , RI986ebc0_33);
and \U$4783 ( \5126 , RI986ecb0_35, \463 );
nor \U$4784 ( \5127 , \5125 , \5126 );
not \U$4785 ( \5128 , \5127 );
or \U$4786 ( \5129 , \5124 , \5128 );
or \U$4787 ( \5130 , \5127 , \454 );
nand \U$4788 ( \5131 , \5129 , \5130 );
xor \U$4789 ( \5132 , \5123 , \5131 );
not \U$4790 ( \5133 , \367 );
and \U$4791 ( \5134 , \376 , RI986ee90_39);
and \U$4792 ( \5135 , RI986eda0_37, \374 );
nor \U$4793 ( \5136 , \5134 , \5135 );
not \U$4794 ( \5137 , \5136 );
or \U$4795 ( \5138 , \5133 , \5137 );
or \U$4796 ( \5139 , \5136 , \367 );
nand \U$4797 ( \5140 , \5138 , \5139 );
and \U$4798 ( \5141 , \5132 , \5140 );
and \U$4799 ( \5142 , \5123 , \5131 );
or \U$4800 ( \5143 , \5141 , \5142 );
not \U$4801 ( \5144 , \345 );
and \U$4802 ( \5145 , \354 , RI986ead0_31);
and \U$4803 ( \5146 , RI986e9e0_29, \352 );
nor \U$4804 ( \5147 , \5145 , \5146 );
not \U$4805 ( \5148 , \5147 );
or \U$4806 ( \5149 , \5144 , \5148 );
or \U$4807 ( \5150 , \5147 , \345 );
nand \U$4808 ( \5151 , \5149 , \5150 );
not \U$4809 ( \5152 , \386 );
and \U$4810 ( \5153 , \395 , RI986e8f0_27);
and \U$4811 ( \5154 , RI986e800_25, \393 );
nor \U$4812 ( \5155 , \5153 , \5154 );
not \U$4813 ( \5156 , \5155 );
or \U$4814 ( \5157 , \5152 , \5156 );
or \U$4815 ( \5158 , \5155 , \386 );
nand \U$4816 ( \5159 , \5157 , \5158 );
xor \U$4817 ( \5160 , \5151 , \5159 );
and \U$4818 ( \5161 , \416 , RI9871500_121);
and \U$4819 ( \5162 , RI98715f0_123, \414 );
nor \U$4820 ( \5163 , \5161 , \5162 );
and \U$4821 ( \5164 , \5163 , \422 );
not \U$4822 ( \5165 , \5163 );
and \U$4823 ( \5166 , \5165 , \421 );
nor \U$4824 ( \5167 , \5164 , \5166 );
and \U$4825 ( \5168 , \5160 , \5167 );
and \U$4826 ( \5169 , \5151 , \5159 );
or \U$4827 ( \5170 , \5168 , \5169 );
xor \U$4828 ( \5171 , \5143 , \5170 );
and \U$4829 ( \5172 , \776 , RI986f250_47);
and \U$4830 ( \5173 , RI986f160_45, \774 );
nor \U$4831 ( \5174 , \5172 , \5173 );
and \U$4832 ( \5175 , \5174 , \474 );
not \U$4833 ( \5176 , \5174 );
and \U$4834 ( \5177 , \5176 , \451 );
nor \U$4835 ( \5178 , \5175 , \5177 );
not \U$4836 ( \5179 , \1301 );
and \U$4837 ( \5180 , \1293 , RI986e530_19);
and \U$4838 ( \5181 , RI986e440_17, \1291 );
nor \U$4839 ( \5182 , \5180 , \5181 );
not \U$4840 ( \5183 , \5182 );
or \U$4841 ( \5184 , \5179 , \5183 );
or \U$4842 ( \5185 , \5182 , \1301 );
nand \U$4843 ( \5186 , \5184 , \5185 );
xor \U$4844 ( \5187 , \5178 , \5186 );
and \U$4845 ( \5188 , \1329 , RI986e710_23);
and \U$4846 ( \5189 , RI986e620_21, \1327 );
nor \U$4847 ( \5190 , \5188 , \5189 );
and \U$4848 ( \5191 , \5190 , \1336 );
not \U$4849 ( \5192 , \5190 );
and \U$4850 ( \5193 , \5192 , \1337 );
nor \U$4851 ( \5194 , \5191 , \5193 );
and \U$4852 ( \5195 , \5187 , \5194 );
and \U$4853 ( \5196 , \5178 , \5186 );
or \U$4854 ( \5197 , \5195 , \5196 );
and \U$4855 ( \5198 , \5171 , \5197 );
and \U$4856 ( \5199 , \5143 , \5170 );
or \U$4857 ( \5200 , \5198 , \5199 );
and \U$4858 ( \5201 , \5116 , \5200 );
and \U$4859 ( \5202 , \5094 , \5115 );
or \U$4860 ( \5203 , \5201 , \5202 );
xor \U$4861 ( \5204 , \5014 , \5203 );
not \U$4862 ( \5205 , \4847 );
xor \U$4863 ( \5206 , \4852 , \4844 );
not \U$4864 ( \5207 , \5206 );
or \U$4865 ( \5208 , \5205 , \5207 );
or \U$4866 ( \5209 , \5206 , \4847 );
nand \U$4867 ( \5210 , \5208 , \5209 );
xor \U$4868 ( \5211 , \4816 , \4823 );
xor \U$4869 ( \5212 , \5211 , \4832 );
xor \U$4870 ( \5213 , \4674 , \4681 );
xor \U$4871 ( \5214 , \5213 , \4690 );
and \U$4872 ( \5215 , \5212 , \5214 );
xor \U$4873 ( \5216 , \4734 , \4741 );
xor \U$4874 ( \5217 , \5216 , \4750 );
xor \U$4875 ( \5218 , \4674 , \4681 );
xor \U$4876 ( \5219 , \5218 , \4690 );
and \U$4877 ( \5220 , \5217 , \5219 );
and \U$4878 ( \5221 , \5212 , \5217 );
or \U$4879 ( \5222 , \5215 , \5220 , \5221 );
xor \U$4880 ( \5223 , \5210 , \5222 );
not \U$4881 ( \5224 , \4885 );
xor \U$4882 ( \5225 , \4877 , \4879 );
not \U$4883 ( \5226 , \5225 );
or \U$4884 ( \5227 , \5224 , \5226 );
or \U$4885 ( \5228 , \5225 , \4885 );
nand \U$4886 ( \5229 , \5227 , \5228 );
and \U$4887 ( \5230 , \5223 , \5229 );
and \U$4888 ( \5231 , \5210 , \5222 );
or \U$4889 ( \5232 , \5230 , \5231 );
and \U$4890 ( \5233 , \5204 , \5232 );
and \U$4891 ( \5234 , \5014 , \5203 );
nor \U$4892 ( \5235 , \5233 , \5234 );
xor \U$4893 ( \5236 , \5009 , \5235 );
xor \U$4894 ( \5237 , \4535 , \4613 );
xor \U$4895 ( \5238 , \5237 , \4624 );
xor \U$4896 ( \5239 , \4454 , \4662 );
xor \U$4897 ( \5240 , \5238 , \5239 );
and \U$4898 ( \5241 , \5236 , \5240 );
and \U$4899 ( \5242 , \5009 , \5235 );
or \U$4900 ( \5243 , \5241 , \5242 );
and \U$4901 ( \5244 , \4984 , \5243 );
and \U$4902 ( \5245 , \4973 , \4983 );
or \U$4903 ( \5246 , \5244 , \5245 );
nor \U$4904 ( \5247 , \4967 , \5246 );
and \U$4905 ( \5248 , \4964 , \5247 );
xor \U$4906 ( \5249 , \5247 , \4964 );
not \U$4907 ( \5250 , \4966 );
not \U$4908 ( \5251 , \5246 );
and \U$4909 ( \5252 , \5250 , \5251 );
and \U$4910 ( \5253 , \4966 , \5246 );
nor \U$4911 ( \5254 , \5252 , \5253 );
xor \U$4912 ( \5255 , \4973 , \4983 );
xor \U$4913 ( \5256 , \5255 , \5243 );
not \U$4914 ( \5257 , \5256 );
xor \U$4915 ( \5258 , \5009 , \5235 );
xor \U$4916 ( \5259 , \5258 , \5240 );
xor \U$4917 ( \5260 , \4856 , \4866 );
xor \U$4918 ( \5261 , \5260 , \4889 );
or \U$4919 ( \5262 , \5259 , \5261 );
not \U$4920 ( \5263 , \5261 );
not \U$4921 ( \5264 , \5259 );
or \U$4922 ( \5265 , \5263 , \5264 );
or \U$4923 ( \5266 , \5104 , \5114 );
nand \U$4924 ( \5267 , \5266 , \5115 );
xor \U$4925 ( \5268 , \5040 , \5063 );
xor \U$4926 ( \5269 , \5268 , \5091 );
and \U$4927 ( \5270 , \5267 , \5269 );
xor \U$4928 ( \5271 , \5143 , \5170 );
xor \U$4929 ( \5272 , \5271 , \5197 );
xor \U$4930 ( \5273 , \5040 , \5063 );
xor \U$4931 ( \5274 , \5273 , \5091 );
and \U$4932 ( \5275 , \5272 , \5274 );
and \U$4933 ( \5276 , \5267 , \5272 );
or \U$4934 ( \5277 , \5270 , \5275 , \5276 );
not \U$4935 ( \5278 , \2034 );
and \U$4936 ( \5279 , \2042 , RI986f700_57);
and \U$4937 ( \5280 , RI986f9d0_63, \2040 );
nor \U$4938 ( \5281 , \5279 , \5280 );
not \U$4939 ( \5282 , \5281 );
or \U$4940 ( \5283 , \5278 , \5282 );
or \U$4941 ( \5284 , \5281 , \2034 );
nand \U$4942 ( \5285 , \5283 , \5284 );
and \U$4943 ( \5286 , \1311 , RI986e620_21);
and \U$4944 ( \5287 , RI986f7f0_59, \1309 );
nor \U$4945 ( \5288 , \5286 , \5287 );
and \U$4946 ( \5289 , \5288 , \1458 );
not \U$4947 ( \5290 , \5288 );
and \U$4948 ( \5291 , \5290 , \1318 );
nor \U$4949 ( \5292 , \5289 , \5291 );
xor \U$4950 ( \5293 , \5285 , \5292 );
and \U$4951 ( \5294 , \2274 , RI986f8e0_61);
and \U$4952 ( \5295 , RI986f430_51, \2272 );
nor \U$4953 ( \5296 , \5294 , \5295 );
and \U$4954 ( \5297 , \5296 , \2030 );
not \U$4955 ( \5298 , \5296 );
and \U$4956 ( \5299 , \5298 , \2031 );
nor \U$4957 ( \5300 , \5297 , \5299 );
and \U$4958 ( \5301 , \5293 , \5300 );
and \U$4959 ( \5302 , \5285 , \5292 );
or \U$4960 ( \5303 , \5301 , \5302 );
and \U$4961 ( \5304 , \4203 , RI986dcc0_1);
and \U$4962 ( \5305 , RI986e170_11, \4201 );
nor \U$4963 ( \5306 , \5304 , \5305 );
and \U$4964 ( \5307 , \5306 , \4207 );
not \U$4965 ( \5308 , \5306 );
and \U$4966 ( \5309 , \5308 , \3922 );
nor \U$4967 ( \5310 , \5307 , \5309 );
and \U$4968 ( \5311 , RI98728b0_163, RI9872928_164);
not \U$4969 ( \5312 , RI9872928_164);
nor \U$4970 ( \5313 , \5312 , RI98729a0_165);
not \U$4971 ( \5314 , RI98729a0_165);
nor \U$4972 ( \5315 , \5314 , RI9872928_164);
or \U$4973 ( \5316 , \5313 , \5315 );
nor \U$4974 ( \5317 , RI98728b0_163, RI9872928_164);
nor \U$4975 ( \5318 , \5311 , \5316 , \5317 );
nand \U$4976 ( \5319 , RI986e350_15, \5318 );
and \U$4977 ( \5320 , \5319 , \5052 );
not \U$4978 ( \5321 , \5319 );
not \U$4979 ( \5322 , \5052 );
and \U$4980 ( \5323 , \5321 , \5322 );
nor \U$4981 ( \5324 , \5320 , \5323 );
xor \U$4982 ( \5325 , \5310 , \5324 );
not \U$4983 ( \5326 , \4519 );
and \U$4984 ( \5327 , \4710 , RI986e080_9);
and \U$4985 ( \5328 , RI986e260_13, \4708 );
nor \U$4986 ( \5329 , \5327 , \5328 );
not \U$4987 ( \5330 , \5329 );
or \U$4988 ( \5331 , \5326 , \5330 );
or \U$4989 ( \5332 , \5329 , \4521 );
nand \U$4990 ( \5333 , \5331 , \5332 );
and \U$4991 ( \5334 , \5325 , \5333 );
and \U$4992 ( \5335 , \5310 , \5324 );
or \U$4993 ( \5336 , \5334 , \5335 );
xor \U$4994 ( \5337 , \5303 , \5336 );
not \U$4995 ( \5338 , \3918 );
and \U$4996 ( \5339 , \3683 , RI986dea0_5);
and \U$4997 ( \5340 , RI986ddb0_3, \3681 );
nor \U$4998 ( \5341 , \5339 , \5340 );
not \U$4999 ( \5342 , \5341 );
or \U$5000 ( \5343 , \5338 , \5342 );
or \U$5001 ( \5344 , \5341 , \3918 );
nand \U$5002 ( \5345 , \5343 , \5344 );
and \U$5003 ( \5346 , \2464 , RI986f340_49);
and \U$5004 ( \5347 , RI986f520_53, \2462 );
nor \U$5005 ( \5348 , \5346 , \5347 );
and \U$5006 ( \5349 , \5348 , \2468 );
not \U$5007 ( \5350 , \5348 );
and \U$5008 ( \5351 , \5350 , \2263 );
nor \U$5009 ( \5352 , \5349 , \5351 );
xor \U$5010 ( \5353 , \5345 , \5352 );
not \U$5011 ( \5354 , \2935 );
and \U$5012 ( \5355 , \3254 , RI986f610_55);
and \U$5013 ( \5356 , RI986df90_7, \3252 );
nor \U$5014 ( \5357 , \5355 , \5356 );
not \U$5015 ( \5358 , \5357 );
or \U$5016 ( \5359 , \5354 , \5358 );
or \U$5017 ( \5360 , \5357 , \2935 );
nand \U$5018 ( \5361 , \5359 , \5360 );
and \U$5019 ( \5362 , \5353 , \5361 );
and \U$5020 ( \5363 , \5345 , \5352 );
or \U$5021 ( \5364 , \5362 , \5363 );
and \U$5022 ( \5365 , \5337 , \5364 );
and \U$5023 ( \5366 , \5303 , \5336 );
or \U$5024 ( \5367 , \5365 , \5366 );
not \U$5025 ( \5368 , \1301 );
and \U$5026 ( \5369 , \1293 , RI986f160_45);
and \U$5027 ( \5370 , RI986e530_19, \1291 );
nor \U$5028 ( \5371 , \5369 , \5370 );
not \U$5029 ( \5372 , \5371 );
or \U$5030 ( \5373 , \5368 , \5372 );
or \U$5031 ( \5374 , \5371 , \1128 );
nand \U$5032 ( \5375 , \5373 , \5374 );
and \U$5033 ( \5376 , \776 , RI986ef80_41);
and \U$5034 ( \5377 , RI986f250_47, \774 );
nor \U$5035 ( \5378 , \5376 , \5377 );
and \U$5036 ( \5379 , \5378 , \474 );
not \U$5037 ( \5380 , \5378 );
and \U$5038 ( \5381 , \5380 , \451 );
nor \U$5039 ( \5382 , \5379 , \5381 );
xor \U$5040 ( \5383 , \5375 , \5382 );
and \U$5041 ( \5384 , \1329 , RI986e440_17);
and \U$5042 ( \5385 , RI986e710_23, \1327 );
nor \U$5043 ( \5386 , \5384 , \5385 );
and \U$5044 ( \5387 , \5386 , \1336 );
not \U$5045 ( \5388 , \5386 );
and \U$5046 ( \5389 , \5388 , \1337 );
nor \U$5047 ( \5390 , \5387 , \5389 );
and \U$5048 ( \5391 , \5383 , \5390 );
and \U$5049 ( \5392 , \5375 , \5382 );
or \U$5050 ( \5393 , \5391 , \5392 );
and \U$5051 ( \5394 , \354 , RI98715f0_123);
and \U$5052 ( \5395 , RI986ead0_31, \352 );
nor \U$5053 ( \5396 , \5394 , \5395 );
not \U$5054 ( \5397 , \5396 );
not \U$5055 ( \5398 , \361 );
and \U$5056 ( \5399 , \5397 , \5398 );
and \U$5057 ( \5400 , \5396 , \361 );
nor \U$5058 ( \5401 , \5399 , \5400 );
and \U$5059 ( \5402 , \416 , RI98717d0_127);
and \U$5060 ( \5403 , RI9871500_121, \414 );
nor \U$5061 ( \5404 , \5402 , \5403 );
and \U$5062 ( \5405 , \5404 , \421 );
not \U$5063 ( \5406 , \5404 );
and \U$5064 ( \5407 , \5406 , \422 );
nor \U$5065 ( \5408 , \5405 , \5407 );
or \U$5066 ( \5409 , \5401 , \5408 );
not \U$5067 ( \5410 , \5408 );
not \U$5068 ( \5411 , \5401 );
or \U$5069 ( \5412 , \5410 , \5411 );
not \U$5070 ( \5413 , \487 );
and \U$5071 ( \5414 , \395 , RI986e9e0_29);
and \U$5072 ( \5415 , RI986e8f0_27, \393 );
nor \U$5073 ( \5416 , \5414 , \5415 );
not \U$5074 ( \5417 , \5416 );
or \U$5075 ( \5418 , \5413 , \5417 );
or \U$5076 ( \5419 , \5416 , \487 );
nand \U$5077 ( \5420 , \5418 , \5419 );
nand \U$5078 ( \5421 , \5412 , \5420 );
nand \U$5079 ( \5422 , \5409 , \5421 );
xor \U$5080 ( \5423 , \5393 , \5422 );
not \U$5081 ( \5424 , \365 );
and \U$5082 ( \5425 , \376 , RI986e800_25);
and \U$5083 ( \5426 , RI986ee90_39, \374 );
nor \U$5084 ( \5427 , \5425 , \5426 );
not \U$5085 ( \5428 , \5427 );
or \U$5086 ( \5429 , \5424 , \5428 );
or \U$5087 ( \5430 , \5427 , \367 );
nand \U$5088 ( \5431 , \5429 , \5430 );
and \U$5089 ( \5432 , \438 , RI986ecb0_35);
and \U$5090 ( \5433 , RI986f070_43, \436 );
nor \U$5091 ( \5434 , \5432 , \5433 );
and \U$5092 ( \5435 , \5434 , \444 );
not \U$5093 ( \5436 , \5434 );
and \U$5094 ( \5437 , \5436 , \443 );
nor \U$5095 ( \5438 , \5435 , \5437 );
xor \U$5096 ( \5439 , \5431 , \5438 );
not \U$5097 ( \5440 , \454 );
and \U$5098 ( \5441 , \465 , RI986eda0_37);
and \U$5099 ( \5442 , RI986ebc0_33, \463 );
nor \U$5100 ( \5443 , \5441 , \5442 );
not \U$5101 ( \5444 , \5443 );
or \U$5102 ( \5445 , \5440 , \5444 );
or \U$5103 ( \5446 , \5443 , \454 );
nand \U$5104 ( \5447 , \5445 , \5446 );
and \U$5105 ( \5448 , \5439 , \5447 );
and \U$5106 ( \5449 , \5431 , \5438 );
or \U$5107 ( \5450 , \5448 , \5449 );
and \U$5108 ( \5451 , \5423 , \5450 );
and \U$5109 ( \5452 , \5393 , \5422 );
or \U$5110 ( \5453 , \5451 , \5452 );
xor \U$5111 ( \5454 , \5367 , \5453 );
not \U$5112 ( \5455 , RI98717d0_127);
nor \U$5113 ( \5456 , \5455 , \407 );
xor \U$5114 ( \5457 , \5123 , \5131 );
xor \U$5115 ( \5458 , \5457 , \5140 );
and \U$5116 ( \5459 , \5456 , \5458 );
xor \U$5117 ( \5460 , \5151 , \5159 );
xor \U$5118 ( \5461 , \5460 , \5167 );
xor \U$5119 ( \5462 , \5123 , \5131 );
xor \U$5120 ( \5463 , \5462 , \5140 );
and \U$5121 ( \5464 , \5461 , \5463 );
and \U$5122 ( \5465 , \5456 , \5461 );
or \U$5123 ( \5466 , \5459 , \5464 , \5465 );
and \U$5124 ( \5467 , \5454 , \5466 );
and \U$5125 ( \5468 , \5367 , \5453 );
or \U$5126 ( \5469 , \5467 , \5468 );
xor \U$5127 ( \5470 , \5277 , \5469 );
xor \U$5128 ( \5471 , \5178 , \5186 );
xor \U$5129 ( \5472 , \5471 , \5194 );
xor \U$5130 ( \5473 , \5072 , \5079 );
xor \U$5131 ( \5474 , \5473 , \5088 );
and \U$5132 ( \5475 , \5472 , \5474 );
xor \U$5133 ( \5476 , \5021 , \5028 );
xor \U$5134 ( \5477 , \5476 , \5037 );
xor \U$5135 ( \5478 , \5072 , \5079 );
xor \U$5136 ( \5479 , \5478 , \5088 );
and \U$5137 ( \5480 , \5477 , \5479 );
and \U$5138 ( \5481 , \5472 , \5477 );
or \U$5139 ( \5482 , \5475 , \5480 , \5481 );
xor \U$5140 ( \5483 , \4701 , \4715 );
xor \U$5141 ( \5484 , \5483 , \4723 );
xor \U$5142 ( \5485 , \5482 , \5484 );
xor \U$5143 ( \5486 , \4674 , \4681 );
xor \U$5144 ( \5487 , \5486 , \4690 );
xor \U$5145 ( \5488 , \5212 , \5217 );
xor \U$5146 ( \5489 , \5487 , \5488 );
and \U$5147 ( \5490 , \5485 , \5489 );
and \U$5148 ( \5491 , \5482 , \5484 );
or \U$5149 ( \5492 , \5490 , \5491 );
and \U$5150 ( \5493 , \5470 , \5492 );
and \U$5151 ( \5494 , \5277 , \5469 );
or \U$5152 ( \5495 , \5493 , \5494 );
xor \U$5153 ( \5496 , \5011 , \5013 );
xor \U$5154 ( \5497 , \5094 , \5115 );
xor \U$5155 ( \5498 , \5497 , \5200 );
and \U$5156 ( \5499 , \5496 , \5498 );
xor \U$5157 ( \5500 , \5210 , \5222 );
xor \U$5158 ( \5501 , \5500 , \5229 );
xor \U$5159 ( \5502 , \5094 , \5115 );
xor \U$5160 ( \5503 , \5502 , \5200 );
and \U$5161 ( \5504 , \5501 , \5503 );
and \U$5162 ( \5505 , \5496 , \5501 );
or \U$5163 ( \5506 , \5499 , \5504 , \5505 );
xor \U$5164 ( \5507 , \5495 , \5506 );
xor \U$5165 ( \5508 , \4989 , \4995 );
xor \U$5166 ( \5509 , \5508 , \5006 );
and \U$5167 ( \5510 , \5507 , \5509 );
and \U$5168 ( \5511 , \5495 , \5506 );
or \U$5169 ( \5512 , \5510 , \5511 );
nand \U$5170 ( \5513 , \5265 , \5512 );
nand \U$5171 ( \5514 , \5262 , \5513 );
nand \U$5172 ( \5515 , \5257 , \5514 );
or \U$5173 ( \5516 , \5254 , \5515 );
xnor \U$5174 ( \5517 , \5515 , \5254 );
not \U$5175 ( \5518 , \5261 );
not \U$5176 ( \5519 , \5512 );
or \U$5177 ( \5520 , \5518 , \5519 );
or \U$5178 ( \5521 , \5512 , \5261 );
nand \U$5179 ( \5522 , \5520 , \5521 );
not \U$5180 ( \5523 , \5522 );
not \U$5181 ( \5524 , \5259 );
and \U$5182 ( \5525 , \5523 , \5524 );
and \U$5183 ( \5526 , \5522 , \5259 );
nor \U$5184 ( \5527 , \5525 , \5526 );
not \U$5185 ( \5528 , \5527 );
xor \U$5186 ( \5529 , \5367 , \5453 );
xor \U$5187 ( \5530 , \5529 , \5466 );
xor \U$5188 ( \5531 , \5482 , \5484 );
xor \U$5189 ( \5532 , \5531 , \5489 );
and \U$5190 ( \5533 , \5530 , \5532 );
xor \U$5191 ( \5534 , \5040 , \5063 );
xor \U$5192 ( \5535 , \5534 , \5091 );
xor \U$5193 ( \5536 , \5267 , \5272 );
xor \U$5194 ( \5537 , \5535 , \5536 );
xor \U$5195 ( \5538 , \5482 , \5484 );
xor \U$5196 ( \5539 , \5538 , \5489 );
and \U$5197 ( \5540 , \5537 , \5539 );
and \U$5198 ( \5541 , \5530 , \5537 );
or \U$5199 ( \5542 , \5533 , \5540 , \5541 );
xor \U$5200 ( \5543 , \5303 , \5336 );
xor \U$5201 ( \5544 , \5543 , \5364 );
xor \U$5202 ( \5545 , \5393 , \5422 );
xor \U$5203 ( \5546 , \5545 , \5450 );
and \U$5204 ( \5547 , \5544 , \5546 );
xor \U$5205 ( \5548 , \5123 , \5131 );
xor \U$5206 ( \5549 , \5548 , \5140 );
xor \U$5207 ( \5550 , \5456 , \5461 );
xor \U$5208 ( \5551 , \5549 , \5550 );
xor \U$5209 ( \5552 , \5393 , \5422 );
xor \U$5210 ( \5553 , \5552 , \5450 );
and \U$5211 ( \5554 , \5551 , \5553 );
and \U$5212 ( \5555 , \5544 , \5551 );
or \U$5213 ( \5556 , \5547 , \5554 , \5555 );
not \U$5214 ( \5557 , \3412 );
and \U$5215 ( \5558 , \3683 , RI986df90_7);
and \U$5216 ( \5559 , RI986dea0_5, \3681 );
nor \U$5217 ( \5560 , \5558 , \5559 );
not \U$5218 ( \5561 , \5560 );
or \U$5219 ( \5562 , \5557 , \5561 );
or \U$5220 ( \5563 , \5560 , \3412 );
nand \U$5221 ( \5564 , \5562 , \5563 );
not \U$5222 ( \5565 , \3406 );
and \U$5223 ( \5566 , \3254 , RI986f520_53);
and \U$5224 ( \5567 , RI986f610_55, \3252 );
nor \U$5225 ( \5568 , \5566 , \5567 );
not \U$5226 ( \5569 , \5568 );
or \U$5227 ( \5570 , \5565 , \5569 );
or \U$5228 ( \5571 , \5568 , \3406 );
nand \U$5229 ( \5572 , \5570 , \5571 );
xor \U$5230 ( \5573 , \5564 , \5572 );
and \U$5231 ( \5574 , \4203 , RI986ddb0_3);
and \U$5232 ( \5575 , RI986dcc0_1, \4201 );
nor \U$5233 ( \5576 , \5574 , \5575 );
and \U$5234 ( \5577 , \5576 , \4207 );
not \U$5235 ( \5578 , \5576 );
and \U$5236 ( \5579 , \5578 , \3922 );
nor \U$5237 ( \5580 , \5577 , \5579 );
and \U$5238 ( \5581 , \5573 , \5580 );
and \U$5239 ( \5582 , \5564 , \5572 );
or \U$5240 ( \5583 , \5581 , \5582 );
and \U$5241 ( \5584 , \5318 , RI986e260_13);
and \U$5242 ( \5585 , RI986e350_15, \5316 );
nor \U$5243 ( \5586 , \5584 , \5585 );
and \U$5244 ( \5587 , \5586 , \5052 );
not \U$5245 ( \5588 , \5586 );
and \U$5246 ( \5589 , \5588 , \5322 );
nor \U$5247 ( \5590 , \5587 , \5589 );
not \U$5248 ( \5591 , RI9872a18_166);
not \U$5249 ( \5592 , RI9872a90_167);
or \U$5250 ( \5593 , \5591 , \5592 );
nand \U$5251 ( \5594 , \5593 , RI98729a0_165);
xor \U$5252 ( \5595 , \5590 , \5594 );
not \U$5253 ( \5596 , \4521 );
and \U$5254 ( \5597 , \4710 , RI986e170_11);
and \U$5255 ( \5598 , RI986e080_9, \4708 );
nor \U$5256 ( \5599 , \5597 , \5598 );
not \U$5257 ( \5600 , \5599 );
or \U$5258 ( \5601 , \5596 , \5600 );
or \U$5259 ( \5602 , \5599 , \4521 );
nand \U$5260 ( \5603 , \5601 , \5602 );
and \U$5261 ( \5604 , \5595 , \5603 );
and \U$5262 ( \5605 , \5590 , \5594 );
or \U$5263 ( \5606 , \5604 , \5605 );
xor \U$5264 ( \5607 , \5583 , \5606 );
and \U$5265 ( \5608 , \2274 , RI986f9d0_63);
and \U$5266 ( \5609 , RI986f8e0_61, \2272 );
nor \U$5267 ( \5610 , \5608 , \5609 );
and \U$5268 ( \5611 , \5610 , \2030 );
not \U$5269 ( \5612 , \5610 );
and \U$5270 ( \5613 , \5612 , \2031 );
nor \U$5271 ( \5614 , \5611 , \5613 );
not \U$5272 ( \5615 , \2034 );
and \U$5273 ( \5616 , \2042 , RI986f7f0_59);
and \U$5274 ( \5617 , RI986f700_57, \2040 );
nor \U$5275 ( \5618 , \5616 , \5617 );
not \U$5276 ( \5619 , \5618 );
or \U$5277 ( \5620 , \5615 , \5619 );
or \U$5278 ( \5621 , \5618 , \2034 );
nand \U$5279 ( \5622 , \5620 , \5621 );
xor \U$5280 ( \5623 , \5614 , \5622 );
and \U$5281 ( \5624 , \2464 , RI986f430_51);
and \U$5282 ( \5625 , RI986f340_49, \2462 );
nor \U$5283 ( \5626 , \5624 , \5625 );
and \U$5284 ( \5627 , \5626 , \2468 );
not \U$5285 ( \5628 , \5626 );
and \U$5286 ( \5629 , \5628 , \2263 );
nor \U$5287 ( \5630 , \5627 , \5629 );
and \U$5288 ( \5631 , \5623 , \5630 );
and \U$5289 ( \5632 , \5614 , \5622 );
or \U$5290 ( \5633 , \5631 , \5632 );
and \U$5291 ( \5634 , \5607 , \5633 );
and \U$5292 ( \5635 , \5583 , \5606 );
or \U$5293 ( \5636 , \5634 , \5635 );
nand \U$5294 ( \5637 , RI98716e0_125, RI9871fc8_144);
not \U$5295 ( \5638 , \5401 );
not \U$5296 ( \5639 , \5420 );
or \U$5297 ( \5640 , \5638 , \5639 );
or \U$5298 ( \5641 , \5401 , \5420 );
nand \U$5299 ( \5642 , \5640 , \5641 );
not \U$5300 ( \5643 , \5642 );
not \U$5301 ( \5644 , \5408 );
and \U$5302 ( \5645 , \5643 , \5644 );
and \U$5303 ( \5646 , \5642 , \5408 );
nor \U$5304 ( \5647 , \5645 , \5646 );
nand \U$5305 ( \5648 , \5637 , \5647 );
xor \U$5306 ( \5649 , \5636 , \5648 );
not \U$5307 ( \5650 , \454 );
and \U$5308 ( \5651 , \465 , RI986ee90_39);
and \U$5309 ( \5652 , RI986eda0_37, \463 );
nor \U$5310 ( \5653 , \5651 , \5652 );
not \U$5311 ( \5654 , \5653 );
or \U$5312 ( \5655 , \5650 , \5654 );
or \U$5313 ( \5656 , \5653 , \456 );
nand \U$5314 ( \5657 , \5655 , \5656 );
and \U$5315 ( \5658 , \776 , RI986f070_43);
and \U$5316 ( \5659 , RI986ef80_41, \774 );
nor \U$5317 ( \5660 , \5658 , \5659 );
and \U$5318 ( \5661 , \5660 , \474 );
not \U$5319 ( \5662 , \5660 );
and \U$5320 ( \5663 , \5662 , \451 );
nor \U$5321 ( \5664 , \5661 , \5663 );
xor \U$5322 ( \5665 , \5657 , \5664 );
and \U$5323 ( \5666 , \438 , RI986ebc0_33);
and \U$5324 ( \5667 , RI986ecb0_35, \436 );
nor \U$5325 ( \5668 , \5666 , \5667 );
and \U$5326 ( \5669 , \5668 , \444 );
not \U$5327 ( \5670 , \5668 );
and \U$5328 ( \5671 , \5670 , \443 );
nor \U$5329 ( \5672 , \5669 , \5671 );
and \U$5330 ( \5673 , \5665 , \5672 );
and \U$5331 ( \5674 , \5657 , \5664 );
or \U$5332 ( \5675 , \5673 , \5674 );
not \U$5333 ( \5676 , \367 );
and \U$5334 ( \5677 , \376 , RI986e8f0_27);
and \U$5335 ( \5678 , RI986e800_25, \374 );
nor \U$5336 ( \5679 , \5677 , \5678 );
not \U$5337 ( \5680 , \5679 );
or \U$5338 ( \5681 , \5676 , \5680 );
or \U$5339 ( \5682 , \5679 , \367 );
nand \U$5340 ( \5683 , \5681 , \5682 );
not \U$5341 ( \5684 , \386 );
and \U$5342 ( \5685 , \395 , RI986ead0_31);
and \U$5343 ( \5686 , RI986e9e0_29, \393 );
nor \U$5344 ( \5687 , \5685 , \5686 );
not \U$5345 ( \5688 , \5687 );
or \U$5346 ( \5689 , \5684 , \5688 );
or \U$5347 ( \5690 , \5687 , \386 );
nand \U$5348 ( \5691 , \5689 , \5690 );
xor \U$5349 ( \5692 , \5683 , \5691 );
not \U$5350 ( \5693 , \361 );
and \U$5351 ( \5694 , \354 , RI9871500_121);
and \U$5352 ( \5695 , RI98715f0_123, \352 );
nor \U$5353 ( \5696 , \5694 , \5695 );
not \U$5354 ( \5697 , \5696 );
or \U$5355 ( \5698 , \5693 , \5697 );
or \U$5356 ( \5699 , \5696 , \345 );
nand \U$5357 ( \5700 , \5698 , \5699 );
and \U$5358 ( \5701 , \5692 , \5700 );
and \U$5359 ( \5702 , \5683 , \5691 );
or \U$5360 ( \5703 , \5701 , \5702 );
xor \U$5361 ( \5704 , \5675 , \5703 );
and \U$5362 ( \5705 , \1311 , RI986e710_23);
and \U$5363 ( \5706 , RI986e620_21, \1309 );
nor \U$5364 ( \5707 , \5705 , \5706 );
and \U$5365 ( \5708 , \5707 , \1458 );
not \U$5366 ( \5709 , \5707 );
and \U$5367 ( \5710 , \5709 , \1318 );
nor \U$5368 ( \5711 , \5708 , \5710 );
not \U$5369 ( \5712 , \1128 );
and \U$5370 ( \5713 , \1293 , RI986f250_47);
and \U$5371 ( \5714 , RI986f160_45, \1291 );
nor \U$5372 ( \5715 , \5713 , \5714 );
not \U$5373 ( \5716 , \5715 );
or \U$5374 ( \5717 , \5712 , \5716 );
or \U$5375 ( \5718 , \5715 , \1301 );
nand \U$5376 ( \5719 , \5717 , \5718 );
xor \U$5377 ( \5720 , \5711 , \5719 );
and \U$5378 ( \5721 , \1329 , RI986e530_19);
and \U$5379 ( \5722 , RI986e440_17, \1327 );
nor \U$5380 ( \5723 , \5721 , \5722 );
and \U$5381 ( \5724 , \5723 , \1336 );
not \U$5382 ( \5725 , \5723 );
and \U$5383 ( \5726 , \5725 , \1337 );
nor \U$5384 ( \5727 , \5724 , \5726 );
and \U$5385 ( \5728 , \5720 , \5727 );
and \U$5386 ( \5729 , \5711 , \5719 );
or \U$5387 ( \5730 , \5728 , \5729 );
and \U$5388 ( \5731 , \5704 , \5730 );
and \U$5389 ( \5732 , \5675 , \5703 );
or \U$5390 ( \5733 , \5731 , \5732 );
and \U$5391 ( \5734 , \5649 , \5733 );
and \U$5392 ( \5735 , \5636 , \5648 );
or \U$5393 ( \5736 , \5734 , \5735 );
xor \U$5394 ( \5737 , \5556 , \5736 );
xor \U$5395 ( \5738 , \5431 , \5438 );
xor \U$5396 ( \5739 , \5738 , \5447 );
xor \U$5397 ( \5740 , \5285 , \5292 );
xor \U$5398 ( \5741 , \5740 , \5300 );
and \U$5399 ( \5742 , \5739 , \5741 );
xor \U$5400 ( \5743 , \5375 , \5382 );
xor \U$5401 ( \5744 , \5743 , \5390 );
xor \U$5402 ( \5745 , \5285 , \5292 );
xor \U$5403 ( \5746 , \5745 , \5300 );
and \U$5404 ( \5747 , \5744 , \5746 );
and \U$5405 ( \5748 , \5739 , \5744 );
or \U$5406 ( \5749 , \5742 , \5747 , \5748 );
xor \U$5407 ( \5750 , \5048 , \5052 );
xor \U$5408 ( \5751 , \5750 , \5060 );
xor \U$5409 ( \5752 , \5749 , \5751 );
xor \U$5410 ( \5753 , \5072 , \5079 );
xor \U$5411 ( \5754 , \5753 , \5088 );
xor \U$5412 ( \5755 , \5472 , \5477 );
xor \U$5413 ( \5756 , \5754 , \5755 );
and \U$5414 ( \5757 , \5752 , \5756 );
and \U$5415 ( \5758 , \5749 , \5751 );
or \U$5416 ( \5759 , \5757 , \5758 );
and \U$5417 ( \5760 , \5737 , \5759 );
and \U$5418 ( \5761 , \5556 , \5736 );
or \U$5419 ( \5762 , \5760 , \5761 );
xor \U$5420 ( \5763 , \5542 , \5762 );
xor \U$5421 ( \5764 , \5094 , \5115 );
xor \U$5422 ( \5765 , \5764 , \5200 );
xor \U$5423 ( \5766 , \5496 , \5501 );
xor \U$5424 ( \5767 , \5765 , \5766 );
and \U$5425 ( \5768 , \5763 , \5767 );
and \U$5426 ( \5769 , \5542 , \5762 );
or \U$5427 ( \5770 , \5768 , \5769 );
xor \U$5428 ( \5771 , \5014 , \5203 );
xor \U$5429 ( \5772 , \5771 , \5232 );
xor \U$5430 ( \5773 , \5770 , \5772 );
xor \U$5431 ( \5774 , \5495 , \5506 );
xor \U$5432 ( \5775 , \5774 , \5509 );
and \U$5433 ( \5776 , \5773 , \5775 );
and \U$5434 ( \5777 , \5770 , \5772 );
or \U$5435 ( \5778 , \5776 , \5777 );
not \U$5436 ( \5779 , \5778 );
and \U$5437 ( \5780 , \5528 , \5779 );
and \U$5438 ( \5781 , \5527 , \5778 );
nor \U$5439 ( \5782 , \5780 , \5781 );
xor \U$5440 ( \5783 , \5636 , \5648 );
xor \U$5441 ( \5784 , \5783 , \5733 );
xor \U$5442 ( \5785 , \5749 , \5751 );
xor \U$5443 ( \5786 , \5785 , \5756 );
and \U$5444 ( \5787 , \5784 , \5786 );
xor \U$5445 ( \5788 , \5393 , \5422 );
xor \U$5446 ( \5789 , \5788 , \5450 );
xor \U$5447 ( \5790 , \5544 , \5551 );
xor \U$5448 ( \5791 , \5789 , \5790 );
xor \U$5449 ( \5792 , \5749 , \5751 );
xor \U$5450 ( \5793 , \5792 , \5756 );
and \U$5451 ( \5794 , \5791 , \5793 );
and \U$5452 ( \5795 , \5784 , \5791 );
or \U$5453 ( \5796 , \5787 , \5794 , \5795 );
xor \U$5454 ( \5797 , \5683 , \5691 );
xor \U$5455 ( \5798 , \5797 , \5700 );
xor \U$5456 ( \5799 , \5657 , \5664 );
xor \U$5457 ( \5800 , \5799 , \5672 );
and \U$5458 ( \5801 , \5798 , \5800 );
xor \U$5459 ( \5802 , \5711 , \5719 );
xor \U$5460 ( \5803 , \5802 , \5727 );
xor \U$5461 ( \5804 , \5657 , \5664 );
xor \U$5462 ( \5805 , \5804 , \5672 );
and \U$5463 ( \5806 , \5803 , \5805 );
and \U$5464 ( \5807 , \5798 , \5803 );
or \U$5465 ( \5808 , \5801 , \5806 , \5807 );
xor \U$5466 ( \5809 , \5345 , \5352 );
xor \U$5467 ( \5810 , \5809 , \5361 );
xor \U$5468 ( \5811 , \5808 , \5810 );
xor \U$5469 ( \5812 , \5590 , \5594 );
xor \U$5470 ( \5813 , \5812 , \5603 );
xor \U$5471 ( \5814 , \5564 , \5572 );
xor \U$5472 ( \5815 , \5814 , \5580 );
and \U$5473 ( \5816 , \5813 , \5815 );
xor \U$5474 ( \5817 , \5614 , \5622 );
xor \U$5475 ( \5818 , \5817 , \5630 );
xor \U$5476 ( \5819 , \5564 , \5572 );
xor \U$5477 ( \5820 , \5819 , \5580 );
and \U$5478 ( \5821 , \5818 , \5820 );
and \U$5479 ( \5822 , \5813 , \5818 );
or \U$5480 ( \5823 , \5816 , \5821 , \5822 );
and \U$5481 ( \5824 , \5811 , \5823 );
and \U$5482 ( \5825 , \5808 , \5810 );
or \U$5483 ( \5826 , \5824 , \5825 );
and \U$5484 ( \5827 , \2042 , RI986e620_21);
and \U$5485 ( \5828 , RI986f7f0_59, \2040 );
nor \U$5486 ( \5829 , \5827 , \5828 );
not \U$5487 ( \5830 , \5829 );
not \U$5488 ( \5831 , \2034 );
and \U$5489 ( \5832 , \5830 , \5831 );
and \U$5490 ( \5833 , \5829 , \2034 );
nor \U$5491 ( \5834 , \5832 , \5833 );
and \U$5492 ( \5835 , \2464 , RI986f8e0_61);
and \U$5493 ( \5836 , RI986f430_51, \2462 );
nor \U$5494 ( \5837 , \5835 , \5836 );
and \U$5495 ( \5838 , \5837 , \2263 );
not \U$5496 ( \5839 , \5837 );
and \U$5497 ( \5840 , \5839 , \2468 );
nor \U$5498 ( \5841 , \5838 , \5840 );
or \U$5499 ( \5842 , \5834 , \5841 );
not \U$5500 ( \5843 , \5841 );
not \U$5501 ( \5844 , \5834 );
or \U$5502 ( \5845 , \5843 , \5844 );
and \U$5503 ( \5846 , \2274 , RI986f700_57);
and \U$5504 ( \5847 , RI986f9d0_63, \2272 );
nor \U$5505 ( \5848 , \5846 , \5847 );
and \U$5506 ( \5849 , \5848 , \2030 );
not \U$5507 ( \5850 , \5848 );
and \U$5508 ( \5851 , \5850 , \2031 );
nor \U$5509 ( \5852 , \5849 , \5851 );
nand \U$5510 ( \5853 , \5845 , \5852 );
nand \U$5511 ( \5854 , \5842 , \5853 );
and \U$5512 ( \5855 , \4710 , RI986dcc0_1);
and \U$5513 ( \5856 , RI986e170_11, \4708 );
nor \U$5514 ( \5857 , \5855 , \5856 );
not \U$5515 ( \5858 , \5857 );
not \U$5516 ( \5859 , \4519 );
and \U$5517 ( \5860 , \5858 , \5859 );
and \U$5518 ( \5861 , \5857 , \4521 );
nor \U$5519 ( \5862 , \5860 , \5861 );
and \U$5520 ( \5863 , \5318 , RI986e080_9);
and \U$5521 ( \5864 , RI986e260_13, \5316 );
nor \U$5522 ( \5865 , \5863 , \5864 );
and \U$5523 ( \5866 , \5865 , \5322 );
not \U$5524 ( \5867 , \5865 );
and \U$5525 ( \5868 , \5867 , \5052 );
nor \U$5526 ( \5869 , \5866 , \5868 );
or \U$5527 ( \5870 , \5862 , \5869 );
not \U$5528 ( \5871 , \5869 );
not \U$5529 ( \5872 , \5862 );
or \U$5530 ( \5873 , \5871 , \5872 );
and \U$5531 ( \5874 , RI98729a0_165, RI9872a90_167);
not \U$5532 ( \5875 , RI9872a18_166);
and \U$5533 ( \5876 , RI9872a90_167, \5875 );
not \U$5534 ( \5877 , RI9872a90_167);
and \U$5535 ( \5878 , \5877 , RI9872a18_166);
or \U$5536 ( \5879 , \5876 , \5878 );
nor \U$5537 ( \5880 , RI98729a0_165, RI9872a90_167);
nor \U$5538 ( \5881 , \5874 , \5879 , \5880 );
nand \U$5539 ( \5882 , RI986e350_15, \5881 );
and \U$5540 ( \5883 , \5882 , \5594 );
not \U$5541 ( \5884 , \5882 );
not \U$5542 ( \5885 , \5594 );
and \U$5543 ( \5886 , \5884 , \5885 );
nor \U$5544 ( \5887 , \5883 , \5886 );
nand \U$5545 ( \5888 , \5873 , \5887 );
nand \U$5546 ( \5889 , \5870 , \5888 );
xor \U$5547 ( \5890 , \5854 , \5889 );
not \U$5548 ( \5891 , \3918 );
and \U$5549 ( \5892 , \3683 , RI986f610_55);
and \U$5550 ( \5893 , RI986df90_7, \3681 );
nor \U$5551 ( \5894 , \5892 , \5893 );
not \U$5552 ( \5895 , \5894 );
or \U$5553 ( \5896 , \5891 , \5895 );
or \U$5554 ( \5897 , \5894 , \3412 );
nand \U$5555 ( \5898 , \5896 , \5897 );
not \U$5556 ( \5899 , \2935 );
and \U$5557 ( \5900 , \3254 , RI986f340_49);
and \U$5558 ( \5901 , RI986f520_53, \3252 );
nor \U$5559 ( \5902 , \5900 , \5901 );
not \U$5560 ( \5903 , \5902 );
or \U$5561 ( \5904 , \5899 , \5903 );
or \U$5562 ( \5905 , \5902 , \2935 );
nand \U$5563 ( \5906 , \5904 , \5905 );
xor \U$5564 ( \5907 , \5898 , \5906 );
and \U$5565 ( \5908 , \4203 , RI986dea0_5);
and \U$5566 ( \5909 , RI986ddb0_3, \4201 );
nor \U$5567 ( \5910 , \5908 , \5909 );
and \U$5568 ( \5911 , \5910 , \4207 );
not \U$5569 ( \5912 , \5910 );
and \U$5570 ( \5913 , \5912 , \3923 );
nor \U$5571 ( \5914 , \5911 , \5913 );
and \U$5572 ( \5915 , \5907 , \5914 );
and \U$5573 ( \5916 , \5898 , \5906 );
or \U$5574 ( \5917 , \5915 , \5916 );
and \U$5575 ( \5918 , \5890 , \5917 );
and \U$5576 ( \5919 , \5854 , \5889 );
or \U$5577 ( \5920 , \5918 , \5919 );
and \U$5578 ( \5921 , \416 , RI98716e0_125);
and \U$5579 ( \5922 , RI98717d0_127, \414 );
nor \U$5580 ( \5923 , \5921 , \5922 );
and \U$5581 ( \5924 , \5923 , \422 );
not \U$5582 ( \5925 , \5923 );
and \U$5583 ( \5926 , \5925 , \421 );
nor \U$5584 ( \5927 , \5924 , \5926 );
not \U$5585 ( \5928 , RI9871410_119);
nor \U$5586 ( \5929 , \5928 , \407 );
xor \U$5587 ( \5930 , \5927 , \5929 );
nand \U$5588 ( \5931 , RI9871320_117, RI9871fc8_144);
and \U$5589 ( \5932 , \416 , RI9871410_119);
and \U$5590 ( \5933 , RI98716e0_125, \414 );
nor \U$5591 ( \5934 , \5932 , \5933 );
and \U$5592 ( \5935 , \5934 , \421 );
not \U$5593 ( \5936 , \5934 );
and \U$5594 ( \5937 , \5936 , \422 );
nor \U$5595 ( \5938 , \5935 , \5937 );
nand \U$5596 ( \5939 , \5931 , \5938 );
and \U$5597 ( \5940 , \5930 , \5939 );
and \U$5598 ( \5941 , \5927 , \5929 );
or \U$5599 ( \5942 , \5940 , \5941 );
xor \U$5600 ( \5943 , \5920 , \5942 );
not \U$5601 ( \5944 , \361 );
and \U$5602 ( \5945 , \354 , RI98717d0_127);
and \U$5603 ( \5946 , RI9871500_121, \352 );
nor \U$5604 ( \5947 , \5945 , \5946 );
not \U$5605 ( \5948 , \5947 );
or \U$5606 ( \5949 , \5944 , \5948 );
or \U$5607 ( \5950 , \5947 , \361 );
nand \U$5608 ( \5951 , \5949 , \5950 );
not \U$5609 ( \5952 , \365 );
and \U$5610 ( \5953 , \376 , RI986e9e0_29);
and \U$5611 ( \5954 , RI986e8f0_27, \374 );
nor \U$5612 ( \5955 , \5953 , \5954 );
not \U$5613 ( \5956 , \5955 );
or \U$5614 ( \5957 , \5952 , \5956 );
or \U$5615 ( \5958 , \5955 , \365 );
nand \U$5616 ( \5959 , \5957 , \5958 );
xor \U$5617 ( \5960 , \5951 , \5959 );
not \U$5618 ( \5961 , \386 );
and \U$5619 ( \5962 , \395 , RI98715f0_123);
and \U$5620 ( \5963 , RI986ead0_31, \393 );
nor \U$5621 ( \5964 , \5962 , \5963 );
not \U$5622 ( \5965 , \5964 );
or \U$5623 ( \5966 , \5961 , \5965 );
or \U$5624 ( \5967 , \5964 , \487 );
nand \U$5625 ( \5968 , \5966 , \5967 );
and \U$5626 ( \5969 , \5960 , \5968 );
and \U$5627 ( \5970 , \5951 , \5959 );
or \U$5628 ( \5971 , \5969 , \5970 );
and \U$5629 ( \5972 , \776 , RI986ecb0_35);
and \U$5630 ( \5973 , RI986f070_43, \774 );
nor \U$5631 ( \5974 , \5972 , \5973 );
and \U$5632 ( \5975 , \5974 , \451 );
not \U$5633 ( \5976 , \5974 );
and \U$5634 ( \5977 , \5976 , \474 );
nor \U$5635 ( \5978 , \5975 , \5977 );
and \U$5636 ( \5979 , \438 , RI986eda0_37);
and \U$5637 ( \5980 , RI986ebc0_33, \436 );
nor \U$5638 ( \5981 , \5979 , \5980 );
and \U$5639 ( \5982 , \5981 , \443 );
not \U$5640 ( \5983 , \5981 );
and \U$5641 ( \5984 , \5983 , \444 );
nor \U$5642 ( \5985 , \5982 , \5984 );
xor \U$5643 ( \5986 , \5978 , \5985 );
and \U$5644 ( \5987 , \465 , RI986e800_25);
and \U$5645 ( \5988 , RI986ee90_39, \463 );
nor \U$5646 ( \5989 , \5987 , \5988 );
not \U$5647 ( \5990 , \5989 );
not \U$5648 ( \5991 , \454 );
and \U$5649 ( \5992 , \5990 , \5991 );
and \U$5650 ( \5993 , \5989 , \454 );
nor \U$5651 ( \5994 , \5992 , \5993 );
and \U$5652 ( \5995 , \5986 , \5994 );
and \U$5653 ( \5996 , \5978 , \5985 );
nor \U$5654 ( \5997 , \5995 , \5996 );
xor \U$5655 ( \5998 , \5971 , \5997 );
and \U$5656 ( \5999 , \1329 , RI986f160_45);
and \U$5657 ( \6000 , RI986e530_19, \1327 );
nor \U$5658 ( \6001 , \5999 , \6000 );
and \U$5659 ( \6002 , \6001 , \1337 );
not \U$5660 ( \6003 , \6001 );
and \U$5661 ( \6004 , \6003 , \1336 );
nor \U$5662 ( \6005 , \6002 , \6004 );
and \U$5663 ( \6006 , \1311 , RI986e440_17);
and \U$5664 ( \6007 , RI986e710_23, \1309 );
nor \U$5665 ( \6008 , \6006 , \6007 );
and \U$5666 ( \6009 , \6008 , \1315 );
not \U$5667 ( \6010 , \6008 );
and \U$5668 ( \6011 , \6010 , \1458 );
nor \U$5669 ( \6012 , \6009 , \6011 );
xor \U$5670 ( \6013 , \6005 , \6012 );
and \U$5671 ( \6014 , \1293 , RI986ef80_41);
and \U$5672 ( \6015 , RI986f250_47, \1291 );
nor \U$5673 ( \6016 , \6014 , \6015 );
not \U$5674 ( \6017 , \6016 );
not \U$5675 ( \6018 , \1301 );
and \U$5676 ( \6019 , \6017 , \6018 );
and \U$5677 ( \6020 , \6016 , \1301 );
nor \U$5678 ( \6021 , \6019 , \6020 );
and \U$5679 ( \6022 , \6013 , \6021 );
and \U$5680 ( \6023 , \6005 , \6012 );
nor \U$5681 ( \6024 , \6022 , \6023 );
and \U$5682 ( \6025 , \5998 , \6024 );
and \U$5683 ( \6026 , \5971 , \5997 );
or \U$5684 ( \6027 , \6025 , \6026 );
and \U$5685 ( \6028 , \5943 , \6027 );
and \U$5686 ( \6029 , \5920 , \5942 );
or \U$5687 ( \6030 , \6028 , \6029 );
xor \U$5688 ( \6031 , \5826 , \6030 );
or \U$5689 ( \6032 , \5647 , \5637 );
nand \U$5690 ( \6033 , \6032 , \5648 );
xor \U$5691 ( \6034 , \5310 , \5324 );
xor \U$5692 ( \6035 , \6034 , \5333 );
xor \U$5693 ( \6036 , \6033 , \6035 );
xor \U$5694 ( \6037 , \5285 , \5292 );
xor \U$5695 ( \6038 , \6037 , \5300 );
xor \U$5696 ( \6039 , \5739 , \5744 );
xor \U$5697 ( \6040 , \6038 , \6039 );
and \U$5698 ( \6041 , \6036 , \6040 );
and \U$5699 ( \6042 , \6033 , \6035 );
or \U$5700 ( \6043 , \6041 , \6042 );
and \U$5701 ( \6044 , \6031 , \6043 );
and \U$5702 ( \6045 , \5826 , \6030 );
or \U$5703 ( \6046 , \6044 , \6045 );
xor \U$5704 ( \6047 , \5796 , \6046 );
xor \U$5705 ( \6048 , \5482 , \5484 );
xor \U$5706 ( \6049 , \6048 , \5489 );
xor \U$5707 ( \6050 , \5530 , \5537 );
xor \U$5708 ( \6051 , \6049 , \6050 );
and \U$5709 ( \6052 , \6047 , \6051 );
and \U$5710 ( \6053 , \5796 , \6046 );
or \U$5711 ( \6054 , \6052 , \6053 );
xor \U$5712 ( \6055 , \5277 , \5469 );
xor \U$5713 ( \6056 , \6055 , \5492 );
xor \U$5714 ( \6057 , \6054 , \6056 );
xor \U$5715 ( \6058 , \5542 , \5762 );
xor \U$5716 ( \6059 , \6058 , \5767 );
and \U$5717 ( \6060 , \6057 , \6059 );
and \U$5718 ( \6061 , \6054 , \6056 );
or \U$5719 ( \6062 , \6060 , \6061 );
xor \U$5720 ( \6063 , \5770 , \5772 );
xor \U$5721 ( \6064 , \6063 , \5775 );
nand \U$5722 ( \6065 , \6062 , \6064 );
or \U$5723 ( \6066 , \5782 , \6065 );
xnor \U$5724 ( \6067 , \6065 , \5782 );
xor \U$5725 ( \6068 , \6062 , \6064 );
xor \U$5726 ( \6069 , \5927 , \5929 );
xor \U$5727 ( \6070 , \6069 , \5939 );
xor \U$5728 ( \6071 , \5971 , \5997 );
xor \U$5729 ( \6072 , \6071 , \6024 );
and \U$5730 ( \6073 , \6070 , \6072 );
xor \U$5731 ( \6074 , \5657 , \5664 );
xor \U$5732 ( \6075 , \6074 , \5672 );
xor \U$5733 ( \6076 , \5798 , \5803 );
xor \U$5734 ( \6077 , \6075 , \6076 );
xor \U$5735 ( \6078 , \5971 , \5997 );
xor \U$5736 ( \6079 , \6078 , \6024 );
and \U$5737 ( \6080 , \6077 , \6079 );
and \U$5738 ( \6081 , \6070 , \6077 );
or \U$5739 ( \6082 , \6073 , \6080 , \6081 );
and \U$5740 ( \6083 , \776 , RI986ebc0_33);
and \U$5741 ( \6084 , RI986ecb0_35, \774 );
nor \U$5742 ( \6085 , \6083 , \6084 );
and \U$5743 ( \6086 , \6085 , \451 );
not \U$5744 ( \6087 , \6085 );
and \U$5745 ( \6088 , \6087 , \474 );
nor \U$5746 ( \6089 , \6086 , \6088 );
not \U$5747 ( \6090 , \6089 );
and \U$5748 ( \6091 , \438 , RI986ee90_39);
and \U$5749 ( \6092 , RI986eda0_37, \436 );
nor \U$5750 ( \6093 , \6091 , \6092 );
and \U$5751 ( \6094 , \6093 , \443 );
not \U$5752 ( \6095 , \6093 );
and \U$5753 ( \6096 , \6095 , \444 );
nor \U$5754 ( \6097 , \6094 , \6096 );
not \U$5755 ( \6098 , \6097 );
and \U$5756 ( \6099 , \6090 , \6098 );
and \U$5757 ( \6100 , \6097 , \6089 );
and \U$5758 ( \6101 , \1293 , RI986f070_43);
and \U$5759 ( \6102 , RI986ef80_41, \1291 );
nor \U$5760 ( \6103 , \6101 , \6102 );
not \U$5761 ( \6104 , \6103 );
not \U$5762 ( \6105 , \1301 );
and \U$5763 ( \6106 , \6104 , \6105 );
and \U$5764 ( \6107 , \6103 , \1128 );
nor \U$5765 ( \6108 , \6106 , \6107 );
nor \U$5766 ( \6109 , \6100 , \6108 );
nor \U$5767 ( \6110 , \6099 , \6109 );
and \U$5768 ( \6111 , \1329 , RI986f250_47);
and \U$5769 ( \6112 , RI986f160_45, \1327 );
nor \U$5770 ( \6113 , \6111 , \6112 );
and \U$5771 ( \6114 , \6113 , \1337 );
not \U$5772 ( \6115 , \6113 );
and \U$5773 ( \6116 , \6115 , \1336 );
nor \U$5774 ( \6117 , \6114 , \6116 );
not \U$5775 ( \6118 , \6117 );
and \U$5776 ( \6119 , \1311 , RI986e530_19);
and \U$5777 ( \6120 , RI986e440_17, \1309 );
nor \U$5778 ( \6121 , \6119 , \6120 );
and \U$5779 ( \6122 , \6121 , \1318 );
not \U$5780 ( \6123 , \6121 );
and \U$5781 ( \6124 , \6123 , \1458 );
nor \U$5782 ( \6125 , \6122 , \6124 );
not \U$5783 ( \6126 , \6125 );
and \U$5784 ( \6127 , \6118 , \6126 );
and \U$5785 ( \6128 , \6125 , \6117 );
and \U$5786 ( \6129 , \2042 , RI986e710_23);
and \U$5787 ( \6130 , RI986e620_21, \2040 );
nor \U$5788 ( \6131 , \6129 , \6130 );
not \U$5789 ( \6132 , \6131 );
not \U$5790 ( \6133 , \2034 );
and \U$5791 ( \6134 , \6132 , \6133 );
and \U$5792 ( \6135 , \6131 , \2034 );
nor \U$5793 ( \6136 , \6134 , \6135 );
nor \U$5794 ( \6137 , \6128 , \6136 );
nor \U$5795 ( \6138 , \6127 , \6137 );
xor \U$5796 ( \6139 , \6110 , \6138 );
and \U$5797 ( \6140 , \465 , RI986e8f0_27);
and \U$5798 ( \6141 , RI986e800_25, \463 );
nor \U$5799 ( \6142 , \6140 , \6141 );
not \U$5800 ( \6143 , \6142 );
not \U$5801 ( \6144 , \456 );
and \U$5802 ( \6145 , \6143 , \6144 );
and \U$5803 ( \6146 , \6142 , \456 );
nor \U$5804 ( \6147 , \6145 , \6146 );
and \U$5805 ( \6148 , \376 , RI986ead0_31);
and \U$5806 ( \6149 , RI986e9e0_29, \374 );
nor \U$5807 ( \6150 , \6148 , \6149 );
not \U$5808 ( \6151 , \6150 );
not \U$5809 ( \6152 , \365 );
and \U$5810 ( \6153 , \6151 , \6152 );
and \U$5811 ( \6154 , \6150 , \365 );
nor \U$5812 ( \6155 , \6153 , \6154 );
xor \U$5813 ( \6156 , \6147 , \6155 );
and \U$5814 ( \6157 , \395 , RI9871500_121);
and \U$5815 ( \6158 , RI98715f0_123, \393 );
nor \U$5816 ( \6159 , \6157 , \6158 );
not \U$5817 ( \6160 , \6159 );
not \U$5818 ( \6161 , \487 );
and \U$5819 ( \6162 , \6160 , \6161 );
and \U$5820 ( \6163 , \6159 , \487 );
nor \U$5821 ( \6164 , \6162 , \6163 );
and \U$5822 ( \6165 , \6156 , \6164 );
and \U$5823 ( \6166 , \6147 , \6155 );
or \U$5824 ( \6167 , \6165 , \6166 );
and \U$5825 ( \6168 , \6139 , \6167 );
and \U$5826 ( \6169 , \6110 , \6138 );
nor \U$5827 ( \6170 , \6168 , \6169 );
and \U$5828 ( \6171 , \5881 , RI986e260_13);
and \U$5829 ( \6172 , RI986e350_15, \5879 );
nor \U$5830 ( \6173 , \6171 , \6172 );
and \U$5831 ( \6174 , \6173 , \5594 );
not \U$5832 ( \6175 , \6173 );
and \U$5833 ( \6176 , \6175 , \5885 );
nor \U$5834 ( \6177 , \6174 , \6176 );
not \U$5835 ( \6178 , \6177 );
and \U$5836 ( \6179 , RI9872b08_168, RI9872b80_169);
nor \U$5837 ( \6180 , \6179 , \5875 );
nand \U$5838 ( \6181 , \6178 , \6180 );
and \U$5839 ( \6182 , \5318 , RI986e170_11);
and \U$5840 ( \6183 , RI986e080_9, \5316 );
nor \U$5841 ( \6184 , \6182 , \6183 );
and \U$5842 ( \6185 , \6184 , \5052 );
not \U$5843 ( \6186 , \6184 );
and \U$5844 ( \6187 , \6186 , \5322 );
nor \U$5845 ( \6188 , \6185 , \6187 );
and \U$5846 ( \6189 , \6181 , \6188 );
not \U$5847 ( \6190 , \6180 );
and \U$5848 ( \6191 , \6190 , \6177 );
nor \U$5849 ( \6192 , \6189 , \6191 );
and \U$5850 ( \6193 , \3683 , RI986f520_53);
and \U$5851 ( \6194 , RI986f610_55, \3681 );
nor \U$5852 ( \6195 , \6193 , \6194 );
not \U$5853 ( \6196 , \6195 );
not \U$5854 ( \6197 , \3918 );
and \U$5855 ( \6198 , \6196 , \6197 );
and \U$5856 ( \6199 , \6195 , \3412 );
nor \U$5857 ( \6200 , \6198 , \6199 );
not \U$5858 ( \6201 , \6200 );
and \U$5859 ( \6202 , \4203 , RI986df90_7);
and \U$5860 ( \6203 , RI986dea0_5, \4201 );
nor \U$5861 ( \6204 , \6202 , \6203 );
and \U$5862 ( \6205 , \6204 , \3923 );
not \U$5863 ( \6206 , \6204 );
and \U$5864 ( \6207 , \6206 , \4207 );
nor \U$5865 ( \6208 , \6205 , \6207 );
not \U$5866 ( \6209 , \6208 );
and \U$5867 ( \6210 , \6201 , \6209 );
and \U$5868 ( \6211 , \6208 , \6200 );
and \U$5869 ( \6212 , \4710 , RI986ddb0_3);
and \U$5870 ( \6213 , RI986dcc0_1, \4708 );
nor \U$5871 ( \6214 , \6212 , \6213 );
not \U$5872 ( \6215 , \6214 );
not \U$5873 ( \6216 , \4519 );
and \U$5874 ( \6217 , \6215 , \6216 );
and \U$5875 ( \6218 , \6214 , \4519 );
nor \U$5876 ( \6219 , \6217 , \6218 );
nor \U$5877 ( \6220 , \6211 , \6219 );
nor \U$5878 ( \6221 , \6210 , \6220 );
xor \U$5879 ( \6222 , \6192 , \6221 );
and \U$5880 ( \6223 , \2274 , RI986f7f0_59);
and \U$5881 ( \6224 , RI986f700_57, \2272 );
nor \U$5882 ( \6225 , \6223 , \6224 );
and \U$5883 ( \6226 , \6225 , \2031 );
not \U$5884 ( \6227 , \6225 );
and \U$5885 ( \6228 , \6227 , \2030 );
nor \U$5886 ( \6229 , \6226 , \6228 );
not \U$5887 ( \6230 , \6229 );
and \U$5888 ( \6231 , \2464 , RI986f9d0_63);
and \U$5889 ( \6232 , RI986f8e0_61, \2462 );
nor \U$5890 ( \6233 , \6231 , \6232 );
and \U$5891 ( \6234 , \6233 , \2263 );
not \U$5892 ( \6235 , \6233 );
and \U$5893 ( \6236 , \6235 , \2468 );
nor \U$5894 ( \6237 , \6234 , \6236 );
not \U$5895 ( \6238 , \6237 );
and \U$5896 ( \6239 , \6230 , \6238 );
and \U$5897 ( \6240 , \6237 , \6229 );
and \U$5898 ( \6241 , \3254 , RI986f430_51);
and \U$5899 ( \6242 , RI986f340_49, \3252 );
nor \U$5900 ( \6243 , \6241 , \6242 );
not \U$5901 ( \6244 , \6243 );
not \U$5902 ( \6245 , \3406 );
and \U$5903 ( \6246 , \6244 , \6245 );
and \U$5904 ( \6247 , \6243 , \2935 );
nor \U$5905 ( \6248 , \6246 , \6247 );
nor \U$5906 ( \6249 , \6240 , \6248 );
nor \U$5907 ( \6250 , \6239 , \6249 );
and \U$5908 ( \6251 , \6222 , \6250 );
and \U$5909 ( \6252 , \6192 , \6221 );
nor \U$5910 ( \6253 , \6251 , \6252 );
xor \U$5911 ( \6254 , \6170 , \6253 );
and \U$5912 ( \6255 , \416 , RI9871320_117);
and \U$5913 ( \6256 , RI9871410_119, \414 );
nor \U$5914 ( \6257 , \6255 , \6256 );
and \U$5915 ( \6258 , \6257 , \421 );
not \U$5916 ( \6259 , \6257 );
and \U$5917 ( \6260 , \6259 , \422 );
nor \U$5918 ( \6261 , \6258 , \6260 );
nand \U$5919 ( \6262 , RI9871140_113, RI9871fc8_144);
or \U$5920 ( \6263 , \6261 , \6262 );
not \U$5921 ( \6264 , \6262 );
not \U$5922 ( \6265 , \6261 );
or \U$5923 ( \6266 , \6264 , \6265 );
not \U$5924 ( \6267 , \361 );
and \U$5925 ( \6268 , \354 , RI98716e0_125);
and \U$5926 ( \6269 , RI98717d0_127, \352 );
nor \U$5927 ( \6270 , \6268 , \6269 );
not \U$5928 ( \6271 , \6270 );
or \U$5929 ( \6272 , \6267 , \6271 );
or \U$5930 ( \6273 , \6270 , \361 );
nand \U$5931 ( \6274 , \6272 , \6273 );
nand \U$5932 ( \6275 , \6266 , \6274 );
nand \U$5933 ( \6276 , \6263 , \6275 );
or \U$5934 ( \6277 , \5938 , \5931 );
nand \U$5935 ( \6278 , \6277 , \5939 );
xor \U$5936 ( \6279 , \6276 , \6278 );
xor \U$5937 ( \6280 , \5951 , \5959 );
xor \U$5938 ( \6281 , \6280 , \5968 );
and \U$5939 ( \6282 , \6279 , \6281 );
and \U$5940 ( \6283 , \6276 , \6278 );
or \U$5941 ( \6284 , \6282 , \6283 );
and \U$5942 ( \6285 , \6254 , \6284 );
and \U$5943 ( \6286 , \6170 , \6253 );
or \U$5944 ( \6287 , \6285 , \6286 );
xor \U$5945 ( \6288 , \6082 , \6287 );
xor \U$5946 ( \6289 , \5978 , \5985 );
xor \U$5947 ( \6290 , \6289 , \5994 );
xor \U$5948 ( \6291 , \6005 , \6012 );
xor \U$5949 ( \6292 , \6291 , \6021 );
xor \U$5950 ( \6293 , \6290 , \6292 );
not \U$5951 ( \6294 , \5841 );
not \U$5952 ( \6295 , \5852 );
or \U$5953 ( \6296 , \6294 , \6295 );
or \U$5954 ( \6297 , \5841 , \5852 );
nand \U$5955 ( \6298 , \6296 , \6297 );
not \U$5956 ( \6299 , \6298 );
not \U$5957 ( \6300 , \5834 );
and \U$5958 ( \6301 , \6299 , \6300 );
and \U$5959 ( \6302 , \6298 , \5834 );
nor \U$5960 ( \6303 , \6301 , \6302 );
and \U$5961 ( \6304 , \6293 , \6303 );
and \U$5962 ( \6305 , \6290 , \6292 );
nor \U$5963 ( \6306 , \6304 , \6305 );
xor \U$5964 ( \6307 , \5898 , \5906 );
xor \U$5965 ( \6308 , \6307 , \5914 );
not \U$5966 ( \6309 , \6308 );
not \U$5967 ( \6310 , \5887 );
not \U$5968 ( \6311 , \5869 );
or \U$5969 ( \6312 , \6310 , \6311 );
or \U$5970 ( \6313 , \5869 , \5887 );
nand \U$5971 ( \6314 , \6312 , \6313 );
not \U$5972 ( \6315 , \6314 );
not \U$5973 ( \6316 , \5862 );
and \U$5974 ( \6317 , \6315 , \6316 );
and \U$5975 ( \6318 , \6314 , \5862 );
nor \U$5976 ( \6319 , \6317 , \6318 );
nor \U$5977 ( \6320 , \6309 , \6319 );
xor \U$5978 ( \6321 , \6306 , \6320 );
xor \U$5979 ( \6322 , \5564 , \5572 );
xor \U$5980 ( \6323 , \6322 , \5580 );
xor \U$5981 ( \6324 , \5813 , \5818 );
xor \U$5982 ( \6325 , \6323 , \6324 );
and \U$5983 ( \6326 , \6321 , \6325 );
and \U$5984 ( \6327 , \6306 , \6320 );
or \U$5985 ( \6328 , \6326 , \6327 );
and \U$5986 ( \6329 , \6288 , \6328 );
and \U$5987 ( \6330 , \6082 , \6287 );
or \U$5988 ( \6331 , \6329 , \6330 );
xor \U$5989 ( \6332 , \5583 , \5606 );
xor \U$5990 ( \6333 , \6332 , \5633 );
xor \U$5991 ( \6334 , \5675 , \5703 );
xor \U$5992 ( \6335 , \6334 , \5730 );
xor \U$5993 ( \6336 , \6333 , \6335 );
xor \U$5994 ( \6337 , \6033 , \6035 );
xor \U$5995 ( \6338 , \6337 , \6040 );
and \U$5996 ( \6339 , \6336 , \6338 );
and \U$5997 ( \6340 , \6333 , \6335 );
or \U$5998 ( \6341 , \6339 , \6340 );
xor \U$5999 ( \6342 , \6331 , \6341 );
xor \U$6000 ( \6343 , \5749 , \5751 );
xor \U$6001 ( \6344 , \6343 , \5756 );
xor \U$6002 ( \6345 , \5784 , \5791 );
xor \U$6003 ( \6346 , \6344 , \6345 );
and \U$6004 ( \6347 , \6342 , \6346 );
and \U$6005 ( \6348 , \6331 , \6341 );
or \U$6006 ( \6349 , \6347 , \6348 );
xor \U$6007 ( \6350 , \5556 , \5736 );
xor \U$6008 ( \6351 , \6350 , \5759 );
xor \U$6009 ( \6352 , \6349 , \6351 );
xor \U$6010 ( \6353 , \5796 , \6046 );
xor \U$6011 ( \6354 , \6353 , \6051 );
and \U$6012 ( \6355 , \6352 , \6354 );
and \U$6013 ( \6356 , \6349 , \6351 );
or \U$6014 ( \6357 , \6355 , \6356 );
xor \U$6015 ( \6358 , \6054 , \6056 );
xor \U$6016 ( \6359 , \6358 , \6059 );
and \U$6017 ( \6360 , \6357 , \6359 );
and \U$6018 ( \6361 , \6068 , \6360 );
xor \U$6019 ( \6362 , \6360 , \6068 );
xor \U$6020 ( \6363 , \6192 , \6221 );
xor \U$6021 ( \6364 , \6363 , \6250 );
xor \U$6022 ( \6365 , \6110 , \6138 );
xor \U$6023 ( \6366 , \6365 , \6167 );
or \U$6024 ( \6367 , \6364 , \6366 );
not \U$6025 ( \6368 , \6366 );
not \U$6026 ( \6369 , \6364 );
or \U$6027 ( \6370 , \6368 , \6369 );
xor \U$6028 ( \6371 , \6276 , \6278 );
xor \U$6029 ( \6372 , \6371 , \6281 );
nand \U$6030 ( \6373 , \6370 , \6372 );
nand \U$6031 ( \6374 , \6367 , \6373 );
xor \U$6032 ( \6375 , \6147 , \6155 );
xor \U$6033 ( \6376 , \6375 , \6164 );
not \U$6034 ( \6377 , \6376 );
and \U$6035 ( \6378 , \416 , RI9871140_113);
and \U$6036 ( \6379 , RI9871320_117, \414 );
nor \U$6037 ( \6380 , \6378 , \6379 );
and \U$6038 ( \6381 , \6380 , \421 );
not \U$6039 ( \6382 , \6380 );
and \U$6040 ( \6383 , \6382 , \422 );
nor \U$6041 ( \6384 , \6381 , \6383 );
nand \U$6042 ( \6385 , RI9871230_115, RI9871fc8_144);
xor \U$6043 ( \6386 , \6384 , \6385 );
and \U$6044 ( \6387 , \354 , RI9871410_119);
and \U$6045 ( \6388 , RI98716e0_125, \352 );
nor \U$6046 ( \6389 , \6387 , \6388 );
not \U$6047 ( \6390 , \6389 );
not \U$6048 ( \6391 , \345 );
and \U$6049 ( \6392 , \6390 , \6391 );
and \U$6050 ( \6393 , \6389 , \361 );
nor \U$6051 ( \6394 , \6392 , \6393 );
and \U$6052 ( \6395 , \6386 , \6394 );
and \U$6053 ( \6396 , \6384 , \6385 );
or \U$6054 ( \6397 , \6395 , \6396 );
not \U$6055 ( \6398 , \6397 );
and \U$6056 ( \6399 , \6377 , \6398 );
and \U$6057 ( \6400 , \6376 , \6397 );
not \U$6058 ( \6401 , \6261 );
not \U$6059 ( \6402 , \6274 );
or \U$6060 ( \6403 , \6401 , \6402 );
or \U$6061 ( \6404 , \6261 , \6274 );
nand \U$6062 ( \6405 , \6403 , \6404 );
not \U$6063 ( \6406 , \6405 );
not \U$6064 ( \6407 , \6262 );
and \U$6065 ( \6408 , \6406 , \6407 );
and \U$6066 ( \6409 , \6405 , \6262 );
nor \U$6067 ( \6410 , \6408 , \6409 );
nor \U$6068 ( \6411 , \6400 , \6410 );
nor \U$6069 ( \6412 , \6399 , \6411 );
not \U$6070 ( \6413 , \4519 );
and \U$6071 ( \6414 , \4710 , RI986dea0_5);
and \U$6072 ( \6415 , RI986ddb0_3, \4708 );
nor \U$6073 ( \6416 , \6414 , \6415 );
not \U$6074 ( \6417 , \6416 );
or \U$6075 ( \6418 , \6413 , \6417 );
or \U$6076 ( \6419 , \6416 , \4519 );
nand \U$6077 ( \6420 , \6418 , \6419 );
not \U$6078 ( \6421 , \3412 );
and \U$6079 ( \6422 , \3683 , RI986f340_49);
and \U$6080 ( \6423 , RI986f520_53, \3681 );
nor \U$6081 ( \6424 , \6422 , \6423 );
not \U$6082 ( \6425 , \6424 );
or \U$6083 ( \6426 , \6421 , \6425 );
or \U$6084 ( \6427 , \6424 , \3918 );
nand \U$6085 ( \6428 , \6426 , \6427 );
xor \U$6086 ( \6429 , \6420 , \6428 );
and \U$6087 ( \6430 , \4203 , RI986f610_55);
and \U$6088 ( \6431 , RI986df90_7, \4201 );
nor \U$6089 ( \6432 , \6430 , \6431 );
and \U$6090 ( \6433 , \6432 , \4207 );
not \U$6091 ( \6434 , \6432 );
and \U$6092 ( \6435 , \6434 , \3923 );
nor \U$6093 ( \6436 , \6433 , \6435 );
and \U$6094 ( \6437 , \6429 , \6436 );
and \U$6095 ( \6438 , \6420 , \6428 );
or \U$6096 ( \6439 , \6437 , \6438 );
and \U$6097 ( \6440 , \5318 , RI986dcc0_1);
and \U$6098 ( \6441 , RI986e170_11, \5316 );
nor \U$6099 ( \6442 , \6440 , \6441 );
and \U$6100 ( \6443 , \6442 , \5052 );
not \U$6101 ( \6444 , \6442 );
and \U$6102 ( \6445 , \6444 , \5322 );
nor \U$6103 ( \6446 , \6443 , \6445 );
and \U$6104 ( \6447 , RI9872a18_166, RI9872b08_168);
not \U$6105 ( \6448 , RI9872b80_169);
and \U$6106 ( \6449 , \6448 , RI9872b08_168);
nor \U$6107 ( \6450 , \6448 , RI9872b08_168);
or \U$6108 ( \6451 , \6449 , \6450 );
nor \U$6109 ( \6452 , RI9872a18_166, RI9872b08_168);
nor \U$6110 ( \6453 , \6447 , \6451 , \6452 );
nand \U$6111 ( \6454 , RI986e350_15, \6453 );
and \U$6112 ( \6455 , \6454 , \6190 );
not \U$6113 ( \6456 , \6454 );
and \U$6114 ( \6457 , \6456 , \6180 );
nor \U$6115 ( \6458 , \6455 , \6457 );
xor \U$6116 ( \6459 , \6446 , \6458 );
and \U$6117 ( \6460 , \5881 , RI986e080_9);
and \U$6118 ( \6461 , RI986e260_13, \5879 );
nor \U$6119 ( \6462 , \6460 , \6461 );
and \U$6120 ( \6463 , \6462 , \5594 );
not \U$6121 ( \6464 , \6462 );
and \U$6122 ( \6465 , \6464 , \5885 );
nor \U$6123 ( \6466 , \6463 , \6465 );
and \U$6124 ( \6467 , \6459 , \6466 );
and \U$6125 ( \6468 , \6446 , \6458 );
or \U$6126 ( \6469 , \6467 , \6468 );
xor \U$6127 ( \6470 , \6439 , \6469 );
and \U$6128 ( \6471 , \2464 , RI986f700_57);
and \U$6129 ( \6472 , RI986f9d0_63, \2462 );
nor \U$6130 ( \6473 , \6471 , \6472 );
and \U$6131 ( \6474 , \6473 , \2468 );
not \U$6132 ( \6475 , \6473 );
and \U$6133 ( \6476 , \6475 , \2263 );
nor \U$6134 ( \6477 , \6474 , \6476 );
and \U$6135 ( \6478 , \2274 , RI986e620_21);
and \U$6136 ( \6479 , RI986f7f0_59, \2272 );
nor \U$6137 ( \6480 , \6478 , \6479 );
and \U$6138 ( \6481 , \6480 , \2030 );
not \U$6139 ( \6482 , \6480 );
and \U$6140 ( \6483 , \6482 , \2031 );
nor \U$6141 ( \6484 , \6481 , \6483 );
xor \U$6142 ( \6485 , \6477 , \6484 );
not \U$6143 ( \6486 , \2935 );
and \U$6144 ( \6487 , \3254 , RI986f8e0_61);
and \U$6145 ( \6488 , RI986f430_51, \3252 );
nor \U$6146 ( \6489 , \6487 , \6488 );
not \U$6147 ( \6490 , \6489 );
or \U$6148 ( \6491 , \6486 , \6490 );
or \U$6149 ( \6492 , \6489 , \2935 );
nand \U$6150 ( \6493 , \6491 , \6492 );
and \U$6151 ( \6494 , \6485 , \6493 );
and \U$6152 ( \6495 , \6477 , \6484 );
or \U$6153 ( \6496 , \6494 , \6495 );
and \U$6154 ( \6497 , \6470 , \6496 );
and \U$6155 ( \6498 , \6439 , \6469 );
nor \U$6156 ( \6499 , \6497 , \6498 );
or \U$6157 ( \6500 , \6412 , \6499 );
not \U$6158 ( \6501 , \6499 );
not \U$6159 ( \6502 , \6412 );
or \U$6160 ( \6503 , \6501 , \6502 );
not \U$6161 ( \6504 , \2034 );
and \U$6162 ( \6505 , \2042 , RI986e440_17);
and \U$6163 ( \6506 , RI986e710_23, \2040 );
nor \U$6164 ( \6507 , \6505 , \6506 );
not \U$6165 ( \6508 , \6507 );
or \U$6166 ( \6509 , \6504 , \6508 );
or \U$6167 ( \6510 , \6507 , \1462 );
nand \U$6168 ( \6511 , \6509 , \6510 );
and \U$6169 ( \6512 , \1329 , RI986ef80_41);
and \U$6170 ( \6513 , RI986f250_47, \1327 );
nor \U$6171 ( \6514 , \6512 , \6513 );
and \U$6172 ( \6515 , \6514 , \1336 );
not \U$6173 ( \6516 , \6514 );
and \U$6174 ( \6517 , \6516 , \1337 );
nor \U$6175 ( \6518 , \6515 , \6517 );
xor \U$6176 ( \6519 , \6511 , \6518 );
and \U$6177 ( \6520 , \1311 , RI986f160_45);
and \U$6178 ( \6521 , RI986e530_19, \1309 );
nor \U$6179 ( \6522 , \6520 , \6521 );
and \U$6180 ( \6523 , \6522 , \1458 );
not \U$6181 ( \6524 , \6522 );
and \U$6182 ( \6525 , \6524 , \1318 );
nor \U$6183 ( \6526 , \6523 , \6525 );
and \U$6184 ( \6527 , \6519 , \6526 );
and \U$6185 ( \6528 , \6511 , \6518 );
or \U$6186 ( \6529 , \6527 , \6528 );
not \U$6187 ( \6530 , \454 );
and \U$6188 ( \6531 , \465 , RI986e9e0_29);
and \U$6189 ( \6532 , RI986e8f0_27, \463 );
nor \U$6190 ( \6533 , \6531 , \6532 );
not \U$6191 ( \6534 , \6533 );
or \U$6192 ( \6535 , \6530 , \6534 );
or \U$6193 ( \6536 , \6533 , \456 );
nand \U$6194 ( \6537 , \6535 , \6536 );
not \U$6195 ( \6538 , \365 );
and \U$6196 ( \6539 , \376 , RI98715f0_123);
and \U$6197 ( \6540 , RI986ead0_31, \374 );
nor \U$6198 ( \6541 , \6539 , \6540 );
not \U$6199 ( \6542 , \6541 );
or \U$6200 ( \6543 , \6538 , \6542 );
or \U$6201 ( \6544 , \6541 , \367 );
nand \U$6202 ( \6545 , \6543 , \6544 );
xor \U$6203 ( \6546 , \6537 , \6545 );
not \U$6204 ( \6547 , \386 );
and \U$6205 ( \6548 , \395 , RI98717d0_127);
and \U$6206 ( \6549 , RI9871500_121, \393 );
nor \U$6207 ( \6550 , \6548 , \6549 );
not \U$6208 ( \6551 , \6550 );
or \U$6209 ( \6552 , \6547 , \6551 );
or \U$6210 ( \6553 , \6550 , \487 );
nand \U$6211 ( \6554 , \6552 , \6553 );
and \U$6212 ( \6555 , \6546 , \6554 );
and \U$6213 ( \6556 , \6537 , \6545 );
or \U$6214 ( \6557 , \6555 , \6556 );
xor \U$6215 ( \6558 , \6529 , \6557 );
not \U$6216 ( \6559 , \1128 );
and \U$6217 ( \6560 , \1293 , RI986ecb0_35);
and \U$6218 ( \6561 , RI986f070_43, \1291 );
nor \U$6219 ( \6562 , \6560 , \6561 );
not \U$6220 ( \6563 , \6562 );
or \U$6221 ( \6564 , \6559 , \6563 );
or \U$6222 ( \6565 , \6562 , \1128 );
nand \U$6223 ( \6566 , \6564 , \6565 );
and \U$6224 ( \6567 , \776 , RI986eda0_37);
and \U$6225 ( \6568 , RI986ebc0_33, \774 );
nor \U$6226 ( \6569 , \6567 , \6568 );
and \U$6227 ( \6570 , \6569 , \474 );
not \U$6228 ( \6571 , \6569 );
and \U$6229 ( \6572 , \6571 , \451 );
nor \U$6230 ( \6573 , \6570 , \6572 );
xor \U$6231 ( \6574 , \6566 , \6573 );
and \U$6232 ( \6575 , \438 , RI986e800_25);
and \U$6233 ( \6576 , RI986ee90_39, \436 );
nor \U$6234 ( \6577 , \6575 , \6576 );
and \U$6235 ( \6578 , \6577 , \444 );
not \U$6236 ( \6579 , \6577 );
and \U$6237 ( \6580 , \6579 , \443 );
nor \U$6238 ( \6581 , \6578 , \6580 );
and \U$6239 ( \6582 , \6574 , \6581 );
and \U$6240 ( \6583 , \6566 , \6573 );
or \U$6241 ( \6584 , \6582 , \6583 );
and \U$6242 ( \6585 , \6558 , \6584 );
and \U$6243 ( \6586 , \6529 , \6557 );
or \U$6244 ( \6587 , \6585 , \6586 );
nand \U$6245 ( \6588 , \6503 , \6587 );
nand \U$6246 ( \6589 , \6500 , \6588 );
xor \U$6247 ( \6590 , \6374 , \6589 );
xor \U$6248 ( \6591 , \6290 , \6292 );
xor \U$6249 ( \6592 , \6591 , \6303 );
not \U$6250 ( \6593 , \6319 );
not \U$6251 ( \6594 , \6308 );
and \U$6252 ( \6595 , \6593 , \6594 );
and \U$6253 ( \6596 , \6319 , \6308 );
nor \U$6254 ( \6597 , \6595 , \6596 );
or \U$6255 ( \6598 , \6592 , \6597 );
not \U$6256 ( \6599 , \6597 );
not \U$6257 ( \6600 , \6592 );
or \U$6258 ( \6601 , \6599 , \6600 );
not \U$6259 ( \6602 , \6097 );
xor \U$6260 ( \6603 , \6089 , \6108 );
not \U$6261 ( \6604 , \6603 );
or \U$6262 ( \6605 , \6602 , \6604 );
or \U$6263 ( \6606 , \6603 , \6097 );
nand \U$6264 ( \6607 , \6605 , \6606 );
not \U$6265 ( \6608 , \6117 );
xor \U$6266 ( \6609 , \6125 , \6136 );
not \U$6267 ( \6610 , \6609 );
or \U$6268 ( \6611 , \6608 , \6610 );
or \U$6269 ( \6612 , \6609 , \6117 );
nand \U$6270 ( \6613 , \6611 , \6612 );
xor \U$6271 ( \6614 , \6607 , \6613 );
not \U$6272 ( \6615 , \6229 );
xor \U$6273 ( \6616 , \6237 , \6248 );
not \U$6274 ( \6617 , \6616 );
or \U$6275 ( \6618 , \6615 , \6617 );
or \U$6276 ( \6619 , \6616 , \6229 );
nand \U$6277 ( \6620 , \6618 , \6619 );
and \U$6278 ( \6621 , \6614 , \6620 );
and \U$6279 ( \6622 , \6607 , \6613 );
or \U$6280 ( \6623 , \6621 , \6622 );
nand \U$6281 ( \6624 , \6601 , \6623 );
nand \U$6282 ( \6625 , \6598 , \6624 );
xor \U$6283 ( \6626 , \6590 , \6625 );
xor \U$6284 ( \6627 , \6306 , \6320 );
xor \U$6285 ( \6628 , \6627 , \6325 );
xor \U$6286 ( \6629 , \5854 , \5889 );
xor \U$6287 ( \6630 , \6629 , \5917 );
xor \U$6288 ( \6631 , \5971 , \5997 );
xor \U$6289 ( \6632 , \6631 , \6024 );
xor \U$6290 ( \6633 , \6070 , \6077 );
xor \U$6291 ( \6634 , \6632 , \6633 );
xor \U$6292 ( \6635 , \6630 , \6634 );
xor \U$6293 ( \6636 , \6628 , \6635 );
xor \U$6294 ( \6637 , \6626 , \6636 );
not \U$6295 ( \6638 , \6637 );
xor \U$6296 ( \6639 , \6446 , \6458 );
xor \U$6297 ( \6640 , \6639 , \6466 );
xor \U$6298 ( \6641 , \6477 , \6484 );
xor \U$6299 ( \6642 , \6641 , \6493 );
and \U$6300 ( \6643 , \6640 , \6642 );
xor \U$6301 ( \6644 , \6420 , \6428 );
xor \U$6302 ( \6645 , \6644 , \6436 );
xor \U$6303 ( \6646 , \6477 , \6484 );
xor \U$6304 ( \6647 , \6646 , \6493 );
and \U$6305 ( \6648 , \6645 , \6647 );
and \U$6306 ( \6649 , \6640 , \6645 );
or \U$6307 ( \6650 , \6643 , \6648 , \6649 );
not \U$6308 ( \6651 , \6200 );
xor \U$6309 ( \6652 , \6208 , \6219 );
not \U$6310 ( \6653 , \6652 );
or \U$6311 ( \6654 , \6651 , \6653 );
or \U$6312 ( \6655 , \6652 , \6200 );
nand \U$6313 ( \6656 , \6654 , \6655 );
xor \U$6314 ( \6657 , \6650 , \6656 );
xor \U$6315 ( \6658 , \6566 , \6573 );
xor \U$6316 ( \6659 , \6658 , \6581 );
xor \U$6317 ( \6660 , \6537 , \6545 );
xor \U$6318 ( \6661 , \6660 , \6554 );
and \U$6319 ( \6662 , \6659 , \6661 );
xor \U$6320 ( \6663 , \6511 , \6518 );
xor \U$6321 ( \6664 , \6663 , \6526 );
xor \U$6322 ( \6665 , \6537 , \6545 );
xor \U$6323 ( \6666 , \6665 , \6554 );
and \U$6324 ( \6667 , \6664 , \6666 );
and \U$6325 ( \6668 , \6659 , \6664 );
or \U$6326 ( \6669 , \6662 , \6667 , \6668 );
and \U$6327 ( \6670 , \6657 , \6669 );
and \U$6328 ( \6671 , \6650 , \6656 );
or \U$6329 ( \6672 , \6670 , \6671 );
not \U$6330 ( \6673 , \3412 );
and \U$6331 ( \6674 , \3683 , RI986f430_51);
and \U$6332 ( \6675 , RI986f340_49, \3681 );
nor \U$6333 ( \6676 , \6674 , \6675 );
not \U$6334 ( \6677 , \6676 );
or \U$6335 ( \6678 , \6673 , \6677 );
or \U$6336 ( \6679 , \6676 , \3918 );
nand \U$6337 ( \6680 , \6678 , \6679 );
and \U$6338 ( \6681 , \2464 , RI986f7f0_59);
and \U$6339 ( \6682 , RI986f700_57, \2462 );
nor \U$6340 ( \6683 , \6681 , \6682 );
and \U$6341 ( \6684 , \6683 , \2468 );
not \U$6342 ( \6685 , \6683 );
and \U$6343 ( \6686 , \6685 , \2263 );
nor \U$6344 ( \6687 , \6684 , \6686 );
xor \U$6345 ( \6688 , \6680 , \6687 );
not \U$6346 ( \6689 , \3406 );
and \U$6347 ( \6690 , \3254 , RI986f9d0_63);
and \U$6348 ( \6691 , RI986f8e0_61, \3252 );
nor \U$6349 ( \6692 , \6690 , \6691 );
not \U$6350 ( \6693 , \6692 );
or \U$6351 ( \6694 , \6689 , \6693 );
or \U$6352 ( \6695 , \6692 , \3406 );
nand \U$6353 ( \6696 , \6694 , \6695 );
and \U$6354 ( \6697 , \6688 , \6696 );
and \U$6355 ( \6698 , \6680 , \6687 );
or \U$6356 ( \6699 , \6697 , \6698 );
and \U$6357 ( \6700 , \6453 , RI986e260_13);
and \U$6358 ( \6701 , RI986e350_15, \6451 );
nor \U$6359 ( \6702 , \6700 , \6701 );
and \U$6360 ( \6703 , \6702 , \6190 );
not \U$6361 ( \6704 , \6702 );
buf \U$6362 ( \6705 , \6180 );
and \U$6363 ( \6706 , \6704 , \6705 );
nor \U$6364 ( \6707 , \6703 , \6706 );
nand \U$6365 ( \6708 , RI9872bf8_170, RI9872c70_171);
and \U$6366 ( \6709 , \6708 , RI9872b80_169);
not \U$6367 ( \6710 , \6709 );
xor \U$6368 ( \6711 , \6707 , \6710 );
and \U$6369 ( \6712 , \5881 , RI986e170_11);
and \U$6370 ( \6713 , RI986e080_9, \5879 );
nor \U$6371 ( \6714 , \6712 , \6713 );
and \U$6372 ( \6715 , \6714 , \5594 );
not \U$6373 ( \6716 , \6714 );
and \U$6374 ( \6717 , \6716 , \5885 );
nor \U$6375 ( \6718 , \6715 , \6717 );
and \U$6376 ( \6719 , \6711 , \6718 );
and \U$6377 ( \6720 , \6707 , \6710 );
or \U$6378 ( \6721 , \6719 , \6720 );
xor \U$6379 ( \6722 , \6699 , \6721 );
and \U$6380 ( \6723 , \4203 , RI986f520_53);
and \U$6381 ( \6724 , RI986f610_55, \4201 );
nor \U$6382 ( \6725 , \6723 , \6724 );
and \U$6383 ( \6726 , \6725 , \3922 );
not \U$6384 ( \6727 , \6725 );
and \U$6385 ( \6728 , \6727 , \4207 );
nor \U$6386 ( \6729 , \6726 , \6728 );
and \U$6387 ( \6730 , \4710 , RI986df90_7);
and \U$6388 ( \6731 , RI986dea0_5, \4708 );
nor \U$6389 ( \6732 , \6730 , \6731 );
not \U$6390 ( \6733 , \6732 );
not \U$6391 ( \6734 , \4519 );
and \U$6392 ( \6735 , \6733 , \6734 );
and \U$6393 ( \6736 , \6732 , \4521 );
nor \U$6394 ( \6737 , \6735 , \6736 );
or \U$6395 ( \6738 , \6729 , \6737 );
not \U$6396 ( \6739 , \6737 );
not \U$6397 ( \6740 , \6729 );
or \U$6398 ( \6741 , \6739 , \6740 );
and \U$6399 ( \6742 , \5318 , RI986ddb0_3);
and \U$6400 ( \6743 , RI986dcc0_1, \5316 );
nor \U$6401 ( \6744 , \6742 , \6743 );
and \U$6402 ( \6745 , \6744 , \5052 );
not \U$6403 ( \6746 , \6744 );
and \U$6404 ( \6747 , \6746 , \5322 );
nor \U$6405 ( \6748 , \6745 , \6747 );
nand \U$6406 ( \6749 , \6741 , \6748 );
nand \U$6407 ( \6750 , \6738 , \6749 );
and \U$6408 ( \6751 , \6722 , \6750 );
and \U$6409 ( \6752 , \6699 , \6721 );
or \U$6410 ( \6753 , \6751 , \6752 );
and \U$6411 ( \6754 , \416 , RI9871230_115);
and \U$6412 ( \6755 , RI9871140_113, \414 );
nor \U$6413 ( \6756 , \6754 , \6755 );
and \U$6414 ( \6757 , \6756 , \421 );
not \U$6415 ( \6758 , \6756 );
and \U$6416 ( \6759 , \6758 , \422 );
nor \U$6417 ( \6760 , \6757 , \6759 );
and \U$6418 ( \6761 , \395 , RI98716e0_125);
and \U$6419 ( \6762 , RI98717d0_127, \393 );
nor \U$6420 ( \6763 , \6761 , \6762 );
not \U$6421 ( \6764 , \6763 );
not \U$6422 ( \6765 , \487 );
and \U$6423 ( \6766 , \6764 , \6765 );
and \U$6424 ( \6767 , \6763 , \386 );
nor \U$6425 ( \6768 , \6766 , \6767 );
xor \U$6426 ( \6769 , \6760 , \6768 );
and \U$6427 ( \6770 , \354 , RI9871320_117);
and \U$6428 ( \6771 , RI9871410_119, \352 );
nor \U$6429 ( \6772 , \6770 , \6771 );
not \U$6430 ( \6773 , \6772 );
not \U$6431 ( \6774 , \345 );
and \U$6432 ( \6775 , \6773 , \6774 );
and \U$6433 ( \6776 , \6772 , \345 );
nor \U$6434 ( \6777 , \6775 , \6776 );
and \U$6435 ( \6778 , \6769 , \6777 );
and \U$6436 ( \6779 , \6760 , \6768 );
or \U$6437 ( \6780 , \6778 , \6779 );
xor \U$6438 ( \6781 , \6384 , \6385 );
xor \U$6439 ( \6782 , \6781 , \6394 );
nand \U$6440 ( \6783 , \6780 , \6782 );
xor \U$6441 ( \6784 , \6753 , \6783 );
and \U$6442 ( \6785 , \1311 , RI986f250_47);
and \U$6443 ( \6786 , RI986f160_45, \1309 );
nor \U$6444 ( \6787 , \6785 , \6786 );
and \U$6445 ( \6788 , \6787 , \1315 );
not \U$6446 ( \6789 , \6787 );
and \U$6447 ( \6790 , \6789 , \1458 );
nor \U$6448 ( \6791 , \6788 , \6790 );
and \U$6449 ( \6792 , \2042 , RI986e530_19);
and \U$6450 ( \6793 , RI986e440_17, \2040 );
nor \U$6451 ( \6794 , \6792 , \6793 );
not \U$6452 ( \6795 , \6794 );
not \U$6453 ( \6796 , \2034 );
and \U$6454 ( \6797 , \6795 , \6796 );
and \U$6455 ( \6798 , \6794 , \1462 );
nor \U$6456 ( \6799 , \6797 , \6798 );
or \U$6457 ( \6800 , \6791 , \6799 );
not \U$6458 ( \6801 , \6799 );
not \U$6459 ( \6802 , \6791 );
or \U$6460 ( \6803 , \6801 , \6802 );
and \U$6461 ( \6804 , \2274 , RI986e710_23);
and \U$6462 ( \6805 , RI986e620_21, \2272 );
nor \U$6463 ( \6806 , \6804 , \6805 );
and \U$6464 ( \6807 , \6806 , \2030 );
not \U$6465 ( \6808 , \6806 );
and \U$6466 ( \6809 , \6808 , \2031 );
nor \U$6467 ( \6810 , \6807 , \6809 );
nand \U$6468 ( \6811 , \6803 , \6810 );
nand \U$6469 ( \6812 , \6800 , \6811 );
and \U$6470 ( \6813 , \465 , RI986ead0_31);
and \U$6471 ( \6814 , RI986e9e0_29, \463 );
nor \U$6472 ( \6815 , \6813 , \6814 );
not \U$6473 ( \6816 , \6815 );
not \U$6474 ( \6817 , \454 );
and \U$6475 ( \6818 , \6816 , \6817 );
and \U$6476 ( \6819 , \6815 , \456 );
nor \U$6477 ( \6820 , \6818 , \6819 );
and \U$6478 ( \6821 , \376 , RI9871500_121);
and \U$6479 ( \6822 , RI98715f0_123, \374 );
nor \U$6480 ( \6823 , \6821 , \6822 );
not \U$6481 ( \6824 , \6823 );
not \U$6482 ( \6825 , \365 );
and \U$6483 ( \6826 , \6824 , \6825 );
and \U$6484 ( \6827 , \6823 , \365 );
nor \U$6485 ( \6828 , \6826 , \6827 );
or \U$6486 ( \6829 , \6820 , \6828 );
not \U$6487 ( \6830 , \6828 );
not \U$6488 ( \6831 , \6820 );
or \U$6489 ( \6832 , \6830 , \6831 );
and \U$6490 ( \6833 , \438 , RI986e8f0_27);
and \U$6491 ( \6834 , RI986e800_25, \436 );
nor \U$6492 ( \6835 , \6833 , \6834 );
and \U$6493 ( \6836 , \6835 , \444 );
not \U$6494 ( \6837 , \6835 );
and \U$6495 ( \6838 , \6837 , \443 );
nor \U$6496 ( \6839 , \6836 , \6838 );
nand \U$6497 ( \6840 , \6832 , \6839 );
nand \U$6498 ( \6841 , \6829 , \6840 );
xor \U$6499 ( \6842 , \6812 , \6841 );
and \U$6500 ( \6843 , \776 , RI986ee90_39);
and \U$6501 ( \6844 , RI986eda0_37, \774 );
nor \U$6502 ( \6845 , \6843 , \6844 );
and \U$6503 ( \6846 , \6845 , \451 );
not \U$6504 ( \6847 , \6845 );
and \U$6505 ( \6848 , \6847 , \474 );
nor \U$6506 ( \6849 , \6846 , \6848 );
and \U$6507 ( \6850 , \1293 , RI986ebc0_33);
and \U$6508 ( \6851 , RI986ecb0_35, \1291 );
nor \U$6509 ( \6852 , \6850 , \6851 );
not \U$6510 ( \6853 , \6852 );
not \U$6511 ( \6854 , \1128 );
and \U$6512 ( \6855 , \6853 , \6854 );
and \U$6513 ( \6856 , \6852 , \1128 );
nor \U$6514 ( \6857 , \6855 , \6856 );
or \U$6515 ( \6858 , \6849 , \6857 );
not \U$6516 ( \6859 , \6857 );
not \U$6517 ( \6860 , \6849 );
or \U$6518 ( \6861 , \6859 , \6860 );
and \U$6519 ( \6862 , \1329 , RI986f070_43);
and \U$6520 ( \6863 , RI986ef80_41, \1327 );
nor \U$6521 ( \6864 , \6862 , \6863 );
and \U$6522 ( \6865 , \6864 , \1336 );
not \U$6523 ( \6866 , \6864 );
and \U$6524 ( \6867 , \6866 , \1337 );
nor \U$6525 ( \6868 , \6865 , \6867 );
nand \U$6526 ( \6869 , \6861 , \6868 );
nand \U$6527 ( \6870 , \6858 , \6869 );
and \U$6528 ( \6871 , \6842 , \6870 );
and \U$6529 ( \6872 , \6812 , \6841 );
or \U$6530 ( \6873 , \6871 , \6872 );
and \U$6531 ( \6874 , \6784 , \6873 );
and \U$6532 ( \6875 , \6753 , \6783 );
or \U$6533 ( \6876 , \6874 , \6875 );
xor \U$6534 ( \6877 , \6672 , \6876 );
not \U$6535 ( \6878 , \6376 );
xor \U$6536 ( \6879 , \6397 , \6410 );
not \U$6537 ( \6880 , \6879 );
or \U$6538 ( \6881 , \6878 , \6880 );
or \U$6539 ( \6882 , \6879 , \6376 );
nand \U$6540 ( \6883 , \6881 , \6882 );
not \U$6541 ( \6884 , \6188 );
and \U$6542 ( \6885 , \6177 , \6180 );
not \U$6543 ( \6886 , \6177 );
and \U$6544 ( \6887 , \6886 , \6190 );
nor \U$6545 ( \6888 , \6885 , \6887 );
not \U$6546 ( \6889 , \6888 );
or \U$6547 ( \6890 , \6884 , \6889 );
or \U$6548 ( \6891 , \6888 , \6188 );
nand \U$6549 ( \6892 , \6890 , \6891 );
xor \U$6550 ( \6893 , \6883 , \6892 );
xor \U$6551 ( \6894 , \6607 , \6613 );
xor \U$6552 ( \6895 , \6894 , \6620 );
and \U$6553 ( \6896 , \6893 , \6895 );
and \U$6554 ( \6897 , \6883 , \6892 );
or \U$6555 ( \6898 , \6896 , \6897 );
and \U$6556 ( \6899 , \6877 , \6898 );
and \U$6557 ( \6900 , \6672 , \6876 );
or \U$6558 ( \6901 , \6899 , \6900 );
xor \U$6559 ( \6902 , \6170 , \6253 );
xor \U$6560 ( \6903 , \6902 , \6284 );
xor \U$6561 ( \6904 , \6901 , \6903 );
not \U$6562 ( \6905 , \6499 );
not \U$6563 ( \6906 , \6587 );
or \U$6564 ( \6907 , \6905 , \6906 );
or \U$6565 ( \6908 , \6587 , \6499 );
nand \U$6566 ( \6909 , \6907 , \6908 );
not \U$6567 ( \6910 , \6909 );
not \U$6568 ( \6911 , \6412 );
and \U$6569 ( \6912 , \6910 , \6911 );
and \U$6570 ( \6913 , \6909 , \6412 );
nor \U$6571 ( \6914 , \6912 , \6913 );
xnor \U$6572 ( \6915 , \6364 , \6366 );
not \U$6573 ( \6916 , \6915 );
not \U$6574 ( \6917 , \6372 );
and \U$6575 ( \6918 , \6916 , \6917 );
and \U$6576 ( \6919 , \6915 , \6372 );
nor \U$6577 ( \6920 , \6918 , \6919 );
xor \U$6578 ( \6921 , \6914 , \6920 );
not \U$6579 ( \6922 , \6623 );
not \U$6580 ( \6923 , \6592 );
or \U$6581 ( \6924 , \6922 , \6923 );
or \U$6582 ( \6925 , \6592 , \6623 );
nand \U$6583 ( \6926 , \6924 , \6925 );
not \U$6584 ( \6927 , \6926 );
not \U$6585 ( \6928 , \6597 );
and \U$6586 ( \6929 , \6927 , \6928 );
and \U$6587 ( \6930 , \6926 , \6597 );
nor \U$6588 ( \6931 , \6929 , \6930 );
and \U$6589 ( \6932 , \6921 , \6931 );
and \U$6590 ( \6933 , \6914 , \6920 );
nor \U$6591 ( \6934 , \6932 , \6933 );
xor \U$6592 ( \6935 , \6904 , \6934 );
not \U$6593 ( \6936 , \6935 );
or \U$6594 ( \6937 , \6638 , \6936 );
or \U$6595 ( \6938 , \6935 , \6637 );
xor \U$6596 ( \6939 , \6914 , \6920 );
xor \U$6597 ( \6940 , \6939 , \6931 );
not \U$6598 ( \6941 , \6799 );
not \U$6599 ( \6942 , \6810 );
or \U$6600 ( \6943 , \6941 , \6942 );
or \U$6601 ( \6944 , \6799 , \6810 );
nand \U$6602 ( \6945 , \6943 , \6944 );
not \U$6603 ( \6946 , \6945 );
not \U$6604 ( \6947 , \6791 );
and \U$6605 ( \6948 , \6946 , \6947 );
and \U$6606 ( \6949 , \6945 , \6791 );
nor \U$6607 ( \6950 , \6948 , \6949 );
not \U$6608 ( \6951 , \6737 );
not \U$6609 ( \6952 , \6748 );
or \U$6610 ( \6953 , \6951 , \6952 );
or \U$6611 ( \6954 , \6737 , \6748 );
nand \U$6612 ( \6955 , \6953 , \6954 );
not \U$6613 ( \6956 , \6955 );
not \U$6614 ( \6957 , \6729 );
and \U$6615 ( \6958 , \6956 , \6957 );
and \U$6616 ( \6959 , \6955 , \6729 );
nor \U$6617 ( \6960 , \6958 , \6959 );
or \U$6618 ( \6961 , \6950 , \6960 );
not \U$6619 ( \6962 , \6960 );
not \U$6620 ( \6963 , \6950 );
or \U$6621 ( \6964 , \6962 , \6963 );
xor \U$6622 ( \6965 , \6680 , \6687 );
xor \U$6623 ( \6966 , \6965 , \6696 );
nand \U$6624 ( \6967 , \6964 , \6966 );
nand \U$6625 ( \6968 , \6961 , \6967 );
not \U$6626 ( \6969 , \6820 );
not \U$6627 ( \6970 , \6839 );
or \U$6628 ( \6971 , \6969 , \6970 );
or \U$6629 ( \6972 , \6820 , \6839 );
nand \U$6630 ( \6973 , \6971 , \6972 );
not \U$6631 ( \6974 , \6973 );
not \U$6632 ( \6975 , \6828 );
and \U$6633 ( \6976 , \6974 , \6975 );
and \U$6634 ( \6977 , \6973 , \6828 );
nor \U$6635 ( \6978 , \6976 , \6977 );
not \U$6636 ( \6979 , \6857 );
not \U$6637 ( \6980 , \6868 );
or \U$6638 ( \6981 , \6979 , \6980 );
or \U$6639 ( \6982 , \6857 , \6868 );
nand \U$6640 ( \6983 , \6981 , \6982 );
not \U$6641 ( \6984 , \6983 );
not \U$6642 ( \6985 , \6849 );
and \U$6643 ( \6986 , \6984 , \6985 );
and \U$6644 ( \6987 , \6983 , \6849 );
nor \U$6645 ( \6988 , \6986 , \6987 );
xor \U$6646 ( \6989 , \6978 , \6988 );
xor \U$6647 ( \6990 , \6760 , \6768 );
xor \U$6648 ( \6991 , \6990 , \6777 );
and \U$6649 ( \6992 , \6989 , \6991 );
and \U$6650 ( \6993 , \6978 , \6988 );
nor \U$6651 ( \6994 , \6992 , \6993 );
xor \U$6652 ( \6995 , \6968 , \6994 );
xor \U$6653 ( \6996 , \6477 , \6484 );
xor \U$6654 ( \6997 , \6996 , \6493 );
xor \U$6655 ( \6998 , \6640 , \6645 );
xor \U$6656 ( \6999 , \6997 , \6998 );
and \U$6657 ( \7000 , \6995 , \6999 );
and \U$6658 ( \7001 , \6968 , \6994 );
or \U$6659 ( \7002 , \7000 , \7001 );
nand \U$6660 ( \7003 , RI9871050_111, RI9871fc8_144);
nand \U$6661 ( \7004 , RI9870c90_103, RI9871fc8_144);
xor \U$6662 ( \7005 , \7003 , \7004 );
and \U$6663 ( \7006 , \395 , RI9871410_119);
and \U$6664 ( \7007 , RI98716e0_125, \393 );
nor \U$6665 ( \7008 , \7006 , \7007 );
not \U$6666 ( \7009 , \7008 );
not \U$6667 ( \7010 , \487 );
and \U$6668 ( \7011 , \7009 , \7010 );
and \U$6669 ( \7012 , \7008 , \487 );
nor \U$6670 ( \7013 , \7011 , \7012 );
not \U$6671 ( \7014 , \7013 );
and \U$6672 ( \7015 , \416 , RI9870c90_103);
and \U$6673 ( \7016 , RI9871230_115, \414 );
nor \U$6674 ( \7017 , \7015 , \7016 );
and \U$6675 ( \7018 , \7017 , \421 );
not \U$6676 ( \7019 , \7017 );
and \U$6677 ( \7020 , \7019 , \422 );
nor \U$6678 ( \7021 , \7018 , \7020 );
not \U$6679 ( \7022 , \7021 );
and \U$6680 ( \7023 , \7014 , \7022 );
and \U$6681 ( \7024 , \7013 , \7021 );
and \U$6682 ( \7025 , \354 , RI9871140_113);
and \U$6683 ( \7026 , RI9871320_117, \352 );
nor \U$6684 ( \7027 , \7025 , \7026 );
not \U$6685 ( \7028 , \7027 );
not \U$6686 ( \7029 , \345 );
and \U$6687 ( \7030 , \7028 , \7029 );
and \U$6688 ( \7031 , \7027 , \361 );
nor \U$6689 ( \7032 , \7030 , \7031 );
nor \U$6690 ( \7033 , \7024 , \7032 );
nor \U$6691 ( \7034 , \7023 , \7033 );
and \U$6692 ( \7035 , \7005 , \7034 );
and \U$6693 ( \7036 , \7003 , \7004 );
or \U$6694 ( \7037 , \7035 , \7036 );
and \U$6695 ( \7038 , \2464 , RI986e620_21);
and \U$6696 ( \7039 , RI986f7f0_59, \2462 );
nor \U$6697 ( \7040 , \7038 , \7039 );
and \U$6698 ( \7041 , \7040 , \2468 );
not \U$6699 ( \7042 , \7040 );
and \U$6700 ( \7043 , \7042 , \2263 );
nor \U$6701 ( \7044 , \7041 , \7043 );
not \U$6702 ( \7045 , \3406 );
and \U$6703 ( \7046 , \3254 , RI986f700_57);
and \U$6704 ( \7047 , RI986f9d0_63, \3252 );
nor \U$6705 ( \7048 , \7046 , \7047 );
not \U$6706 ( \7049 , \7048 );
or \U$6707 ( \7050 , \7045 , \7049 );
or \U$6708 ( \7051 , \7048 , \2935 );
nand \U$6709 ( \7052 , \7050 , \7051 );
xor \U$6710 ( \7053 , \7044 , \7052 );
not \U$6711 ( \7054 , \3412 );
and \U$6712 ( \7055 , \3683 , RI986f8e0_61);
and \U$6713 ( \7056 , RI986f430_51, \3681 );
nor \U$6714 ( \7057 , \7055 , \7056 );
not \U$6715 ( \7058 , \7057 );
or \U$6716 ( \7059 , \7054 , \7058 );
or \U$6717 ( \7060 , \7057 , \3412 );
nand \U$6718 ( \7061 , \7059 , \7060 );
and \U$6719 ( \7062 , \7053 , \7061 );
and \U$6720 ( \7063 , \7044 , \7052 );
or \U$6721 ( \7064 , \7062 , \7063 );
and \U$6722 ( \7065 , \5881 , RI986dcc0_1);
and \U$6723 ( \7066 , RI986e170_11, \5879 );
nor \U$6724 ( \7067 , \7065 , \7066 );
and \U$6725 ( \7068 , \7067 , \5594 );
not \U$6726 ( \7069 , \7067 );
and \U$6727 ( \7070 , \7069 , \5885 );
nor \U$6728 ( \7071 , \7068 , \7070 );
and \U$6729 ( \7072 , RI9872b80_169, RI9872c70_171);
not \U$6730 ( \7073 , RI9872c70_171);
nor \U$6731 ( \7074 , \7073 , RI9872bf8_170);
not \U$6732 ( \7075 , RI9872bf8_170);
nor \U$6733 ( \7076 , \7075 , RI9872c70_171);
or \U$6734 ( \7077 , \7074 , \7076 );
nor \U$6735 ( \7078 , RI9872b80_169, RI9872c70_171);
nor \U$6736 ( \7079 , \7072 , \7077 , \7078 );
nand \U$6737 ( \7080 , RI986e350_15, \7079 );
and \U$6738 ( \7081 , \7080 , \6710 );
not \U$6739 ( \7082 , \7080 );
and \U$6740 ( \7083 , \7082 , \6709 );
nor \U$6741 ( \7084 , \7081 , \7083 );
xor \U$6742 ( \7085 , \7071 , \7084 );
and \U$6743 ( \7086 , \6453 , RI986e080_9);
and \U$6744 ( \7087 , RI986e260_13, \6451 );
nor \U$6745 ( \7088 , \7086 , \7087 );
and \U$6746 ( \7089 , \7088 , \6190 );
not \U$6747 ( \7090 , \7088 );
and \U$6748 ( \7091 , \7090 , \6705 );
nor \U$6749 ( \7092 , \7089 , \7091 );
and \U$6750 ( \7093 , \7085 , \7092 );
and \U$6751 ( \7094 , \7071 , \7084 );
or \U$6752 ( \7095 , \7093 , \7094 );
xor \U$6753 ( \7096 , \7064 , \7095 );
and \U$6754 ( \7097 , \4203 , RI986f340_49);
and \U$6755 ( \7098 , RI986f520_53, \4201 );
nor \U$6756 ( \7099 , \7097 , \7098 );
and \U$6757 ( \7100 , \7099 , \4207 );
not \U$6758 ( \7101 , \7099 );
and \U$6759 ( \7102 , \7101 , \3922 );
nor \U$6760 ( \7103 , \7100 , \7102 );
not \U$6761 ( \7104 , \4521 );
and \U$6762 ( \7105 , \4710 , RI986f610_55);
and \U$6763 ( \7106 , RI986df90_7, \4708 );
nor \U$6764 ( \7107 , \7105 , \7106 );
not \U$6765 ( \7108 , \7107 );
or \U$6766 ( \7109 , \7104 , \7108 );
or \U$6767 ( \7110 , \7107 , \4519 );
nand \U$6768 ( \7111 , \7109 , \7110 );
xor \U$6769 ( \7112 , \7103 , \7111 );
and \U$6770 ( \7113 , \5318 , RI986dea0_5);
and \U$6771 ( \7114 , RI986ddb0_3, \5316 );
nor \U$6772 ( \7115 , \7113 , \7114 );
and \U$6773 ( \7116 , \7115 , \5052 );
not \U$6774 ( \7117 , \7115 );
and \U$6775 ( \7118 , \7117 , \5322 );
nor \U$6776 ( \7119 , \7116 , \7118 );
and \U$6777 ( \7120 , \7112 , \7119 );
and \U$6778 ( \7121 , \7103 , \7111 );
or \U$6779 ( \7122 , \7120 , \7121 );
and \U$6780 ( \7123 , \7096 , \7122 );
and \U$6781 ( \7124 , \7064 , \7095 );
nor \U$6782 ( \7125 , \7123 , \7124 );
xor \U$6783 ( \7126 , \7037 , \7125 );
and \U$6784 ( \7127 , \776 , RI986e800_25);
and \U$6785 ( \7128 , RI986ee90_39, \774 );
nor \U$6786 ( \7129 , \7127 , \7128 );
and \U$6787 ( \7130 , \7129 , \474 );
not \U$6788 ( \7131 , \7129 );
and \U$6789 ( \7132 , \7131 , \451 );
nor \U$6790 ( \7133 , \7130 , \7132 );
not \U$6791 ( \7134 , \1128 );
and \U$6792 ( \7135 , \1293 , RI986eda0_37);
and \U$6793 ( \7136 , RI986ebc0_33, \1291 );
nor \U$6794 ( \7137 , \7135 , \7136 );
not \U$6795 ( \7138 , \7137 );
or \U$6796 ( \7139 , \7134 , \7138 );
or \U$6797 ( \7140 , \7137 , \1301 );
nand \U$6798 ( \7141 , \7139 , \7140 );
xor \U$6799 ( \7142 , \7133 , \7141 );
and \U$6800 ( \7143 , \1329 , RI986ecb0_35);
and \U$6801 ( \7144 , RI986f070_43, \1327 );
nor \U$6802 ( \7145 , \7143 , \7144 );
and \U$6803 ( \7146 , \7145 , \1336 );
not \U$6804 ( \7147 , \7145 );
and \U$6805 ( \7148 , \7147 , \1337 );
nor \U$6806 ( \7149 , \7146 , \7148 );
and \U$6807 ( \7150 , \7142 , \7149 );
and \U$6808 ( \7151 , \7133 , \7141 );
or \U$6809 ( \7152 , \7150 , \7151 );
not \U$6810 ( \7153 , \367 );
and \U$6811 ( \7154 , \376 , RI98717d0_127);
and \U$6812 ( \7155 , RI9871500_121, \374 );
nor \U$6813 ( \7156 , \7154 , \7155 );
not \U$6814 ( \7157 , \7156 );
or \U$6815 ( \7158 , \7153 , \7157 );
or \U$6816 ( \7159 , \7156 , \365 );
nand \U$6817 ( \7160 , \7158 , \7159 );
and \U$6818 ( \7161 , \438 , RI986e9e0_29);
and \U$6819 ( \7162 , RI986e8f0_27, \436 );
nor \U$6820 ( \7163 , \7161 , \7162 );
and \U$6821 ( \7164 , \7163 , \444 );
not \U$6822 ( \7165 , \7163 );
and \U$6823 ( \7166 , \7165 , \443 );
nor \U$6824 ( \7167 , \7164 , \7166 );
xor \U$6825 ( \7168 , \7160 , \7167 );
not \U$6826 ( \7169 , \454 );
and \U$6827 ( \7170 , \465 , RI98715f0_123);
and \U$6828 ( \7171 , RI986ead0_31, \463 );
nor \U$6829 ( \7172 , \7170 , \7171 );
not \U$6830 ( \7173 , \7172 );
or \U$6831 ( \7174 , \7169 , \7173 );
or \U$6832 ( \7175 , \7172 , \456 );
nand \U$6833 ( \7176 , \7174 , \7175 );
and \U$6834 ( \7177 , \7168 , \7176 );
and \U$6835 ( \7178 , \7160 , \7167 );
or \U$6836 ( \7179 , \7177 , \7178 );
xor \U$6837 ( \7180 , \7152 , \7179 );
and \U$6838 ( \7181 , \1311 , RI986ef80_41);
and \U$6839 ( \7182 , RI986f250_47, \1309 );
nor \U$6840 ( \7183 , \7181 , \7182 );
and \U$6841 ( \7184 , \7183 , \1458 );
not \U$6842 ( \7185 , \7183 );
and \U$6843 ( \7186 , \7185 , \1318 );
nor \U$6844 ( \7187 , \7184 , \7186 );
not \U$6845 ( \7188 , \2034 );
and \U$6846 ( \7189 , \2042 , RI986f160_45);
and \U$6847 ( \7190 , RI986e530_19, \2040 );
nor \U$6848 ( \7191 , \7189 , \7190 );
not \U$6849 ( \7192 , \7191 );
or \U$6850 ( \7193 , \7188 , \7192 );
or \U$6851 ( \7194 , \7191 , \1462 );
nand \U$6852 ( \7195 , \7193 , \7194 );
xor \U$6853 ( \7196 , \7187 , \7195 );
and \U$6854 ( \7197 , \2274 , RI986e440_17);
and \U$6855 ( \7198 , RI986e710_23, \2272 );
nor \U$6856 ( \7199 , \7197 , \7198 );
and \U$6857 ( \7200 , \7199 , \2030 );
not \U$6858 ( \7201 , \7199 );
and \U$6859 ( \7202 , \7201 , \2031 );
nor \U$6860 ( \7203 , \7200 , \7202 );
and \U$6861 ( \7204 , \7196 , \7203 );
and \U$6862 ( \7205 , \7187 , \7195 );
or \U$6863 ( \7206 , \7204 , \7205 );
and \U$6864 ( \7207 , \7180 , \7206 );
and \U$6865 ( \7208 , \7152 , \7179 );
nor \U$6866 ( \7209 , \7207 , \7208 );
and \U$6867 ( \7210 , \7126 , \7209 );
and \U$6868 ( \7211 , \7037 , \7125 );
nor \U$6869 ( \7212 , \7210 , \7211 );
xor \U$6870 ( \7213 , \7002 , \7212 );
or \U$6871 ( \7214 , \6782 , \6780 );
nand \U$6872 ( \7215 , \7214 , \6783 );
xor \U$6873 ( \7216 , \6812 , \6841 );
xor \U$6874 ( \7217 , \7216 , \6870 );
and \U$6875 ( \7218 , \7215 , \7217 );
xor \U$6876 ( \7219 , \6537 , \6545 );
xor \U$6877 ( \7220 , \7219 , \6554 );
xor \U$6878 ( \7221 , \6659 , \6664 );
xor \U$6879 ( \7222 , \7220 , \7221 );
xor \U$6880 ( \7223 , \6812 , \6841 );
xor \U$6881 ( \7224 , \7223 , \6870 );
and \U$6882 ( \7225 , \7222 , \7224 );
and \U$6883 ( \7226 , \7215 , \7222 );
or \U$6884 ( \7227 , \7218 , \7225 , \7226 );
and \U$6885 ( \7228 , \7213 , \7227 );
and \U$6886 ( \7229 , \7002 , \7212 );
nor \U$6887 ( \7230 , \7228 , \7229 );
or \U$6888 ( \7231 , \6940 , \7230 );
not \U$6889 ( \7232 , \7230 );
not \U$6890 ( \7233 , \6940 );
or \U$6891 ( \7234 , \7232 , \7233 );
xor \U$6892 ( \7235 , \6529 , \6557 );
xor \U$6893 ( \7236 , \7235 , \6584 );
xor \U$6894 ( \7237 , \6439 , \6469 );
xor \U$6895 ( \7238 , \7237 , \6496 );
xor \U$6896 ( \7239 , \7236 , \7238 );
xor \U$6897 ( \7240 , \6883 , \6892 );
xor \U$6898 ( \7241 , \7240 , \6895 );
and \U$6899 ( \7242 , \7239 , \7241 );
and \U$6900 ( \7243 , \7236 , \7238 );
or \U$6901 ( \7244 , \7242 , \7243 );
nand \U$6902 ( \7245 , \7234 , \7244 );
nand \U$6903 ( \7246 , \7231 , \7245 );
nand \U$6904 ( \7247 , \6938 , \7246 );
nand \U$6905 ( \7248 , \6937 , \7247 );
xor \U$6906 ( \7249 , \6374 , \6589 );
and \U$6907 ( \7250 , \7249 , \6625 );
and \U$6908 ( \7251 , \6374 , \6589 );
or \U$6909 ( \7252 , \7250 , \7251 );
xor \U$6910 ( \7253 , \5808 , \5810 );
xor \U$6911 ( \7254 , \7253 , \5823 );
xor \U$6912 ( \7255 , \7252 , \7254 );
xor \U$6913 ( \7256 , \6306 , \6320 );
xor \U$6914 ( \7257 , \7256 , \6325 );
and \U$6915 ( \7258 , \6630 , \7257 );
xor \U$6916 ( \7259 , \6306 , \6320 );
xor \U$6917 ( \7260 , \7259 , \6325 );
and \U$6918 ( \7261 , \6634 , \7260 );
and \U$6919 ( \7262 , \6630 , \6634 );
or \U$6920 ( \7263 , \7258 , \7261 , \7262 );
xor \U$6921 ( \7264 , \7255 , \7263 );
xor \U$6922 ( \7265 , \7248 , \7264 );
xor \U$6923 ( \7266 , \6901 , \6903 );
and \U$6924 ( \7267 , \7266 , \6934 );
and \U$6925 ( \7268 , \6901 , \6903 );
or \U$6926 ( \7269 , \7267 , \7268 );
and \U$6927 ( \7270 , \6626 , \6636 );
xor \U$6928 ( \7271 , \7269 , \7270 );
xor \U$6929 ( \7272 , \6333 , \6335 );
xor \U$6930 ( \7273 , \7272 , \6338 );
xor \U$6931 ( \7274 , \5920 , \5942 );
xor \U$6932 ( \7275 , \7274 , \6027 );
xor \U$6933 ( \7276 , \6082 , \6287 );
xor \U$6934 ( \7277 , \7276 , \6328 );
xor \U$6935 ( \7278 , \7275 , \7277 );
xor \U$6936 ( \7279 , \7273 , \7278 );
xor \U$6937 ( \7280 , \7271 , \7279 );
and \U$6938 ( \7281 , \7265 , \7280 );
and \U$6939 ( \7282 , \7248 , \7264 );
or \U$6940 ( \7283 , \7281 , \7282 );
not \U$6941 ( \7284 , \7283 );
xor \U$6942 ( \7285 , \7269 , \7270 );
and \U$6943 ( \7286 , \7285 , \7279 );
and \U$6944 ( \7287 , \7269 , \7270 );
or \U$6945 ( \7288 , \7286 , \7287 );
xor \U$6946 ( \7289 , \6331 , \6341 );
xor \U$6947 ( \7290 , \7289 , \6346 );
xor \U$6948 ( \7291 , \7288 , \7290 );
xor \U$6949 ( \7292 , \5826 , \6030 );
xor \U$6950 ( \7293 , \7292 , \6043 );
xor \U$6951 ( \7294 , \7252 , \7254 );
and \U$6952 ( \7295 , \7294 , \7263 );
and \U$6953 ( \7296 , \7252 , \7254 );
or \U$6954 ( \7297 , \7295 , \7296 );
xor \U$6955 ( \7298 , \7293 , \7297 );
xor \U$6956 ( \7299 , \6333 , \6335 );
xor \U$6957 ( \7300 , \7299 , \6338 );
and \U$6958 ( \7301 , \7275 , \7300 );
xor \U$6959 ( \7302 , \6333 , \6335 );
xor \U$6960 ( \7303 , \7302 , \6338 );
and \U$6961 ( \7304 , \7277 , \7303 );
and \U$6962 ( \7305 , \7275 , \7277 );
or \U$6963 ( \7306 , \7301 , \7304 , \7305 );
xor \U$6964 ( \7307 , \7298 , \7306 );
xor \U$6965 ( \7308 , \7291 , \7307 );
not \U$6966 ( \7309 , \7308 );
or \U$6967 ( \7310 , \7284 , \7309 );
xor \U$6968 ( \7311 , \6699 , \6721 );
xor \U$6969 ( \7312 , \7311 , \6750 );
xor \U$6970 ( \7313 , \6968 , \6994 );
xor \U$6971 ( \7314 , \7313 , \6999 );
and \U$6972 ( \7315 , \7312 , \7314 );
xor \U$6973 ( \7316 , \6812 , \6841 );
xor \U$6974 ( \7317 , \7316 , \6870 );
xor \U$6975 ( \7318 , \7215 , \7222 );
xor \U$6976 ( \7319 , \7317 , \7318 );
xor \U$6977 ( \7320 , \6968 , \6994 );
xor \U$6978 ( \7321 , \7320 , \6999 );
and \U$6979 ( \7322 , \7319 , \7321 );
and \U$6980 ( \7323 , \7312 , \7319 );
or \U$6981 ( \7324 , \7315 , \7322 , \7323 );
xor \U$6982 ( \7325 , \6650 , \6656 );
xor \U$6983 ( \7326 , \7325 , \6669 );
and \U$6984 ( \7327 , \7324 , \7326 );
not \U$6985 ( \7328 , \7324 );
not \U$6986 ( \7329 , \7326 );
and \U$6987 ( \7330 , \7328 , \7329 );
xor \U$6988 ( \7331 , \7071 , \7084 );
xor \U$6989 ( \7332 , \7331 , \7092 );
xor \U$6990 ( \7333 , \7044 , \7052 );
xor \U$6991 ( \7334 , \7333 , \7061 );
and \U$6992 ( \7335 , \7332 , \7334 );
xor \U$6993 ( \7336 , \7103 , \7111 );
xor \U$6994 ( \7337 , \7336 , \7119 );
xor \U$6995 ( \7338 , \7044 , \7052 );
xor \U$6996 ( \7339 , \7338 , \7061 );
and \U$6997 ( \7340 , \7337 , \7339 );
and \U$6998 ( \7341 , \7332 , \7337 );
or \U$6999 ( \7342 , \7335 , \7340 , \7341 );
xor \U$7000 ( \7343 , \6707 , \6710 );
xor \U$7001 ( \7344 , \7343 , \6718 );
xor \U$7002 ( \7345 , \7342 , \7344 );
xor \U$7003 ( \7346 , \7133 , \7141 );
xor \U$7004 ( \7347 , \7346 , \7149 );
xor \U$7005 ( \7348 , \7160 , \7167 );
xor \U$7006 ( \7349 , \7348 , \7176 );
and \U$7007 ( \7350 , \7347 , \7349 );
xor \U$7008 ( \7351 , \7187 , \7195 );
xor \U$7009 ( \7352 , \7351 , \7203 );
xor \U$7010 ( \7353 , \7160 , \7167 );
xor \U$7011 ( \7354 , \7353 , \7176 );
and \U$7012 ( \7355 , \7352 , \7354 );
and \U$7013 ( \7356 , \7347 , \7352 );
or \U$7014 ( \7357 , \7350 , \7355 , \7356 );
and \U$7015 ( \7358 , \7345 , \7357 );
and \U$7016 ( \7359 , \7342 , \7344 );
or \U$7017 ( \7360 , \7358 , \7359 );
and \U$7018 ( \7361 , \2464 , RI986e710_23);
and \U$7019 ( \7362 , RI986e620_21, \2462 );
nor \U$7020 ( \7363 , \7361 , \7362 );
and \U$7021 ( \7364 , \7363 , \2468 );
not \U$7022 ( \7365 , \7363 );
and \U$7023 ( \7366 , \7365 , \2263 );
nor \U$7024 ( \7367 , \7364 , \7366 );
not \U$7025 ( \7368 , \2034 );
and \U$7026 ( \7369 , \2042 , RI986f250_47);
and \U$7027 ( \7370 , RI986f160_45, \2040 );
nor \U$7028 ( \7371 , \7369 , \7370 );
not \U$7029 ( \7372 , \7371 );
or \U$7030 ( \7373 , \7368 , \7372 );
or \U$7031 ( \7374 , \7371 , \2034 );
nand \U$7032 ( \7375 , \7373 , \7374 );
xor \U$7033 ( \7376 , \7367 , \7375 );
and \U$7034 ( \7377 , \2274 , RI986e530_19);
and \U$7035 ( \7378 , RI986e440_17, \2272 );
nor \U$7036 ( \7379 , \7377 , \7378 );
and \U$7037 ( \7380 , \7379 , \2030 );
not \U$7038 ( \7381 , \7379 );
and \U$7039 ( \7382 , \7381 , \2031 );
nor \U$7040 ( \7383 , \7380 , \7382 );
and \U$7041 ( \7384 , \7376 , \7383 );
and \U$7042 ( \7385 , \7367 , \7375 );
or \U$7043 ( \7386 , \7384 , \7385 );
and \U$7044 ( \7387 , \438 , RI986ead0_31);
and \U$7045 ( \7388 , RI986e9e0_29, \436 );
nor \U$7046 ( \7389 , \7387 , \7388 );
and \U$7047 ( \7390 , \7389 , \444 );
not \U$7048 ( \7391 , \7389 );
and \U$7049 ( \7392 , \7391 , \443 );
nor \U$7050 ( \7393 , \7390 , \7392 );
and \U$7051 ( \7394 , \776 , RI986e8f0_27);
and \U$7052 ( \7395 , RI986e800_25, \774 );
nor \U$7053 ( \7396 , \7394 , \7395 );
and \U$7054 ( \7397 , \7396 , \474 );
not \U$7055 ( \7398 , \7396 );
and \U$7056 ( \7399 , \7398 , \451 );
nor \U$7057 ( \7400 , \7397 , \7399 );
xor \U$7058 ( \7401 , \7393 , \7400 );
not \U$7059 ( \7402 , \456 );
and \U$7060 ( \7403 , \465 , RI9871500_121);
and \U$7061 ( \7404 , RI98715f0_123, \463 );
nor \U$7062 ( \7405 , \7403 , \7404 );
not \U$7063 ( \7406 , \7405 );
or \U$7064 ( \7407 , \7402 , \7406 );
or \U$7065 ( \7408 , \7405 , \456 );
nand \U$7066 ( \7409 , \7407 , \7408 );
and \U$7067 ( \7410 , \7401 , \7409 );
and \U$7068 ( \7411 , \7393 , \7400 );
or \U$7069 ( \7412 , \7410 , \7411 );
xor \U$7070 ( \7413 , \7386 , \7412 );
and \U$7071 ( \7414 , \1329 , RI986ebc0_33);
and \U$7072 ( \7415 , RI986ecb0_35, \1327 );
nor \U$7073 ( \7416 , \7414 , \7415 );
and \U$7074 ( \7417 , \7416 , \1336 );
not \U$7075 ( \7418 , \7416 );
and \U$7076 ( \7419 , \7418 , \1337 );
nor \U$7077 ( \7420 , \7417 , \7419 );
not \U$7078 ( \7421 , \1128 );
and \U$7079 ( \7422 , \1293 , RI986ee90_39);
and \U$7080 ( \7423 , RI986eda0_37, \1291 );
nor \U$7081 ( \7424 , \7422 , \7423 );
not \U$7082 ( \7425 , \7424 );
or \U$7083 ( \7426 , \7421 , \7425 );
or \U$7084 ( \7427 , \7424 , \1128 );
nand \U$7085 ( \7428 , \7426 , \7427 );
xor \U$7086 ( \7429 , \7420 , \7428 );
and \U$7087 ( \7430 , \1311 , RI986f070_43);
and \U$7088 ( \7431 , RI986ef80_41, \1309 );
nor \U$7089 ( \7432 , \7430 , \7431 );
and \U$7090 ( \7433 , \7432 , \1458 );
not \U$7091 ( \7434 , \7432 );
and \U$7092 ( \7435 , \7434 , \1315 );
nor \U$7093 ( \7436 , \7433 , \7435 );
and \U$7094 ( \7437 , \7429 , \7436 );
and \U$7095 ( \7438 , \7420 , \7428 );
or \U$7096 ( \7439 , \7437 , \7438 );
and \U$7097 ( \7440 , \7413 , \7439 );
and \U$7098 ( \7441 , \7386 , \7412 );
or \U$7099 ( \7442 , \7440 , \7441 );
and \U$7100 ( \7443 , \4203 , RI986f430_51);
and \U$7101 ( \7444 , RI986f340_49, \4201 );
nor \U$7102 ( \7445 , \7443 , \7444 );
and \U$7103 ( \7446 , \7445 , \4207 );
not \U$7104 ( \7447 , \7445 );
and \U$7105 ( \7448 , \7447 , \3922 );
nor \U$7106 ( \7449 , \7446 , \7448 );
not \U$7107 ( \7450 , \3406 );
and \U$7108 ( \7451 , \3254 , RI986f7f0_59);
and \U$7109 ( \7452 , RI986f700_57, \3252 );
nor \U$7110 ( \7453 , \7451 , \7452 );
not \U$7111 ( \7454 , \7453 );
or \U$7112 ( \7455 , \7450 , \7454 );
or \U$7113 ( \7456 , \7453 , \3406 );
nand \U$7114 ( \7457 , \7455 , \7456 );
xor \U$7115 ( \7458 , \7449 , \7457 );
not \U$7116 ( \7459 , \3918 );
and \U$7117 ( \7460 , \3683 , RI986f9d0_63);
and \U$7118 ( \7461 , RI986f8e0_61, \3681 );
nor \U$7119 ( \7462 , \7460 , \7461 );
not \U$7120 ( \7463 , \7462 );
or \U$7121 ( \7464 , \7459 , \7463 );
or \U$7122 ( \7465 , \7462 , \3918 );
nand \U$7123 ( \7466 , \7464 , \7465 );
and \U$7124 ( \7467 , \7458 , \7466 );
and \U$7125 ( \7468 , \7449 , \7457 );
or \U$7126 ( \7469 , \7467 , \7468 );
and \U$7127 ( \7470 , \6453 , RI986e170_11);
and \U$7128 ( \7471 , RI986e080_9, \6451 );
nor \U$7129 ( \7472 , \7470 , \7471 );
and \U$7130 ( \7473 , \7472 , \6190 );
not \U$7131 ( \7474 , \7472 );
and \U$7132 ( \7475 , \7474 , \6705 );
nor \U$7133 ( \7476 , \7473 , \7475 );
not \U$7134 ( \7477 , RI9872d60_173);
not \U$7135 ( \7478 , RI9872ce8_172);
or \U$7136 ( \7479 , \7477 , \7478 );
nand \U$7137 ( \7480 , \7479 , RI9872bf8_170);
xor \U$7138 ( \7481 , \7476 , \7480 );
and \U$7139 ( \7482 , \7079 , RI986e260_13);
and \U$7140 ( \7483 , RI986e350_15, \7077 );
nor \U$7141 ( \7484 , \7482 , \7483 );
and \U$7142 ( \7485 , \7484 , \6710 );
not \U$7143 ( \7486 , \7484 );
and \U$7144 ( \7487 , \7486 , \6709 );
nor \U$7145 ( \7488 , \7485 , \7487 );
and \U$7146 ( \7489 , \7481 , \7488 );
and \U$7147 ( \7490 , \7476 , \7480 );
or \U$7148 ( \7491 , \7489 , \7490 );
xor \U$7149 ( \7492 , \7469 , \7491 );
and \U$7150 ( \7493 , \5318 , RI986df90_7);
and \U$7151 ( \7494 , RI986dea0_5, \5316 );
nor \U$7152 ( \7495 , \7493 , \7494 );
and \U$7153 ( \7496 , \7495 , \5052 );
not \U$7154 ( \7497 , \7495 );
and \U$7155 ( \7498 , \7497 , \5322 );
nor \U$7156 ( \7499 , \7496 , \7498 );
not \U$7157 ( \7500 , \4519 );
and \U$7158 ( \7501 , \4710 , RI986f520_53);
and \U$7159 ( \7502 , RI986f610_55, \4708 );
nor \U$7160 ( \7503 , \7501 , \7502 );
not \U$7161 ( \7504 , \7503 );
or \U$7162 ( \7505 , \7500 , \7504 );
or \U$7163 ( \7506 , \7503 , \4521 );
nand \U$7164 ( \7507 , \7505 , \7506 );
xor \U$7165 ( \7508 , \7499 , \7507 );
and \U$7166 ( \7509 , \5881 , RI986ddb0_3);
and \U$7167 ( \7510 , RI986dcc0_1, \5879 );
nor \U$7168 ( \7511 , \7509 , \7510 );
and \U$7169 ( \7512 , \7511 , \5594 );
not \U$7170 ( \7513 , \7511 );
and \U$7171 ( \7514 , \7513 , \5885 );
nor \U$7172 ( \7515 , \7512 , \7514 );
and \U$7173 ( \7516 , \7508 , \7515 );
and \U$7174 ( \7517 , \7499 , \7507 );
or \U$7175 ( \7518 , \7516 , \7517 );
and \U$7176 ( \7519 , \7492 , \7518 );
and \U$7177 ( \7520 , \7469 , \7491 );
or \U$7178 ( \7521 , \7519 , \7520 );
xor \U$7179 ( \7522 , \7442 , \7521 );
not \U$7180 ( \7523 , \345 );
and \U$7181 ( \7524 , \354 , RI9871230_115);
and \U$7182 ( \7525 , RI9871140_113, \352 );
nor \U$7183 ( \7526 , \7524 , \7525 );
not \U$7184 ( \7527 , \7526 );
or \U$7185 ( \7528 , \7523 , \7527 );
or \U$7186 ( \7529 , \7526 , \345 );
nand \U$7187 ( \7530 , \7528 , \7529 );
not \U$7188 ( \7531 , \367 );
and \U$7189 ( \7532 , \376 , RI98716e0_125);
and \U$7190 ( \7533 , RI98717d0_127, \374 );
nor \U$7191 ( \7534 , \7532 , \7533 );
not \U$7192 ( \7535 , \7534 );
or \U$7193 ( \7536 , \7531 , \7535 );
or \U$7194 ( \7537 , \7534 , \365 );
nand \U$7195 ( \7538 , \7536 , \7537 );
xor \U$7196 ( \7539 , \7530 , \7538 );
not \U$7197 ( \7540 , \386 );
and \U$7198 ( \7541 , \395 , RI9871320_117);
and \U$7199 ( \7542 , RI9871410_119, \393 );
nor \U$7200 ( \7543 , \7541 , \7542 );
not \U$7201 ( \7544 , \7543 );
or \U$7202 ( \7545 , \7540 , \7544 );
or \U$7203 ( \7546 , \7543 , \487 );
nand \U$7204 ( \7547 , \7545 , \7546 );
and \U$7205 ( \7548 , \7539 , \7547 );
and \U$7206 ( \7549 , \7530 , \7538 );
or \U$7207 ( \7550 , \7548 , \7549 );
xor \U$7208 ( \7551 , \7550 , \7003 );
not \U$7209 ( \7552 , \7021 );
xor \U$7210 ( \7553 , \7013 , \7032 );
not \U$7211 ( \7554 , \7553 );
or \U$7212 ( \7555 , \7552 , \7554 );
or \U$7213 ( \7556 , \7553 , \7021 );
nand \U$7214 ( \7557 , \7555 , \7556 );
and \U$7215 ( \7558 , \7551 , \7557 );
and \U$7216 ( \7559 , \7550 , \7003 );
or \U$7217 ( \7560 , \7558 , \7559 );
and \U$7218 ( \7561 , \7522 , \7560 );
and \U$7219 ( \7562 , \7442 , \7521 );
or \U$7220 ( \7563 , \7561 , \7562 );
and \U$7221 ( \7564 , \7360 , \7563 );
not \U$7222 ( \7565 , \7360 );
not \U$7223 ( \7566 , \7563 );
and \U$7224 ( \7567 , \7565 , \7566 );
not \U$7225 ( \7568 , \6950 );
not \U$7226 ( \7569 , \6966 );
or \U$7227 ( \7570 , \7568 , \7569 );
or \U$7228 ( \7571 , \6950 , \6966 );
nand \U$7229 ( \7572 , \7570 , \7571 );
not \U$7230 ( \7573 , \7572 );
not \U$7231 ( \7574 , \6960 );
and \U$7232 ( \7575 , \7573 , \7574 );
and \U$7233 ( \7576 , \7572 , \6960 );
nor \U$7234 ( \7577 , \7575 , \7576 );
xor \U$7235 ( \7578 , \7003 , \7004 );
xor \U$7236 ( \7579 , \7578 , \7034 );
xor \U$7237 ( \7580 , \7577 , \7579 );
xor \U$7238 ( \7581 , \6978 , \6988 );
xor \U$7239 ( \7582 , \7581 , \6991 );
and \U$7240 ( \7583 , \7580 , \7582 );
and \U$7241 ( \7584 , \7577 , \7579 );
or \U$7242 ( \7585 , \7583 , \7584 );
nor \U$7243 ( \7586 , \7567 , \7585 );
nor \U$7244 ( \7587 , \7564 , \7586 );
nor \U$7245 ( \7588 , \7330 , \7587 );
nor \U$7246 ( \7589 , \7327 , \7588 );
xor \U$7247 ( \7590 , \6672 , \6876 );
xor \U$7248 ( \7591 , \7590 , \6898 );
not \U$7249 ( \7592 , \7591 );
or \U$7250 ( \7593 , \7589 , \7592 );
not \U$7251 ( \7594 , \7592 );
not \U$7252 ( \7595 , \7589 );
or \U$7253 ( \7596 , \7594 , \7595 );
xor \U$7254 ( \7597 , \6753 , \6783 );
xor \U$7255 ( \7598 , \7597 , \6873 );
xor \U$7256 ( \7599 , \7236 , \7238 );
xor \U$7257 ( \7600 , \7599 , \7241 );
and \U$7258 ( \7601 , \7598 , \7600 );
xor \U$7259 ( \7602 , \7002 , \7212 );
xor \U$7260 ( \7603 , \7602 , \7227 );
xor \U$7261 ( \7604 , \7236 , \7238 );
xor \U$7262 ( \7605 , \7604 , \7241 );
and \U$7263 ( \7606 , \7603 , \7605 );
and \U$7264 ( \7607 , \7598 , \7603 );
or \U$7265 ( \7608 , \7601 , \7606 , \7607 );
nand \U$7266 ( \7609 , \7596 , \7608 );
nand \U$7267 ( \7610 , \7593 , \7609 );
not \U$7268 ( \7611 , \7610 );
not \U$7269 ( \7612 , \7589 );
not \U$7270 ( \7613 , \7608 );
and \U$7271 ( \7614 , \7612 , \7613 );
and \U$7272 ( \7615 , \7589 , \7608 );
nor \U$7273 ( \7616 , \7614 , \7615 );
not \U$7274 ( \7617 , \7616 );
not \U$7275 ( \7618 , \7591 );
and \U$7276 ( \7619 , \7617 , \7618 );
and \U$7277 ( \7620 , \7616 , \7591 );
nor \U$7278 ( \7621 , \7619 , \7620 );
not \U$7279 ( \7622 , \7244 );
not \U$7280 ( \7623 , \7230 );
or \U$7281 ( \7624 , \7622 , \7623 );
or \U$7282 ( \7625 , \7230 , \7244 );
nand \U$7283 ( \7626 , \7624 , \7625 );
not \U$7284 ( \7627 , \7626 );
not \U$7285 ( \7628 , \6940 );
and \U$7286 ( \7629 , \7627 , \7628 );
and \U$7287 ( \7630 , \7626 , \6940 );
nor \U$7288 ( \7631 , \7629 , \7630 );
xor \U$7289 ( \7632 , \7621 , \7631 );
xor \U$7290 ( \7633 , \7236 , \7238 );
xor \U$7291 ( \7634 , \7633 , \7241 );
xor \U$7292 ( \7635 , \7598 , \7603 );
xor \U$7293 ( \7636 , \7634 , \7635 );
not \U$7294 ( \7637 , \7587 );
not \U$7295 ( \7638 , \7324 );
or \U$7296 ( \7639 , \7637 , \7638 );
or \U$7297 ( \7640 , \7324 , \7587 );
nand \U$7298 ( \7641 , \7639 , \7640 );
xor \U$7299 ( \7642 , \7326 , \7641 );
and \U$7300 ( \7643 , \7636 , \7642 );
not \U$7301 ( \7644 , \7636 );
not \U$7302 ( \7645 , \7642 );
and \U$7303 ( \7646 , \7644 , \7645 );
xor \U$7304 ( \7647 , \7367 , \7375 );
xor \U$7305 ( \7648 , \7647 , \7383 );
xor \U$7306 ( \7649 , \7420 , \7428 );
xor \U$7307 ( \7650 , \7649 , \7436 );
and \U$7308 ( \7651 , \7648 , \7650 );
xor \U$7309 ( \7652 , \7449 , \7457 );
xor \U$7310 ( \7653 , \7652 , \7466 );
xor \U$7311 ( \7654 , \7420 , \7428 );
xor \U$7312 ( \7655 , \7654 , \7436 );
and \U$7313 ( \7656 , \7653 , \7655 );
and \U$7314 ( \7657 , \7648 , \7653 );
or \U$7315 ( \7658 , \7651 , \7656 , \7657 );
xor \U$7316 ( \7659 , \7530 , \7538 );
xor \U$7317 ( \7660 , \7659 , \7547 );
not \U$7318 ( \7661 , RI9870ba0_101);
nor \U$7319 ( \7662 , \7661 , \407 );
xor \U$7320 ( \7663 , \7660 , \7662 );
xor \U$7321 ( \7664 , \7393 , \7400 );
xor \U$7322 ( \7665 , \7664 , \7409 );
and \U$7323 ( \7666 , \7663 , \7665 );
and \U$7324 ( \7667 , \7660 , \7662 );
or \U$7325 ( \7668 , \7666 , \7667 );
xor \U$7326 ( \7669 , \7658 , \7668 );
xor \U$7327 ( \7670 , \7044 , \7052 );
xor \U$7328 ( \7671 , \7670 , \7061 );
xor \U$7329 ( \7672 , \7332 , \7337 );
xor \U$7330 ( \7673 , \7671 , \7672 );
and \U$7331 ( \7674 , \7669 , \7673 );
and \U$7332 ( \7675 , \7658 , \7668 );
or \U$7333 ( \7676 , \7674 , \7675 );
and \U$7334 ( \7677 , \4203 , RI986f8e0_61);
and \U$7335 ( \7678 , RI986f430_51, \4201 );
nor \U$7336 ( \7679 , \7677 , \7678 );
and \U$7337 ( \7680 , \7679 , \4207 );
not \U$7338 ( \7681 , \7679 );
and \U$7339 ( \7682 , \7681 , \3923 );
nor \U$7340 ( \7683 , \7680 , \7682 );
not \U$7341 ( \7684 , \2935 );
and \U$7342 ( \7685 , \3254 , RI986e620_21);
and \U$7343 ( \7686 , RI986f7f0_59, \3252 );
nor \U$7344 ( \7687 , \7685 , \7686 );
not \U$7345 ( \7688 , \7687 );
or \U$7346 ( \7689 , \7684 , \7688 );
or \U$7347 ( \7690 , \7687 , \2935 );
nand \U$7348 ( \7691 , \7689 , \7690 );
xor \U$7349 ( \7692 , \7683 , \7691 );
not \U$7350 ( \7693 , \3918 );
and \U$7351 ( \7694 , \3683 , RI986f700_57);
and \U$7352 ( \7695 , RI986f9d0_63, \3681 );
nor \U$7353 ( \7696 , \7694 , \7695 );
not \U$7354 ( \7697 , \7696 );
or \U$7355 ( \7698 , \7693 , \7697 );
or \U$7356 ( \7699 , \7696 , \3412 );
nand \U$7357 ( \7700 , \7698 , \7699 );
and \U$7358 ( \7701 , \7692 , \7700 );
and \U$7359 ( \7702 , \7683 , \7691 );
or \U$7360 ( \7703 , \7701 , \7702 );
and \U$7361 ( \7704 , \6453 , RI986dcc0_1);
and \U$7362 ( \7705 , RI986e170_11, \6451 );
nor \U$7363 ( \7706 , \7704 , \7705 );
and \U$7364 ( \7707 , \7706 , \6180 );
not \U$7365 ( \7708 , \7706 );
and \U$7366 ( \7709 , \7708 , \6190 );
nor \U$7367 ( \7710 , \7707 , \7709 );
and \U$7368 ( \7711 , \7079 , RI986e080_9);
and \U$7369 ( \7712 , RI986e260_13, \7077 );
nor \U$7370 ( \7713 , \7711 , \7712 );
and \U$7371 ( \7714 , \7713 , \6709 );
not \U$7372 ( \7715 , \7713 );
and \U$7373 ( \7716 , \7715 , \6710 );
nor \U$7374 ( \7717 , \7714 , \7716 );
or \U$7375 ( \7718 , \7710 , \7717 );
not \U$7376 ( \7719 , \7717 );
not \U$7377 ( \7720 , \7710 );
or \U$7378 ( \7721 , \7719 , \7720 );
and \U$7379 ( \7722 , RI9872bf8_170, RI9872ce8_172);
not \U$7380 ( \7723 , RI9872ce8_172);
nor \U$7381 ( \7724 , \7723 , RI9872d60_173);
not \U$7382 ( \7725 , RI9872d60_173);
nor \U$7383 ( \7726 , \7725 , RI9872ce8_172);
or \U$7384 ( \7727 , \7724 , \7726 );
nor \U$7385 ( \7728 , RI9872bf8_170, RI9872ce8_172);
nor \U$7386 ( \7729 , \7722 , \7727 , \7728 );
nand \U$7387 ( \7730 , RI986e350_15, \7729 );
and \U$7388 ( \7731 , \7730 , \7480 );
not \U$7389 ( \7732 , \7730 );
not \U$7390 ( \7733 , \7480 );
and \U$7391 ( \7734 , \7732 , \7733 );
nor \U$7392 ( \7735 , \7731 , \7734 );
nand \U$7393 ( \7736 , \7721 , \7735 );
nand \U$7394 ( \7737 , \7718 , \7736 );
xor \U$7395 ( \7738 , \7703 , \7737 );
and \U$7396 ( \7739 , \5881 , RI986dea0_5);
and \U$7397 ( \7740 , RI986ddb0_3, \5879 );
nor \U$7398 ( \7741 , \7739 , \7740 );
and \U$7399 ( \7742 , \7741 , \5594 );
not \U$7400 ( \7743 , \7741 );
and \U$7401 ( \7744 , \7743 , \5885 );
nor \U$7402 ( \7745 , \7742 , \7744 );
not \U$7403 ( \7746 , \4519 );
and \U$7404 ( \7747 , \4710 , RI986f340_49);
and \U$7405 ( \7748 , RI986f520_53, \4708 );
nor \U$7406 ( \7749 , \7747 , \7748 );
not \U$7407 ( \7750 , \7749 );
or \U$7408 ( \7751 , \7746 , \7750 );
or \U$7409 ( \7752 , \7749 , \4519 );
nand \U$7410 ( \7753 , \7751 , \7752 );
xor \U$7411 ( \7754 , \7745 , \7753 );
and \U$7412 ( \7755 , \5318 , RI986f610_55);
and \U$7413 ( \7756 , RI986df90_7, \5316 );
nor \U$7414 ( \7757 , \7755 , \7756 );
and \U$7415 ( \7758 , \7757 , \5052 );
not \U$7416 ( \7759 , \7757 );
and \U$7417 ( \7760 , \7759 , \5322 );
nor \U$7418 ( \7761 , \7758 , \7760 );
and \U$7419 ( \7762 , \7754 , \7761 );
and \U$7420 ( \7763 , \7745 , \7753 );
or \U$7421 ( \7764 , \7762 , \7763 );
and \U$7422 ( \7765 , \7738 , \7764 );
and \U$7423 ( \7766 , \7703 , \7737 );
or \U$7424 ( \7767 , \7765 , \7766 );
nand \U$7425 ( \7768 , RI9870e70_107, RI9871fc8_144);
and \U$7426 ( \7769 , \416 , RI9870ba0_101);
and \U$7427 ( \7770 , RI9871050_111, \414 );
nor \U$7428 ( \7771 , \7769 , \7770 );
and \U$7429 ( \7772 , \7771 , \421 );
not \U$7430 ( \7773 , \7771 );
and \U$7431 ( \7774 , \7773 , \422 );
nor \U$7432 ( \7775 , \7772 , \7774 );
nand \U$7433 ( \7776 , \7768 , \7775 );
and \U$7434 ( \7777 , \416 , RI9871050_111);
and \U$7435 ( \7778 , RI9870c90_103, \414 );
nor \U$7436 ( \7779 , \7777 , \7778 );
and \U$7437 ( \7780 , \7779 , \422 );
not \U$7438 ( \7781 , \7779 );
and \U$7439 ( \7782 , \7781 , \421 );
nor \U$7440 ( \7783 , \7780 , \7782 );
xor \U$7441 ( \7784 , \7776 , \7783 );
not \U$7442 ( \7785 , \365 );
and \U$7443 ( \7786 , \376 , RI9871410_119);
and \U$7444 ( \7787 , RI98716e0_125, \374 );
nor \U$7445 ( \7788 , \7786 , \7787 );
not \U$7446 ( \7789 , \7788 );
or \U$7447 ( \7790 , \7785 , \7789 );
or \U$7448 ( \7791 , \7788 , \365 );
nand \U$7449 ( \7792 , \7790 , \7791 );
not \U$7450 ( \7793 , \386 );
and \U$7451 ( \7794 , \395 , RI9871140_113);
and \U$7452 ( \7795 , RI9871320_117, \393 );
nor \U$7453 ( \7796 , \7794 , \7795 );
not \U$7454 ( \7797 , \7796 );
or \U$7455 ( \7798 , \7793 , \7797 );
or \U$7456 ( \7799 , \7796 , \487 );
nand \U$7457 ( \7800 , \7798 , \7799 );
xor \U$7458 ( \7801 , \7792 , \7800 );
not \U$7459 ( \7802 , \345 );
and \U$7460 ( \7803 , \354 , RI9870c90_103);
and \U$7461 ( \7804 , RI9871230_115, \352 );
nor \U$7462 ( \7805 , \7803 , \7804 );
not \U$7463 ( \7806 , \7805 );
or \U$7464 ( \7807 , \7802 , \7806 );
or \U$7465 ( \7808 , \7805 , \361 );
nand \U$7466 ( \7809 , \7807 , \7808 );
and \U$7467 ( \7810 , \7801 , \7809 );
and \U$7468 ( \7811 , \7792 , \7800 );
or \U$7469 ( \7812 , \7810 , \7811 );
and \U$7470 ( \7813 , \7784 , \7812 );
and \U$7471 ( \7814 , \7776 , \7783 );
or \U$7472 ( \7815 , \7813 , \7814 );
xor \U$7473 ( \7816 , \7767 , \7815 );
and \U$7474 ( \7817 , \2464 , RI986e440_17);
and \U$7475 ( \7818 , RI986e710_23, \2462 );
nor \U$7476 ( \7819 , \7817 , \7818 );
and \U$7477 ( \7820 , \7819 , \2468 );
not \U$7478 ( \7821 , \7819 );
and \U$7479 ( \7822 , \7821 , \2263 );
nor \U$7480 ( \7823 , \7820 , \7822 );
not \U$7481 ( \7824 , \1462 );
and \U$7482 ( \7825 , \2042 , RI986ef80_41);
and \U$7483 ( \7826 , RI986f250_47, \2040 );
nor \U$7484 ( \7827 , \7825 , \7826 );
not \U$7485 ( \7828 , \7827 );
or \U$7486 ( \7829 , \7824 , \7828 );
or \U$7487 ( \7830 , \7827 , \2034 );
nand \U$7488 ( \7831 , \7829 , \7830 );
xor \U$7489 ( \7832 , \7823 , \7831 );
and \U$7490 ( \7833 , \2274 , RI986f160_45);
and \U$7491 ( \7834 , RI986e530_19, \2272 );
nor \U$7492 ( \7835 , \7833 , \7834 );
and \U$7493 ( \7836 , \7835 , \2030 );
not \U$7494 ( \7837 , \7835 );
and \U$7495 ( \7838 , \7837 , \2031 );
nor \U$7496 ( \7839 , \7836 , \7838 );
and \U$7497 ( \7840 , \7832 , \7839 );
and \U$7498 ( \7841 , \7823 , \7831 );
or \U$7499 ( \7842 , \7840 , \7841 );
and \U$7500 ( \7843 , \1293 , RI986e800_25);
and \U$7501 ( \7844 , RI986ee90_39, \1291 );
nor \U$7502 ( \7845 , \7843 , \7844 );
not \U$7503 ( \7846 , \7845 );
not \U$7504 ( \7847 , \1128 );
and \U$7505 ( \7848 , \7846 , \7847 );
and \U$7506 ( \7849 , \7845 , \1128 );
nor \U$7507 ( \7850 , \7848 , \7849 );
and \U$7508 ( \7851 , \1329 , RI986eda0_37);
and \U$7509 ( \7852 , RI986ebc0_33, \1327 );
nor \U$7510 ( \7853 , \7851 , \7852 );
and \U$7511 ( \7854 , \7853 , \1337 );
not \U$7512 ( \7855 , \7853 );
and \U$7513 ( \7856 , \7855 , \1336 );
nor \U$7514 ( \7857 , \7854 , \7856 );
or \U$7515 ( \7858 , \7850 , \7857 );
not \U$7516 ( \7859 , \7857 );
not \U$7517 ( \7860 , \7850 );
or \U$7518 ( \7861 , \7859 , \7860 );
and \U$7519 ( \7862 , \1311 , RI986ecb0_35);
and \U$7520 ( \7863 , RI986f070_43, \1309 );
nor \U$7521 ( \7864 , \7862 , \7863 );
and \U$7522 ( \7865 , \7864 , \1458 );
not \U$7523 ( \7866 , \7864 );
and \U$7524 ( \7867 , \7866 , \1315 );
nor \U$7525 ( \7868 , \7865 , \7867 );
nand \U$7526 ( \7869 , \7861 , \7868 );
nand \U$7527 ( \7870 , \7858 , \7869 );
xor \U$7528 ( \7871 , \7842 , \7870 );
and \U$7529 ( \7872 , \438 , RI98715f0_123);
and \U$7530 ( \7873 , RI986ead0_31, \436 );
nor \U$7531 ( \7874 , \7872 , \7873 );
and \U$7532 ( \7875 , \7874 , \443 );
not \U$7533 ( \7876 , \7874 );
and \U$7534 ( \7877 , \7876 , \444 );
nor \U$7535 ( \7878 , \7875 , \7877 );
and \U$7536 ( \7879 , \465 , RI98717d0_127);
and \U$7537 ( \7880 , RI9871500_121, \463 );
nor \U$7538 ( \7881 , \7879 , \7880 );
not \U$7539 ( \7882 , \7881 );
not \U$7540 ( \7883 , \456 );
and \U$7541 ( \7884 , \7882 , \7883 );
and \U$7542 ( \7885 , \7881 , \454 );
nor \U$7543 ( \7886 , \7884 , \7885 );
or \U$7544 ( \7887 , \7878 , \7886 );
not \U$7545 ( \7888 , \7886 );
not \U$7546 ( \7889 , \7878 );
or \U$7547 ( \7890 , \7888 , \7889 );
and \U$7548 ( \7891 , \776 , RI986e9e0_29);
and \U$7549 ( \7892 , RI986e8f0_27, \774 );
nor \U$7550 ( \7893 , \7891 , \7892 );
and \U$7551 ( \7894 , \7893 , \474 );
not \U$7552 ( \7895 , \7893 );
and \U$7553 ( \7896 , \7895 , \451 );
nor \U$7554 ( \7897 , \7894 , \7896 );
nand \U$7555 ( \7898 , \7890 , \7897 );
nand \U$7556 ( \7899 , \7887 , \7898 );
and \U$7557 ( \7900 , \7871 , \7899 );
and \U$7558 ( \7901 , \7842 , \7870 );
or \U$7559 ( \7902 , \7900 , \7901 );
and \U$7560 ( \7903 , \7816 , \7902 );
and \U$7561 ( \7904 , \7767 , \7815 );
or \U$7562 ( \7905 , \7903 , \7904 );
xor \U$7563 ( \7906 , \7676 , \7905 );
xor \U$7564 ( \7907 , \7386 , \7412 );
xor \U$7565 ( \7908 , \7907 , \7439 );
xor \U$7566 ( \7909 , \7550 , \7003 );
xor \U$7567 ( \7910 , \7909 , \7557 );
and \U$7568 ( \7911 , \7908 , \7910 );
xor \U$7569 ( \7912 , \7160 , \7167 );
xor \U$7570 ( \7913 , \7912 , \7176 );
xor \U$7571 ( \7914 , \7347 , \7352 );
xor \U$7572 ( \7915 , \7913 , \7914 );
xor \U$7573 ( \7916 , \7550 , \7003 );
xor \U$7574 ( \7917 , \7916 , \7557 );
and \U$7575 ( \7918 , \7915 , \7917 );
and \U$7576 ( \7919 , \7908 , \7915 );
or \U$7577 ( \7920 , \7911 , \7918 , \7919 );
and \U$7578 ( \7921 , \7906 , \7920 );
and \U$7579 ( \7922 , \7676 , \7905 );
nor \U$7580 ( \7923 , \7921 , \7922 );
not \U$7581 ( \7924 , \7923 );
xor \U$7582 ( \7925 , \7037 , \7125 );
xor \U$7583 ( \7926 , \7925 , \7209 );
not \U$7584 ( \7927 , \7926 );
and \U$7585 ( \7928 , \7924 , \7927 );
and \U$7586 ( \7929 , \7923 , \7926 );
xor \U$7587 ( \7930 , \7152 , \7179 );
xor \U$7588 ( \7931 , \7930 , \7206 );
xor \U$7589 ( \7932 , \7064 , \7095 );
xor \U$7590 ( \7933 , \7932 , \7122 );
and \U$7591 ( \7934 , \7931 , \7933 );
not \U$7592 ( \7935 , \7933 );
not \U$7593 ( \7936 , \7931 );
and \U$7594 ( \7937 , \7935 , \7936 );
xor \U$7595 ( \7938 , \7577 , \7579 );
xor \U$7596 ( \7939 , \7938 , \7582 );
nor \U$7597 ( \7940 , \7937 , \7939 );
nor \U$7598 ( \7941 , \7934 , \7940 );
nor \U$7599 ( \7942 , \7929 , \7941 );
nor \U$7600 ( \7943 , \7928 , \7942 );
nor \U$7601 ( \7944 , \7646 , \7943 );
nor \U$7602 ( \7945 , \7643 , \7944 );
and \U$7603 ( \7946 , \7632 , \7945 );
and \U$7604 ( \7947 , \7621 , \7631 );
or \U$7605 ( \7948 , \7946 , \7947 );
not \U$7606 ( \7949 , \7948 );
or \U$7607 ( \7950 , \7611 , \7949 );
or \U$7608 ( \7951 , \7948 , \7610 );
nand \U$7609 ( \7952 , \7950 , \7951 );
not \U$7610 ( \7953 , \7952 );
xnor \U$7611 ( \7954 , \7246 , \6935 );
not \U$7612 ( \7955 , \7954 );
not \U$7613 ( \7956 , \6637 );
and \U$7614 ( \7957 , \7955 , \7956 );
and \U$7615 ( \7958 , \7954 , \6637 );
nor \U$7616 ( \7959 , \7957 , \7958 );
not \U$7617 ( \7960 , \7959 );
and \U$7618 ( \7961 , \7953 , \7960 );
and \U$7619 ( \7962 , \7952 , \7959 );
nor \U$7620 ( \7963 , \7961 , \7962 );
xor \U$7621 ( \7964 , \7621 , \7631 );
xor \U$7622 ( \7965 , \7964 , \7945 );
not \U$7623 ( \7966 , \7965 );
xor \U$7624 ( \7967 , \7683 , \7691 );
xor \U$7625 ( \7968 , \7967 , \7700 );
xor \U$7626 ( \7969 , \7823 , \7831 );
xor \U$7627 ( \7970 , \7969 , \7839 );
and \U$7628 ( \7971 , \7968 , \7970 );
xor \U$7629 ( \7972 , \7745 , \7753 );
xor \U$7630 ( \7973 , \7972 , \7761 );
xor \U$7631 ( \7974 , \7823 , \7831 );
xor \U$7632 ( \7975 , \7974 , \7839 );
and \U$7633 ( \7976 , \7973 , \7975 );
and \U$7634 ( \7977 , \7968 , \7973 );
or \U$7635 ( \7978 , \7971 , \7976 , \7977 );
xor \U$7636 ( \7979 , \7499 , \7507 );
xor \U$7637 ( \7980 , \7979 , \7515 );
xor \U$7638 ( \7981 , \7978 , \7980 );
not \U$7639 ( \7982 , \7878 );
not \U$7640 ( \7983 , \7897 );
or \U$7641 ( \7984 , \7982 , \7983 );
or \U$7642 ( \7985 , \7878 , \7897 );
nand \U$7643 ( \7986 , \7984 , \7985 );
not \U$7644 ( \7987 , \7986 );
not \U$7645 ( \7988 , \7886 );
and \U$7646 ( \7989 , \7987 , \7988 );
and \U$7647 ( \7990 , \7986 , \7886 );
nor \U$7648 ( \7991 , \7989 , \7990 );
not \U$7649 ( \7992 , \7857 );
not \U$7650 ( \7993 , \7868 );
or \U$7651 ( \7994 , \7992 , \7993 );
or \U$7652 ( \7995 , \7857 , \7868 );
nand \U$7653 ( \7996 , \7994 , \7995 );
not \U$7654 ( \7997 , \7996 );
not \U$7655 ( \7998 , \7850 );
and \U$7656 ( \7999 , \7997 , \7998 );
and \U$7657 ( \8000 , \7996 , \7850 );
nor \U$7658 ( \8001 , \7999 , \8000 );
or \U$7659 ( \8002 , \7991 , \8001 );
not \U$7660 ( \8003 , \8001 );
not \U$7661 ( \8004 , \7991 );
or \U$7662 ( \8005 , \8003 , \8004 );
xor \U$7663 ( \8006 , \7792 , \7800 );
xor \U$7664 ( \8007 , \8006 , \7809 );
nand \U$7665 ( \8008 , \8005 , \8007 );
nand \U$7666 ( \8009 , \8002 , \8008 );
and \U$7667 ( \8010 , \7981 , \8009 );
and \U$7668 ( \8011 , \7978 , \7980 );
or \U$7669 ( \8012 , \8010 , \8011 );
and \U$7670 ( \8013 , \3683 , RI986f7f0_59);
and \U$7671 ( \8014 , RI986f700_57, \3681 );
nor \U$7672 ( \8015 , \8013 , \8014 );
not \U$7673 ( \8016 , \8015 );
not \U$7674 ( \8017 , \3412 );
and \U$7675 ( \8018 , \8016 , \8017 );
and \U$7676 ( \8019 , \8015 , \3412 );
nor \U$7677 ( \8020 , \8018 , \8019 );
and \U$7678 ( \8021 , \4203 , RI986f9d0_63);
and \U$7679 ( \8022 , RI986f8e0_61, \4201 );
nor \U$7680 ( \8023 , \8021 , \8022 );
and \U$7681 ( \8024 , \8023 , \3922 );
not \U$7682 ( \8025 , \8023 );
and \U$7683 ( \8026 , \8025 , \4207 );
nor \U$7684 ( \8027 , \8024 , \8026 );
xor \U$7685 ( \8028 , \8020 , \8027 );
and \U$7686 ( \8029 , \4710 , RI986f430_51);
and \U$7687 ( \8030 , RI986f340_49, \4708 );
nor \U$7688 ( \8031 , \8029 , \8030 );
not \U$7689 ( \8032 , \8031 );
not \U$7690 ( \8033 , \4519 );
and \U$7691 ( \8034 , \8032 , \8033 );
and \U$7692 ( \8035 , \8031 , \4519 );
nor \U$7693 ( \8036 , \8034 , \8035 );
and \U$7694 ( \8037 , \8028 , \8036 );
and \U$7695 ( \8038 , \8020 , \8027 );
or \U$7696 ( \8039 , \8037 , \8038 );
and \U$7697 ( \8040 , \7079 , RI986e170_11);
and \U$7698 ( \8041 , RI986e080_9, \7077 );
nor \U$7699 ( \8042 , \8040 , \8041 );
and \U$7700 ( \8043 , \8042 , \6709 );
not \U$7701 ( \8044 , \8042 );
and \U$7702 ( \8045 , \8044 , \6710 );
nor \U$7703 ( \8046 , \8043 , \8045 );
not \U$7704 ( \8047 , RI9872e50_175);
not \U$7705 ( \8048 , RI9872dd8_174);
or \U$7706 ( \8049 , \8047 , \8048 );
nand \U$7707 ( \8050 , \8049 , RI9872d60_173);
not \U$7708 ( \8051 , \8050 );
xor \U$7709 ( \8052 , \8046 , \8051 );
and \U$7710 ( \8053 , \7729 , RI986e260_13);
and \U$7711 ( \8054 , RI986e350_15, \7727 );
nor \U$7712 ( \8055 , \8053 , \8054 );
and \U$7713 ( \8056 , \8055 , \7733 );
not \U$7714 ( \8057 , \8055 );
and \U$7715 ( \8058 , \8057 , \7480 );
nor \U$7716 ( \8059 , \8056 , \8058 );
and \U$7717 ( \8060 , \8052 , \8059 );
and \U$7718 ( \8061 , \8046 , \8051 );
or \U$7719 ( \8062 , \8060 , \8061 );
xor \U$7720 ( \8063 , \8039 , \8062 );
and \U$7721 ( \8064 , \5881 , RI986df90_7);
and \U$7722 ( \8065 , RI986dea0_5, \5879 );
nor \U$7723 ( \8066 , \8064 , \8065 );
and \U$7724 ( \8067 , \8066 , \5885 );
not \U$7725 ( \8068 , \8066 );
and \U$7726 ( \8069 , \8068 , \5594 );
nor \U$7727 ( \8070 , \8067 , \8069 );
and \U$7728 ( \8071 , \5318 , RI986f520_53);
and \U$7729 ( \8072 , RI986f610_55, \5316 );
nor \U$7730 ( \8073 , \8071 , \8072 );
and \U$7731 ( \8074 , \8073 , \5322 );
not \U$7732 ( \8075 , \8073 );
and \U$7733 ( \8076 , \8075 , \5052 );
nor \U$7734 ( \8077 , \8074 , \8076 );
xor \U$7735 ( \8078 , \8070 , \8077 );
and \U$7736 ( \8079 , \6453 , RI986ddb0_3);
and \U$7737 ( \8080 , RI986dcc0_1, \6451 );
nor \U$7738 ( \8081 , \8079 , \8080 );
and \U$7739 ( \8082 , \8081 , \6180 );
not \U$7740 ( \8083 , \8081 );
and \U$7741 ( \8084 , \8083 , \6190 );
nor \U$7742 ( \8085 , \8082 , \8084 );
and \U$7743 ( \8086 , \8078 , \8085 );
and \U$7744 ( \8087 , \8070 , \8077 );
or \U$7745 ( \8088 , \8086 , \8087 );
and \U$7746 ( \8089 , \8063 , \8088 );
and \U$7747 ( \8090 , \8039 , \8062 );
or \U$7748 ( \8091 , \8089 , \8090 );
and \U$7749 ( \8092 , \3254 , RI986e710_23);
and \U$7750 ( \8093 , RI986e620_21, \3252 );
nor \U$7751 ( \8094 , \8092 , \8093 );
not \U$7752 ( \8095 , \8094 );
not \U$7753 ( \8096 , \2935 );
and \U$7754 ( \8097 , \8095 , \8096 );
and \U$7755 ( \8098 , \8094 , \2935 );
nor \U$7756 ( \8099 , \8097 , \8098 );
and \U$7757 ( \8100 , \2274 , RI986f250_47);
and \U$7758 ( \8101 , RI986f160_45, \2272 );
nor \U$7759 ( \8102 , \8100 , \8101 );
and \U$7760 ( \8103 , \8102 , \2031 );
not \U$7761 ( \8104 , \8102 );
and \U$7762 ( \8105 , \8104 , \2030 );
nor \U$7763 ( \8106 , \8103 , \8105 );
xor \U$7764 ( \8107 , \8099 , \8106 );
and \U$7765 ( \8108 , \2464 , RI986e530_19);
and \U$7766 ( \8109 , RI986e440_17, \2462 );
nor \U$7767 ( \8110 , \8108 , \8109 );
and \U$7768 ( \8111 , \8110 , \2263 );
not \U$7769 ( \8112 , \8110 );
and \U$7770 ( \8113 , \8112 , \2468 );
nor \U$7771 ( \8114 , \8111 , \8113 );
and \U$7772 ( \8115 , \8107 , \8114 );
and \U$7773 ( \8116 , \8099 , \8106 );
or \U$7774 ( \8117 , \8115 , \8116 );
and \U$7775 ( \8118 , \2042 , RI986f070_43);
and \U$7776 ( \8119 , RI986ef80_41, \2040 );
nor \U$7777 ( \8120 , \8118 , \8119 );
not \U$7778 ( \8121 , \8120 );
not \U$7779 ( \8122 , \1462 );
and \U$7780 ( \8123 , \8121 , \8122 );
and \U$7781 ( \8124 , \8120 , \2034 );
nor \U$7782 ( \8125 , \8123 , \8124 );
and \U$7783 ( \8126 , \1329 , RI986ee90_39);
and \U$7784 ( \8127 , RI986eda0_37, \1327 );
nor \U$7785 ( \8128 , \8126 , \8127 );
and \U$7786 ( \8129 , \8128 , \1337 );
not \U$7787 ( \8130 , \8128 );
and \U$7788 ( \8131 , \8130 , \1336 );
nor \U$7789 ( \8132 , \8129 , \8131 );
xor \U$7790 ( \8133 , \8125 , \8132 );
and \U$7791 ( \8134 , \1311 , RI986ebc0_33);
and \U$7792 ( \8135 , RI986ecb0_35, \1309 );
nor \U$7793 ( \8136 , \8134 , \8135 );
and \U$7794 ( \8137 , \8136 , \1318 );
not \U$7795 ( \8138 , \8136 );
and \U$7796 ( \8139 , \8138 , \1458 );
nor \U$7797 ( \8140 , \8137 , \8139 );
and \U$7798 ( \8141 , \8133 , \8140 );
and \U$7799 ( \8142 , \8125 , \8132 );
or \U$7800 ( \8143 , \8141 , \8142 );
xor \U$7801 ( \8144 , \8117 , \8143 );
and \U$7802 ( \8145 , \438 , RI9871500_121);
and \U$7803 ( \8146 , RI98715f0_123, \436 );
nor \U$7804 ( \8147 , \8145 , \8146 );
and \U$7805 ( \8148 , \8147 , \443 );
not \U$7806 ( \8149 , \8147 );
and \U$7807 ( \8150 , \8149 , \444 );
nor \U$7808 ( \8151 , \8148 , \8150 );
and \U$7809 ( \8152 , \776 , RI986ead0_31);
and \U$7810 ( \8153 , RI986e9e0_29, \774 );
nor \U$7811 ( \8154 , \8152 , \8153 );
and \U$7812 ( \8155 , \8154 , \451 );
not \U$7813 ( \8156 , \8154 );
and \U$7814 ( \8157 , \8156 , \474 );
nor \U$7815 ( \8158 , \8155 , \8157 );
xor \U$7816 ( \8159 , \8151 , \8158 );
and \U$7817 ( \8160 , \1293 , RI986e8f0_27);
and \U$7818 ( \8161 , RI986e800_25, \1291 );
nor \U$7819 ( \8162 , \8160 , \8161 );
not \U$7820 ( \8163 , \8162 );
not \U$7821 ( \8164 , \1128 );
and \U$7822 ( \8165 , \8163 , \8164 );
and \U$7823 ( \8166 , \8162 , \1301 );
nor \U$7824 ( \8167 , \8165 , \8166 );
and \U$7825 ( \8168 , \8159 , \8167 );
and \U$7826 ( \8169 , \8151 , \8158 );
or \U$7827 ( \8170 , \8168 , \8169 );
and \U$7828 ( \8171 , \8144 , \8170 );
and \U$7829 ( \8172 , \8117 , \8143 );
or \U$7830 ( \8173 , \8171 , \8172 );
or \U$7831 ( \8174 , \8091 , \8173 );
not \U$7832 ( \8175 , \8091 );
not \U$7833 ( \8176 , \8173 );
or \U$7834 ( \8177 , \8175 , \8176 );
and \U$7835 ( \8178 , \395 , RI9871230_115);
and \U$7836 ( \8179 , RI9871140_113, \393 );
nor \U$7837 ( \8180 , \8178 , \8179 );
not \U$7838 ( \8181 , \8180 );
not \U$7839 ( \8182 , \386 );
and \U$7840 ( \8183 , \8181 , \8182 );
and \U$7841 ( \8184 , \8180 , \487 );
nor \U$7842 ( \8185 , \8183 , \8184 );
and \U$7843 ( \8186 , \465 , RI98716e0_125);
and \U$7844 ( \8187 , RI98717d0_127, \463 );
nor \U$7845 ( \8188 , \8186 , \8187 );
not \U$7846 ( \8189 , \8188 );
not \U$7847 ( \8190 , \454 );
and \U$7848 ( \8191 , \8189 , \8190 );
and \U$7849 ( \8192 , \8188 , \456 );
nor \U$7850 ( \8193 , \8191 , \8192 );
xor \U$7851 ( \8194 , \8185 , \8193 );
and \U$7852 ( \8195 , \376 , RI9871320_117);
and \U$7853 ( \8196 , RI9871410_119, \374 );
nor \U$7854 ( \8197 , \8195 , \8196 );
not \U$7855 ( \8198 , \8197 );
not \U$7856 ( \8199 , \365 );
and \U$7857 ( \8200 , \8198 , \8199 );
and \U$7858 ( \8201 , \8197 , \367 );
nor \U$7859 ( \8202 , \8200 , \8201 );
and \U$7860 ( \8203 , \8194 , \8202 );
and \U$7861 ( \8204 , \8185 , \8193 );
or \U$7862 ( \8205 , \8203 , \8204 );
and \U$7863 ( \8206 , \416 , RI9870e70_107);
and \U$7864 ( \8207 , RI9870ba0_101, \414 );
nor \U$7865 ( \8208 , \8206 , \8207 );
and \U$7866 ( \8209 , \8208 , \421 );
not \U$7867 ( \8210 , \8208 );
and \U$7868 ( \8211 , \8210 , \422 );
nor \U$7869 ( \8212 , \8209 , \8211 );
nand \U$7870 ( \8213 , RI98709c0_97, RI9871fc8_144);
xor \U$7871 ( \8214 , \8212 , \8213 );
and \U$7872 ( \8215 , \354 , RI9871050_111);
and \U$7873 ( \8216 , RI9870c90_103, \352 );
nor \U$7874 ( \8217 , \8215 , \8216 );
not \U$7875 ( \8218 , \8217 );
not \U$7876 ( \8219 , \345 );
and \U$7877 ( \8220 , \8218 , \8219 );
and \U$7878 ( \8221 , \8217 , \361 );
nor \U$7879 ( \8222 , \8220 , \8221 );
and \U$7880 ( \8223 , \8214 , \8222 );
and \U$7881 ( \8224 , \8212 , \8213 );
or \U$7882 ( \8225 , \8223 , \8224 );
or \U$7883 ( \8226 , \8205 , \8225 );
not \U$7884 ( \8227 , \8225 );
not \U$7885 ( \8228 , \8205 );
or \U$7886 ( \8229 , \8227 , \8228 );
or \U$7887 ( \8230 , \7775 , \7768 );
nand \U$7888 ( \8231 , \8230 , \7776 );
nand \U$7889 ( \8232 , \8229 , \8231 );
nand \U$7890 ( \8233 , \8226 , \8232 );
nand \U$7891 ( \8234 , \8177 , \8233 );
nand \U$7892 ( \8235 , \8174 , \8234 );
xor \U$7893 ( \8236 , \8012 , \8235 );
xor \U$7894 ( \8237 , \7476 , \7480 );
xor \U$7895 ( \8238 , \8237 , \7488 );
xor \U$7896 ( \8239 , \7660 , \7662 );
xor \U$7897 ( \8240 , \8239 , \7665 );
and \U$7898 ( \8241 , \8238 , \8240 );
xor \U$7899 ( \8242 , \7420 , \7428 );
xor \U$7900 ( \8243 , \8242 , \7436 );
xor \U$7901 ( \8244 , \7648 , \7653 );
xor \U$7902 ( \8245 , \8243 , \8244 );
xor \U$7903 ( \8246 , \7660 , \7662 );
xor \U$7904 ( \8247 , \8246 , \7665 );
and \U$7905 ( \8248 , \8245 , \8247 );
and \U$7906 ( \8249 , \8238 , \8245 );
or \U$7907 ( \8250 , \8241 , \8248 , \8249 );
and \U$7908 ( \8251 , \8236 , \8250 );
and \U$7909 ( \8252 , \8012 , \8235 );
or \U$7910 ( \8253 , \8251 , \8252 );
xor \U$7911 ( \8254 , \7342 , \7344 );
xor \U$7912 ( \8255 , \8254 , \7357 );
xor \U$7913 ( \8256 , \8253 , \8255 );
xor \U$7914 ( \8257 , \7776 , \7783 );
xor \U$7915 ( \8258 , \8257 , \7812 );
xor \U$7916 ( \8259 , \7703 , \7737 );
xor \U$7917 ( \8260 , \8259 , \7764 );
and \U$7918 ( \8261 , \8258 , \8260 );
xor \U$7919 ( \8262 , \7842 , \7870 );
xor \U$7920 ( \8263 , \8262 , \7899 );
xor \U$7921 ( \8264 , \7703 , \7737 );
xor \U$7922 ( \8265 , \8264 , \7764 );
and \U$7923 ( \8266 , \8263 , \8265 );
and \U$7924 ( \8267 , \8258 , \8263 );
or \U$7925 ( \8268 , \8261 , \8266 , \8267 );
xor \U$7926 ( \8269 , \7469 , \7491 );
xor \U$7927 ( \8270 , \8269 , \7518 );
xor \U$7928 ( \8271 , \8268 , \8270 );
xor \U$7929 ( \8272 , \7550 , \7003 );
xor \U$7930 ( \8273 , \8272 , \7557 );
xor \U$7931 ( \8274 , \7908 , \7915 );
xor \U$7932 ( \8275 , \8273 , \8274 );
and \U$7933 ( \8276 , \8271 , \8275 );
and \U$7934 ( \8277 , \8268 , \8270 );
or \U$7935 ( \8278 , \8276 , \8277 );
and \U$7936 ( \8279 , \8256 , \8278 );
and \U$7937 ( \8280 , \8253 , \8255 );
or \U$7938 ( \8281 , \8279 , \8280 );
xor \U$7939 ( \8282 , \6968 , \6994 );
xor \U$7940 ( \8283 , \8282 , \6999 );
xor \U$7941 ( \8284 , \7312 , \7319 );
xor \U$7942 ( \8285 , \8283 , \8284 );
xor \U$7943 ( \8286 , \8281 , \8285 );
xor \U$7944 ( \8287 , \7931 , \7933 );
not \U$7945 ( \8288 , \8287 );
not \U$7946 ( \8289 , \7939 );
or \U$7947 ( \8290 , \8288 , \8289 );
or \U$7948 ( \8291 , \7939 , \8287 );
nand \U$7949 ( \8292 , \8290 , \8291 );
xor \U$7950 ( \8293 , \7442 , \7521 );
xor \U$7951 ( \8294 , \8293 , \7560 );
xor \U$7952 ( \8295 , \8292 , \8294 );
xor \U$7953 ( \8296 , \7676 , \7905 );
xor \U$7954 ( \8297 , \8296 , \7920 );
and \U$7955 ( \8298 , \8295 , \8297 );
and \U$7956 ( \8299 , \8292 , \8294 );
or \U$7957 ( \8300 , \8298 , \8299 );
and \U$7958 ( \8301 , \8286 , \8300 );
and \U$7959 ( \8302 , \8281 , \8285 );
or \U$7960 ( \8303 , \8301 , \8302 );
not \U$7961 ( \8304 , \7585 );
xor \U$7962 ( \8305 , \7563 , \7360 );
not \U$7963 ( \8306 , \8305 );
or \U$7964 ( \8307 , \8304 , \8306 );
or \U$7965 ( \8308 , \8305 , \7585 );
nand \U$7966 ( \8309 , \8307 , \8308 );
not \U$7967 ( \8310 , \7926 );
xor \U$7968 ( \8311 , \7941 , \7923 );
not \U$7969 ( \8312 , \8311 );
or \U$7970 ( \8313 , \8310 , \8312 );
or \U$7971 ( \8314 , \8311 , \7926 );
nand \U$7972 ( \8315 , \8313 , \8314 );
and \U$7973 ( \8316 , \8309 , \8315 );
xor \U$7974 ( \8317 , \8303 , \8316 );
not \U$7975 ( \8318 , \7636 );
not \U$7976 ( \8319 , \7642 );
not \U$7977 ( \8320 , \7943 );
and \U$7978 ( \8321 , \8319 , \8320 );
and \U$7979 ( \8322 , \7642 , \7943 );
nor \U$7980 ( \8323 , \8321 , \8322 );
not \U$7981 ( \8324 , \8323 );
or \U$7982 ( \8325 , \8318 , \8324 );
or \U$7983 ( \8326 , \8323 , \7636 );
nand \U$7984 ( \8327 , \8325 , \8326 );
and \U$7985 ( \8328 , \8317 , \8327 );
and \U$7986 ( \8329 , \8303 , \8316 );
or \U$7987 ( \8330 , \8328 , \8329 );
nand \U$7988 ( \8331 , \7966 , \8330 );
or \U$7989 ( \8332 , \7963 , \8331 );
xnor \U$7990 ( \8333 , \8331 , \7963 );
and \U$7991 ( \8334 , \2274 , RI986ef80_41);
and \U$7992 ( \8335 , RI986f250_47, \2272 );
nor \U$7993 ( \8336 , \8334 , \8335 );
and \U$7994 ( \8337 , \8336 , \2031 );
not \U$7995 ( \8338 , \8336 );
and \U$7996 ( \8339 , \8338 , \2030 );
nor \U$7997 ( \8340 , \8337 , \8339 );
not \U$7998 ( \8341 , \8340 );
and \U$7999 ( \8342 , \2464 , RI986f160_45);
and \U$8000 ( \8343 , RI986e530_19, \2462 );
nor \U$8001 ( \8344 , \8342 , \8343 );
and \U$8002 ( \8345 , \8344 , \2263 );
not \U$8003 ( \8346 , \8344 );
and \U$8004 ( \8347 , \8346 , \2468 );
nor \U$8005 ( \8348 , \8345 , \8347 );
not \U$8006 ( \8349 , \8348 );
and \U$8007 ( \8350 , \8341 , \8349 );
and \U$8008 ( \8351 , \8348 , \8340 );
and \U$8009 ( \8352 , \3254 , RI986e440_17);
and \U$8010 ( \8353 , RI986e710_23, \3252 );
nor \U$8011 ( \8354 , \8352 , \8353 );
not \U$8012 ( \8355 , \8354 );
not \U$8013 ( \8356 , \2935 );
and \U$8014 ( \8357 , \8355 , \8356 );
and \U$8015 ( \8358 , \8354 , \3406 );
nor \U$8016 ( \8359 , \8357 , \8358 );
nor \U$8017 ( \8360 , \8351 , \8359 );
nor \U$8018 ( \8361 , \8350 , \8360 );
and \U$8019 ( \8362 , \1311 , RI986eda0_37);
and \U$8020 ( \8363 , RI986ebc0_33, \1309 );
nor \U$8021 ( \8364 , \8362 , \8363 );
and \U$8022 ( \8365 , \8364 , \1315 );
not \U$8023 ( \8366 , \8364 );
and \U$8024 ( \8367 , \8366 , \1458 );
nor \U$8025 ( \8368 , \8365 , \8367 );
and \U$8026 ( \8369 , \1329 , RI986e800_25);
and \U$8027 ( \8370 , RI986ee90_39, \1327 );
nor \U$8028 ( \8371 , \8369 , \8370 );
and \U$8029 ( \8372 , \8371 , \1337 );
not \U$8030 ( \8373 , \8371 );
and \U$8031 ( \8374 , \8373 , \1336 );
nor \U$8032 ( \8375 , \8372 , \8374 );
xor \U$8033 ( \8376 , \8368 , \8375 );
and \U$8034 ( \8377 , \2042 , RI986ecb0_35);
and \U$8035 ( \8378 , RI986f070_43, \2040 );
nor \U$8036 ( \8379 , \8377 , \8378 );
not \U$8037 ( \8380 , \8379 );
not \U$8038 ( \8381 , \2034 );
and \U$8039 ( \8382 , \8380 , \8381 );
and \U$8040 ( \8383 , \8379 , \2034 );
nor \U$8041 ( \8384 , \8382 , \8383 );
and \U$8042 ( \8385 , \8376 , \8384 );
and \U$8043 ( \8386 , \8368 , \8375 );
or \U$8044 ( \8387 , \8385 , \8386 );
xor \U$8045 ( \8388 , \8361 , \8387 );
and \U$8046 ( \8389 , \776 , RI98715f0_123);
and \U$8047 ( \8390 , RI986ead0_31, \774 );
nor \U$8048 ( \8391 , \8389 , \8390 );
and \U$8049 ( \8392 , \8391 , \451 );
not \U$8050 ( \8393 , \8391 );
and \U$8051 ( \8394 , \8393 , \474 );
nor \U$8052 ( \8395 , \8392 , \8394 );
not \U$8053 ( \8396 , \8395 );
and \U$8054 ( \8397 , \438 , RI98717d0_127);
and \U$8055 ( \8398 , RI9871500_121, \436 );
nor \U$8056 ( \8399 , \8397 , \8398 );
and \U$8057 ( \8400 , \8399 , \443 );
not \U$8058 ( \8401 , \8399 );
and \U$8059 ( \8402 , \8401 , \444 );
nor \U$8060 ( \8403 , \8400 , \8402 );
not \U$8061 ( \8404 , \8403 );
and \U$8062 ( \8405 , \8396 , \8404 );
and \U$8063 ( \8406 , \8403 , \8395 );
and \U$8064 ( \8407 , \1293 , RI986e9e0_29);
and \U$8065 ( \8408 , RI986e8f0_27, \1291 );
nor \U$8066 ( \8409 , \8407 , \8408 );
not \U$8067 ( \8410 , \8409 );
not \U$8068 ( \8411 , \1128 );
and \U$8069 ( \8412 , \8410 , \8411 );
and \U$8070 ( \8413 , \8409 , \1128 );
nor \U$8071 ( \8414 , \8412 , \8413 );
nor \U$8072 ( \8415 , \8406 , \8414 );
nor \U$8073 ( \8416 , \8405 , \8415 );
and \U$8074 ( \8417 , \8388 , \8416 );
and \U$8075 ( \8418 , \8361 , \8387 );
or \U$8076 ( \8419 , \8417 , \8418 );
and \U$8077 ( \8420 , \5881 , RI986f610_55);
and \U$8078 ( \8421 , RI986df90_7, \5879 );
nor \U$8079 ( \8422 , \8420 , \8421 );
and \U$8080 ( \8423 , \8422 , \5594 );
not \U$8081 ( \8424 , \8422 );
and \U$8082 ( \8425 , \8424 , \5885 );
nor \U$8083 ( \8426 , \8423 , \8425 );
and \U$8084 ( \8427 , \6453 , RI986dea0_5);
and \U$8085 ( \8428 , RI986ddb0_3, \6451 );
nor \U$8086 ( \8429 , \8427 , \8428 );
and \U$8087 ( \8430 , \8429 , \6190 );
not \U$8088 ( \8431 , \8429 );
and \U$8089 ( \8432 , \8431 , \6705 );
nor \U$8090 ( \8433 , \8430 , \8432 );
xor \U$8091 ( \8434 , \8426 , \8433 );
and \U$8092 ( \8435 , \5318 , RI986f340_49);
and \U$8093 ( \8436 , RI986f520_53, \5316 );
nor \U$8094 ( \8437 , \8435 , \8436 );
and \U$8095 ( \8438 , \8437 , \5052 );
not \U$8096 ( \8439 , \8437 );
and \U$8097 ( \8440 , \8439 , \5322 );
nor \U$8098 ( \8441 , \8438 , \8440 );
and \U$8099 ( \8442 , \8434 , \8441 );
and \U$8100 ( \8443 , \8426 , \8433 );
nor \U$8101 ( \8444 , \8442 , \8443 );
and \U$8102 ( \8445 , \4710 , RI986f8e0_61);
and \U$8103 ( \8446 , RI986f430_51, \4708 );
nor \U$8104 ( \8447 , \8445 , \8446 );
not \U$8105 ( \8448 , \8447 );
not \U$8106 ( \8449 , \4521 );
and \U$8107 ( \8450 , \8448 , \8449 );
and \U$8108 ( \8451 , \8447 , \4519 );
nor \U$8109 ( \8452 , \8450 , \8451 );
and \U$8110 ( \8453 , \3683 , RI986e620_21);
and \U$8111 ( \8454 , RI986f7f0_59, \3681 );
nor \U$8112 ( \8455 , \8453 , \8454 );
not \U$8113 ( \8456 , \8455 );
not \U$8114 ( \8457 , \3918 );
and \U$8115 ( \8458 , \8456 , \8457 );
and \U$8116 ( \8459 , \8455 , \3918 );
nor \U$8117 ( \8460 , \8458 , \8459 );
xor \U$8118 ( \8461 , \8452 , \8460 );
and \U$8119 ( \8462 , \4203 , RI986f700_57);
and \U$8120 ( \8463 , RI986f9d0_63, \4201 );
nor \U$8121 ( \8464 , \8462 , \8463 );
and \U$8122 ( \8465 , \8464 , \3923 );
not \U$8123 ( \8466 , \8464 );
and \U$8124 ( \8467 , \8466 , \4207 );
nor \U$8125 ( \8468 , \8465 , \8467 );
and \U$8126 ( \8469 , \8461 , \8468 );
and \U$8127 ( \8470 , \8452 , \8460 );
or \U$8128 ( \8471 , \8469 , \8470 );
xor \U$8129 ( \8472 , \8444 , \8471 );
and \U$8130 ( \8473 , \7079 , RI986dcc0_1);
and \U$8131 ( \8474 , RI986e170_11, \7077 );
nor \U$8132 ( \8475 , \8473 , \8474 );
and \U$8133 ( \8476 , \8475 , \6709 );
not \U$8134 ( \8477 , \8475 );
and \U$8135 ( \8478 , \8477 , \6710 );
nor \U$8136 ( \8479 , \8476 , \8478 );
and \U$8137 ( \8480 , RI9872d60_173, RI9872dd8_174);
not \U$8138 ( \8481 , RI9872e50_175);
and \U$8139 ( \8482 , \8481 , RI9872dd8_174);
nor \U$8140 ( \8483 , \8481 , RI9872dd8_174);
or \U$8141 ( \8484 , \8482 , \8483 );
nor \U$8142 ( \8485 , RI9872d60_173, RI9872dd8_174);
nor \U$8143 ( \8486 , \8480 , \8484 , \8485 );
nand \U$8144 ( \8487 , RI986e350_15, \8486 );
and \U$8145 ( \8488 , \8487 , \8051 );
not \U$8146 ( \8489 , \8487 );
and \U$8147 ( \8490 , \8489 , \8050 );
nor \U$8148 ( \8491 , \8488 , \8490 );
xor \U$8149 ( \8492 , \8479 , \8491 );
and \U$8150 ( \8493 , \7729 , RI986e080_9);
and \U$8151 ( \8494 , RI986e260_13, \7727 );
nor \U$8152 ( \8495 , \8493 , \8494 );
and \U$8153 ( \8496 , \8495 , \7733 );
not \U$8154 ( \8497 , \8495 );
and \U$8155 ( \8498 , \8497 , \7480 );
nor \U$8156 ( \8499 , \8496 , \8498 );
and \U$8157 ( \8500 , \8492 , \8499 );
and \U$8158 ( \8501 , \8479 , \8491 );
or \U$8159 ( \8502 , \8500 , \8501 );
and \U$8160 ( \8503 , \8472 , \8502 );
and \U$8161 ( \8504 , \8444 , \8471 );
or \U$8162 ( \8505 , \8503 , \8504 );
xor \U$8163 ( \8506 , \8419 , \8505 );
and \U$8164 ( \8507 , \376 , RI9871140_113);
and \U$8165 ( \8508 , RI9871320_117, \374 );
nor \U$8166 ( \8509 , \8507 , \8508 );
not \U$8167 ( \8510 , \8509 );
not \U$8168 ( \8511 , \367 );
and \U$8169 ( \8512 , \8510 , \8511 );
and \U$8170 ( \8513 , \8509 , \365 );
nor \U$8171 ( \8514 , \8512 , \8513 );
not \U$8172 ( \8515 , \8514 );
and \U$8173 ( \8516 , \395 , RI9870c90_103);
and \U$8174 ( \8517 , RI9871230_115, \393 );
nor \U$8175 ( \8518 , \8516 , \8517 );
not \U$8176 ( \8519 , \8518 );
not \U$8177 ( \8520 , \386 );
and \U$8178 ( \8521 , \8519 , \8520 );
and \U$8179 ( \8522 , \8518 , \487 );
nor \U$8180 ( \8523 , \8521 , \8522 );
not \U$8181 ( \8524 , \8523 );
and \U$8182 ( \8525 , \8515 , \8524 );
and \U$8183 ( \8526 , \8523 , \8514 );
and \U$8184 ( \8527 , \465 , RI9871410_119);
and \U$8185 ( \8528 , RI98716e0_125, \463 );
nor \U$8186 ( \8529 , \8527 , \8528 );
not \U$8187 ( \8530 , \8529 );
not \U$8188 ( \8531 , \454 );
and \U$8189 ( \8532 , \8530 , \8531 );
and \U$8190 ( \8533 , \8529 , \456 );
nor \U$8191 ( \8534 , \8532 , \8533 );
nor \U$8192 ( \8535 , \8526 , \8534 );
nor \U$8193 ( \8536 , \8525 , \8535 );
and \U$8194 ( \8537 , \354 , RI9870ba0_101);
and \U$8195 ( \8538 , RI9871050_111, \352 );
nor \U$8196 ( \8539 , \8537 , \8538 );
not \U$8197 ( \8540 , \8539 );
not \U$8198 ( \8541 , \361 );
and \U$8199 ( \8542 , \8540 , \8541 );
and \U$8200 ( \8543 , \8539 , \361 );
nor \U$8201 ( \8544 , \8542 , \8543 );
nand \U$8202 ( \8545 , RI9870d80_105, RI9871fc8_144);
xor \U$8203 ( \8546 , \8544 , \8545 );
and \U$8204 ( \8547 , \416 , RI98709c0_97);
and \U$8205 ( \8548 , RI9870e70_107, \414 );
nor \U$8206 ( \8549 , \8547 , \8548 );
and \U$8207 ( \8550 , \8549 , \421 );
not \U$8208 ( \8551 , \8549 );
and \U$8209 ( \8552 , \8551 , \422 );
nor \U$8210 ( \8553 , \8550 , \8552 );
and \U$8211 ( \8554 , \8546 , \8553 );
and \U$8212 ( \8555 , \8544 , \8545 );
or \U$8213 ( \8556 , \8554 , \8555 );
xor \U$8214 ( \8557 , \8536 , \8556 );
xor \U$8215 ( \8558 , \8212 , \8213 );
xor \U$8216 ( \8559 , \8558 , \8222 );
and \U$8217 ( \8560 , \8557 , \8559 );
and \U$8218 ( \8561 , \8536 , \8556 );
or \U$8219 ( \8562 , \8560 , \8561 );
xor \U$8220 ( \8563 , \8506 , \8562 );
xor \U$8221 ( \8564 , \8125 , \8132 );
xor \U$8222 ( \8565 , \8564 , \8140 );
xor \U$8223 ( \8566 , \8185 , \8193 );
xor \U$8224 ( \8567 , \8566 , \8202 );
xor \U$8225 ( \8568 , \8565 , \8567 );
xor \U$8226 ( \8569 , \8151 , \8158 );
xor \U$8227 ( \8570 , \8569 , \8167 );
and \U$8228 ( \8571 , \8568 , \8570 );
and \U$8229 ( \8572 , \8565 , \8567 );
or \U$8230 ( \8573 , \8571 , \8572 );
not \U$8231 ( \8574 , \7735 );
not \U$8232 ( \8575 , \7717 );
or \U$8233 ( \8576 , \8574 , \8575 );
or \U$8234 ( \8577 , \7717 , \7735 );
nand \U$8235 ( \8578 , \8576 , \8577 );
not \U$8236 ( \8579 , \8578 );
not \U$8237 ( \8580 , \7710 );
and \U$8238 ( \8581 , \8579 , \8580 );
and \U$8239 ( \8582 , \8578 , \7710 );
nor \U$8240 ( \8583 , \8581 , \8582 );
xor \U$8241 ( \8584 , \8573 , \8583 );
xor \U$8242 ( \8585 , \8099 , \8106 );
xor \U$8243 ( \8586 , \8585 , \8114 );
xor \U$8244 ( \8587 , \8070 , \8077 );
xor \U$8245 ( \8588 , \8587 , \8085 );
and \U$8246 ( \8589 , \8586 , \8588 );
xor \U$8247 ( \8590 , \8020 , \8027 );
xor \U$8248 ( \8591 , \8590 , \8036 );
xor \U$8249 ( \8592 , \8070 , \8077 );
xor \U$8250 ( \8593 , \8592 , \8085 );
and \U$8251 ( \8594 , \8591 , \8593 );
and \U$8252 ( \8595 , \8586 , \8591 );
or \U$8253 ( \8596 , \8589 , \8594 , \8595 );
xor \U$8254 ( \8597 , \8584 , \8596 );
and \U$8255 ( \8598 , \8563 , \8597 );
not \U$8256 ( \8599 , \8007 );
not \U$8257 ( \8600 , \8001 );
or \U$8258 ( \8601 , \8599 , \8600 );
or \U$8259 ( \8602 , \8001 , \8007 );
nand \U$8260 ( \8603 , \8601 , \8602 );
not \U$8261 ( \8604 , \8603 );
not \U$8262 ( \8605 , \7991 );
and \U$8263 ( \8606 , \8604 , \8605 );
and \U$8264 ( \8607 , \8603 , \7991 );
nor \U$8265 ( \8608 , \8606 , \8607 );
not \U$8266 ( \8609 , \8608 );
xor \U$8267 ( \8610 , \7823 , \7831 );
xor \U$8268 ( \8611 , \8610 , \7839 );
xor \U$8269 ( \8612 , \7968 , \7973 );
xor \U$8270 ( \8613 , \8611 , \8612 );
not \U$8271 ( \8614 , \8613 );
or \U$8272 ( \8615 , \8609 , \8614 );
or \U$8273 ( \8616 , \8608 , \8613 );
nand \U$8274 ( \8617 , \8615 , \8616 );
not \U$8275 ( \8618 , \8617 );
xnor \U$8276 ( \8619 , \8225 , \8205 );
not \U$8277 ( \8620 , \8619 );
not \U$8278 ( \8621 , \8231 );
and \U$8279 ( \8622 , \8620 , \8621 );
and \U$8280 ( \8623 , \8619 , \8231 );
nor \U$8281 ( \8624 , \8622 , \8623 );
not \U$8282 ( \8625 , \8624 );
and \U$8283 ( \8626 , \8618 , \8625 );
and \U$8284 ( \8627 , \8617 , \8624 );
nor \U$8285 ( \8628 , \8626 , \8627 );
xor \U$8286 ( \8629 , \8573 , \8583 );
xor \U$8287 ( \8630 , \8629 , \8596 );
and \U$8288 ( \8631 , \8628 , \8630 );
and \U$8289 ( \8632 , \8563 , \8628 );
or \U$8290 ( \8633 , \8598 , \8631 , \8632 );
xor \U$8291 ( \8634 , \8117 , \8143 );
xor \U$8292 ( \8635 , \8634 , \8170 );
xor \U$8293 ( \8636 , \8039 , \8062 );
xor \U$8294 ( \8637 , \8636 , \8088 );
xor \U$8295 ( \8638 , \8635 , \8637 );
xor \U$8296 ( \8639 , \8444 , \8471 );
xor \U$8297 ( \8640 , \8639 , \8502 );
xor \U$8298 ( \8641 , \8536 , \8556 );
xor \U$8299 ( \8642 , \8641 , \8559 );
xor \U$8300 ( \8643 , \8640 , \8642 );
xor \U$8301 ( \8644 , \8361 , \8387 );
xor \U$8302 ( \8645 , \8644 , \8416 );
and \U$8303 ( \8646 , \8643 , \8645 );
and \U$8304 ( \8647 , \8640 , \8642 );
or \U$8305 ( \8648 , \8646 , \8647 );
and \U$8306 ( \8649 , \8638 , \8648 );
and \U$8307 ( \8650 , \8635 , \8637 );
or \U$8308 ( \8651 , \8649 , \8650 );
or \U$8309 ( \8652 , \8633 , \8651 );
not \U$8310 ( \8653 , \8651 );
not \U$8311 ( \8654 , \8633 );
or \U$8312 ( \8655 , \8653 , \8654 );
and \U$8313 ( \8656 , \1311 , RI986ee90_39);
and \U$8314 ( \8657 , RI986eda0_37, \1309 );
nor \U$8315 ( \8658 , \8656 , \8657 );
and \U$8316 ( \8659 , \8658 , \1315 );
not \U$8317 ( \8660 , \8658 );
and \U$8318 ( \8661 , \8660 , \1458 );
nor \U$8319 ( \8662 , \8659 , \8661 );
not \U$8320 ( \8663 , \8662 );
and \U$8321 ( \8664 , \2042 , RI986ebc0_33);
and \U$8322 ( \8665 , RI986ecb0_35, \2040 );
nor \U$8323 ( \8666 , \8664 , \8665 );
not \U$8324 ( \8667 , \8666 );
not \U$8325 ( \8668 , \2034 );
and \U$8326 ( \8669 , \8667 , \8668 );
and \U$8327 ( \8670 , \8666 , \2034 );
nor \U$8328 ( \8671 , \8669 , \8670 );
not \U$8329 ( \8672 , \8671 );
and \U$8330 ( \8673 , \8663 , \8672 );
and \U$8331 ( \8674 , \8671 , \8662 );
and \U$8332 ( \8675 , \2274 , RI986f070_43);
and \U$8333 ( \8676 , RI986ef80_41, \2272 );
nor \U$8334 ( \8677 , \8675 , \8676 );
and \U$8335 ( \8678 , \8677 , \2031 );
not \U$8336 ( \8679 , \8677 );
and \U$8337 ( \8680 , \8679 , \2030 );
nor \U$8338 ( \8681 , \8678 , \8680 );
nor \U$8339 ( \8682 , \8674 , \8681 );
nor \U$8340 ( \8683 , \8673 , \8682 );
and \U$8341 ( \8684 , \776 , RI9871500_121);
and \U$8342 ( \8685 , RI98715f0_123, \774 );
nor \U$8343 ( \8686 , \8684 , \8685 );
and \U$8344 ( \8687 , \8686 , \451 );
not \U$8345 ( \8688 , \8686 );
and \U$8346 ( \8689 , \8688 , \474 );
nor \U$8347 ( \8690 , \8687 , \8689 );
not \U$8348 ( \8691 , \8690 );
and \U$8349 ( \8692 , \1293 , RI986ead0_31);
and \U$8350 ( \8693 , RI986e9e0_29, \1291 );
nor \U$8351 ( \8694 , \8692 , \8693 );
not \U$8352 ( \8695 , \8694 );
not \U$8353 ( \8696 , \1128 );
and \U$8354 ( \8697 , \8695 , \8696 );
and \U$8355 ( \8698 , \8694 , \1128 );
nor \U$8356 ( \8699 , \8697 , \8698 );
not \U$8357 ( \8700 , \8699 );
and \U$8358 ( \8701 , \8691 , \8700 );
and \U$8359 ( \8702 , \8699 , \8690 );
and \U$8360 ( \8703 , \1329 , RI986e8f0_27);
and \U$8361 ( \8704 , RI986e800_25, \1327 );
nor \U$8362 ( \8705 , \8703 , \8704 );
and \U$8363 ( \8706 , \8705 , \1337 );
not \U$8364 ( \8707 , \8705 );
and \U$8365 ( \8708 , \8707 , \1336 );
nor \U$8366 ( \8709 , \8706 , \8708 );
nor \U$8367 ( \8710 , \8702 , \8709 );
nor \U$8368 ( \8711 , \8701 , \8710 );
xor \U$8369 ( \8712 , \8683 , \8711 );
not \U$8370 ( \8713 , \3406 );
and \U$8371 ( \8714 , \3254 , RI986e530_19);
and \U$8372 ( \8715 , RI986e440_17, \3252 );
nor \U$8373 ( \8716 , \8714 , \8715 );
not \U$8374 ( \8717 , \8716 );
or \U$8375 ( \8718 , \8713 , \8717 );
or \U$8376 ( \8719 , \8716 , \3406 );
nand \U$8377 ( \8720 , \8718 , \8719 );
not \U$8378 ( \8721 , \3412 );
and \U$8379 ( \8722 , \3683 , RI986e710_23);
and \U$8380 ( \8723 , RI986e620_21, \3681 );
nor \U$8381 ( \8724 , \8722 , \8723 );
not \U$8382 ( \8725 , \8724 );
or \U$8383 ( \8726 , \8721 , \8725 );
or \U$8384 ( \8727 , \8724 , \3412 );
nand \U$8385 ( \8728 , \8726 , \8727 );
xor \U$8386 ( \8729 , \8720 , \8728 );
and \U$8387 ( \8730 , \2464 , RI986f250_47);
and \U$8388 ( \8731 , RI986f160_45, \2462 );
nor \U$8389 ( \8732 , \8730 , \8731 );
and \U$8390 ( \8733 , \8732 , \2468 );
not \U$8391 ( \8734 , \8732 );
and \U$8392 ( \8735 , \8734 , \2263 );
nor \U$8393 ( \8736 , \8733 , \8735 );
and \U$8394 ( \8737 , \8729 , \8736 );
and \U$8395 ( \8738 , \8720 , \8728 );
nor \U$8396 ( \8739 , \8737 , \8738 );
and \U$8397 ( \8740 , \8712 , \8739 );
and \U$8398 ( \8741 , \8683 , \8711 );
or \U$8399 ( \8742 , \8740 , \8741 );
and \U$8400 ( \8743 , \465 , RI9871320_117);
and \U$8401 ( \8744 , RI9871410_119, \463 );
nor \U$8402 ( \8745 , \8743 , \8744 );
not \U$8403 ( \8746 , \8745 );
not \U$8404 ( \8747 , \454 );
and \U$8405 ( \8748 , \8746 , \8747 );
and \U$8406 ( \8749 , \8745 , \456 );
nor \U$8407 ( \8750 , \8748 , \8749 );
and \U$8408 ( \8751 , \376 , RI9871230_115);
and \U$8409 ( \8752 , RI9871140_113, \374 );
nor \U$8410 ( \8753 , \8751 , \8752 );
not \U$8411 ( \8754 , \8753 );
not \U$8412 ( \8755 , \367 );
and \U$8413 ( \8756 , \8754 , \8755 );
and \U$8414 ( \8757 , \8753 , \367 );
nor \U$8415 ( \8758 , \8756 , \8757 );
or \U$8416 ( \8759 , \8750 , \8758 );
not \U$8417 ( \8760 , \8758 );
not \U$8418 ( \8761 , \8750 );
or \U$8419 ( \8762 , \8760 , \8761 );
and \U$8420 ( \8763 , \438 , RI98716e0_125);
and \U$8421 ( \8764 , RI98717d0_127, \436 );
nor \U$8422 ( \8765 , \8763 , \8764 );
and \U$8423 ( \8766 , \8765 , \444 );
not \U$8424 ( \8767 , \8765 );
and \U$8425 ( \8768 , \8767 , \443 );
nor \U$8426 ( \8769 , \8766 , \8768 );
nand \U$8427 ( \8770 , \8762 , \8769 );
nand \U$8428 ( \8771 , \8759 , \8770 );
and \U$8429 ( \8772 , \395 , RI9871050_111);
and \U$8430 ( \8773 , RI9870c90_103, \393 );
nor \U$8431 ( \8774 , \8772 , \8773 );
not \U$8432 ( \8775 , \8774 );
not \U$8433 ( \8776 , \386 );
and \U$8434 ( \8777 , \8775 , \8776 );
and \U$8435 ( \8778 , \8774 , \386 );
nor \U$8436 ( \8779 , \8777 , \8778 );
and \U$8437 ( \8780 , \416 , RI9870d80_105);
and \U$8438 ( \8781 , RI98709c0_97, \414 );
nor \U$8439 ( \8782 , \8780 , \8781 );
and \U$8440 ( \8783 , \8782 , \421 );
not \U$8441 ( \8784 , \8782 );
and \U$8442 ( \8785 , \8784 , \422 );
nor \U$8443 ( \8786 , \8783 , \8785 );
or \U$8444 ( \8787 , \8779 , \8786 );
not \U$8445 ( \8788 , \8786 );
not \U$8446 ( \8789 , \8779 );
or \U$8447 ( \8790 , \8788 , \8789 );
not \U$8448 ( \8791 , \345 );
and \U$8449 ( \8792 , \354 , RI9870e70_107);
and \U$8450 ( \8793 , RI9870ba0_101, \352 );
nor \U$8451 ( \8794 , \8792 , \8793 );
not \U$8452 ( \8795 , \8794 );
or \U$8453 ( \8796 , \8791 , \8795 );
or \U$8454 ( \8797 , \8794 , \361 );
nand \U$8455 ( \8798 , \8796 , \8797 );
nand \U$8456 ( \8799 , \8790 , \8798 );
nand \U$8457 ( \8800 , \8787 , \8799 );
nor \U$8458 ( \8801 , \8771 , \8800 );
xor \U$8459 ( \8802 , \8742 , \8801 );
and \U$8460 ( \8803 , \7079 , RI986ddb0_3);
and \U$8461 ( \8804 , RI986dcc0_1, \7077 );
nor \U$8462 ( \8805 , \8803 , \8804 );
and \U$8463 ( \8806 , \8805 , \6709 );
not \U$8464 ( \8807 , \8805 );
and \U$8465 ( \8808 , \8807 , \6710 );
nor \U$8466 ( \8809 , \8806 , \8808 );
and \U$8467 ( \8810 , \5881 , RI986f520_53);
and \U$8468 ( \8811 , RI986f610_55, \5879 );
nor \U$8469 ( \8812 , \8810 , \8811 );
and \U$8470 ( \8813 , \8812 , \5885 );
not \U$8471 ( \8814 , \8812 );
and \U$8472 ( \8815 , \8814 , \5594 );
nor \U$8473 ( \8816 , \8813 , \8815 );
xor \U$8474 ( \8817 , \8809 , \8816 );
and \U$8475 ( \8818 , \6453 , RI986df90_7);
and \U$8476 ( \8819 , RI986dea0_5, \6451 );
nor \U$8477 ( \8820 , \8818 , \8819 );
and \U$8478 ( \8821 , \8820 , \6180 );
not \U$8479 ( \8822 , \8820 );
and \U$8480 ( \8823 , \8822 , \6190 );
nor \U$8481 ( \8824 , \8821 , \8823 );
and \U$8482 ( \8825 , \8817 , \8824 );
and \U$8483 ( \8826 , \8809 , \8816 );
or \U$8484 ( \8827 , \8825 , \8826 );
and \U$8485 ( \8828 , \8486 , RI986e260_13);
and \U$8486 ( \8829 , RI986e350_15, \8484 );
nor \U$8487 ( \8830 , \8828 , \8829 );
and \U$8488 ( \8831 , \8830 , \8051 );
not \U$8489 ( \8832 , \8830 );
and \U$8490 ( \8833 , \8832 , \8050 );
nor \U$8491 ( \8834 , \8831 , \8833 );
nand \U$8492 ( \8835 , RI9872f40_177, RI9872ec8_176);
and \U$8493 ( \8836 , \8835 , RI9872e50_175);
xor \U$8494 ( \8837 , \8834 , \8836 );
and \U$8495 ( \8838 , \7729 , RI986e170_11);
and \U$8496 ( \8839 , RI986e080_9, \7727 );
nor \U$8497 ( \8840 , \8838 , \8839 );
and \U$8498 ( \8841 , \8840 , \7733 );
not \U$8499 ( \8842 , \8840 );
and \U$8500 ( \8843 , \8842 , \7480 );
nor \U$8501 ( \8844 , \8841 , \8843 );
and \U$8502 ( \8845 , \8837 , \8844 );
and \U$8503 ( \8846 , \8834 , \8836 );
or \U$8504 ( \8847 , \8845 , \8846 );
xor \U$8505 ( \8848 , \8827 , \8847 );
and \U$8506 ( \8849 , \5318 , RI986f430_51);
and \U$8507 ( \8850 , RI986f340_49, \5316 );
nor \U$8508 ( \8851 , \8849 , \8850 );
and \U$8509 ( \8852 , \8851 , \5322 );
not \U$8510 ( \8853 , \8851 );
and \U$8511 ( \8854 , \8853 , \5052 );
nor \U$8512 ( \8855 , \8852 , \8854 );
and \U$8513 ( \8856 , \4203 , RI986f7f0_59);
and \U$8514 ( \8857 , RI986f700_57, \4201 );
nor \U$8515 ( \8858 , \8856 , \8857 );
and \U$8516 ( \8859 , \8858 , \3922 );
not \U$8517 ( \8860 , \8858 );
and \U$8518 ( \8861 , \8860 , \4207 );
nor \U$8519 ( \8862 , \8859 , \8861 );
xor \U$8520 ( \8863 , \8855 , \8862 );
and \U$8521 ( \8864 , \4710 , RI986f9d0_63);
and \U$8522 ( \8865 , RI986f8e0_61, \4708 );
nor \U$8523 ( \8866 , \8864 , \8865 );
not \U$8524 ( \8867 , \8866 );
not \U$8525 ( \8868 , \4521 );
and \U$8526 ( \8869 , \8867 , \8868 );
and \U$8527 ( \8870 , \8866 , \4521 );
nor \U$8528 ( \8871 , \8869 , \8870 );
and \U$8529 ( \8872 , \8863 , \8871 );
and \U$8530 ( \8873 , \8855 , \8862 );
or \U$8531 ( \8874 , \8872 , \8873 );
and \U$8532 ( \8875 , \8848 , \8874 );
and \U$8533 ( \8876 , \8827 , \8847 );
or \U$8534 ( \8877 , \8875 , \8876 );
and \U$8535 ( \8878 , \8802 , \8877 );
and \U$8536 ( \8879 , \8742 , \8801 );
or \U$8537 ( \8880 , \8878 , \8879 );
xor \U$8538 ( \8881 , \8368 , \8375 );
xor \U$8539 ( \8882 , \8881 , \8384 );
xor \U$8540 ( \8883 , \8452 , \8460 );
xor \U$8541 ( \8884 , \8883 , \8468 );
or \U$8542 ( \8885 , \8882 , \8884 );
not \U$8543 ( \8886 , \8884 );
not \U$8544 ( \8887 , \8882 );
or \U$8545 ( \8888 , \8886 , \8887 );
not \U$8546 ( \8889 , \8340 );
xor \U$8547 ( \8890 , \8348 , \8359 );
not \U$8548 ( \8891 , \8890 );
or \U$8549 ( \8892 , \8889 , \8891 );
or \U$8550 ( \8893 , \8890 , \8340 );
nand \U$8551 ( \8894 , \8892 , \8893 );
nand \U$8552 ( \8895 , \8888 , \8894 );
nand \U$8553 ( \8896 , \8885 , \8895 );
xor \U$8554 ( \8897 , \8479 , \8491 );
xor \U$8555 ( \8898 , \8897 , \8499 );
not \U$8556 ( \8899 , \8898 );
xor \U$8557 ( \8900 , \8426 , \8433 );
xor \U$8558 ( \8901 , \8900 , \8441 );
nand \U$8559 ( \8902 , \8899 , \8901 );
not \U$8560 ( \8903 , \8902 );
and \U$8561 ( \8904 , \8896 , \8903 );
not \U$8562 ( \8905 , \8896 );
not \U$8563 ( \8906 , \8903 );
and \U$8564 ( \8907 , \8905 , \8906 );
not \U$8565 ( \8908 , \8403 );
xor \U$8566 ( \8909 , \8395 , \8414 );
not \U$8567 ( \8910 , \8909 );
or \U$8568 ( \8911 , \8908 , \8910 );
or \U$8569 ( \8912 , \8909 , \8403 );
nand \U$8570 ( \8913 , \8911 , \8912 );
not \U$8571 ( \8914 , \8523 );
xor \U$8572 ( \8915 , \8534 , \8514 );
not \U$8573 ( \8916 , \8915 );
or \U$8574 ( \8917 , \8914 , \8916 );
or \U$8575 ( \8918 , \8915 , \8523 );
nand \U$8576 ( \8919 , \8917 , \8918 );
and \U$8577 ( \8920 , \8913 , \8919 );
not \U$8578 ( \8921 , \8919 );
not \U$8579 ( \8922 , \8913 );
and \U$8580 ( \8923 , \8921 , \8922 );
xor \U$8581 ( \8924 , \8544 , \8545 );
xor \U$8582 ( \8925 , \8924 , \8553 );
nor \U$8583 ( \8926 , \8923 , \8925 );
nor \U$8584 ( \8927 , \8920 , \8926 );
nor \U$8585 ( \8928 , \8907 , \8927 );
nor \U$8586 ( \8929 , \8904 , \8928 );
xor \U$8587 ( \8930 , \8880 , \8929 );
xor \U$8588 ( \8931 , \8046 , \8051 );
xor \U$8589 ( \8932 , \8931 , \8059 );
xor \U$8590 ( \8933 , \8565 , \8567 );
xor \U$8591 ( \8934 , \8933 , \8570 );
and \U$8592 ( \8935 , \8932 , \8934 );
xor \U$8593 ( \8936 , \8070 , \8077 );
xor \U$8594 ( \8937 , \8936 , \8085 );
xor \U$8595 ( \8938 , \8586 , \8591 );
xor \U$8596 ( \8939 , \8937 , \8938 );
xor \U$8597 ( \8940 , \8565 , \8567 );
xor \U$8598 ( \8941 , \8940 , \8570 );
and \U$8599 ( \8942 , \8939 , \8941 );
and \U$8600 ( \8943 , \8932 , \8939 );
or \U$8601 ( \8944 , \8935 , \8942 , \8943 );
and \U$8602 ( \8945 , \8930 , \8944 );
and \U$8603 ( \8946 , \8880 , \8929 );
nor \U$8604 ( \8947 , \8945 , \8946 );
nand \U$8605 ( \8948 , \8655 , \8947 );
nand \U$8606 ( \8949 , \8652 , \8948 );
xor \U$8607 ( \8950 , \8573 , \8583 );
and \U$8608 ( \8951 , \8950 , \8596 );
and \U$8609 ( \8952 , \8573 , \8583 );
or \U$8610 ( \8953 , \8951 , \8952 );
xor \U$8611 ( \8954 , \8419 , \8505 );
and \U$8612 ( \8955 , \8954 , \8562 );
and \U$8613 ( \8956 , \8419 , \8505 );
or \U$8614 ( \8957 , \8955 , \8956 );
xnor \U$8615 ( \8958 , \8953 , \8957 );
not \U$8616 ( \8959 , \8958 );
or \U$8617 ( \8960 , \8608 , \8624 );
not \U$8618 ( \8961 , \8624 );
not \U$8619 ( \8962 , \8608 );
or \U$8620 ( \8963 , \8961 , \8962 );
nand \U$8621 ( \8964 , \8963 , \8613 );
nand \U$8622 ( \8965 , \8960 , \8964 );
not \U$8623 ( \8966 , \8965 );
and \U$8624 ( \8967 , \8959 , \8966 );
and \U$8625 ( \8968 , \8958 , \8965 );
nor \U$8626 ( \8969 , \8967 , \8968 );
xnor \U$8627 ( \8970 , \8091 , \8173 );
not \U$8628 ( \8971 , \8970 );
not \U$8629 ( \8972 , \8233 );
and \U$8630 ( \8973 , \8971 , \8972 );
and \U$8631 ( \8974 , \8970 , \8233 );
nor \U$8632 ( \8975 , \8973 , \8974 );
or \U$8633 ( \8976 , \8969 , \8975 );
not \U$8634 ( \8977 , \8975 );
not \U$8635 ( \8978 , \8969 );
or \U$8636 ( \8979 , \8977 , \8978 );
xor \U$8637 ( \8980 , \7978 , \7980 );
xor \U$8638 ( \8981 , \8980 , \8009 );
xor \U$8639 ( \8982 , \7703 , \7737 );
xor \U$8640 ( \8983 , \8982 , \7764 );
xor \U$8641 ( \8984 , \8258 , \8263 );
xor \U$8642 ( \8985 , \8983 , \8984 );
xor \U$8643 ( \8986 , \7660 , \7662 );
xor \U$8644 ( \8987 , \8986 , \7665 );
xor \U$8645 ( \8988 , \8238 , \8245 );
xor \U$8646 ( \8989 , \8987 , \8988 );
xor \U$8647 ( \8990 , \8985 , \8989 );
xor \U$8648 ( \8991 , \8981 , \8990 );
nand \U$8649 ( \8992 , \8979 , \8991 );
nand \U$8650 ( \8993 , \8976 , \8992 );
xor \U$8651 ( \8994 , \8949 , \8993 );
xor \U$8652 ( \8995 , \8268 , \8270 );
xor \U$8653 ( \8996 , \8995 , \8275 );
xor \U$8654 ( \8997 , \7767 , \7815 );
xor \U$8655 ( \8998 , \8997 , \7902 );
xor \U$8656 ( \8999 , \8012 , \8235 );
xor \U$8657 ( \9000 , \8999 , \8250 );
xor \U$8658 ( \9001 , \8998 , \9000 );
xor \U$8659 ( \9002 , \8996 , \9001 );
and \U$8660 ( \9003 , \8994 , \9002 );
and \U$8661 ( \9004 , \8949 , \8993 );
or \U$8662 ( \9005 , \9003 , \9004 );
xor \U$8663 ( \9006 , \8253 , \8255 );
xor \U$8664 ( \9007 , \9006 , \8278 );
xor \U$8665 ( \9008 , \9005 , \9007 );
or \U$8666 ( \9009 , \8957 , \8953 );
not \U$8667 ( \9010 , \8953 );
not \U$8668 ( \9011 , \8957 );
or \U$8669 ( \9012 , \9010 , \9011 );
nand \U$8670 ( \9013 , \9012 , \8965 );
nand \U$8671 ( \9014 , \9009 , \9013 );
xor \U$8672 ( \9015 , \7658 , \7668 );
xor \U$8673 ( \9016 , \9015 , \7673 );
xor \U$8674 ( \9017 , \9014 , \9016 );
xor \U$8675 ( \9018 , \7978 , \7980 );
xor \U$8676 ( \9019 , \9018 , \8009 );
and \U$8677 ( \9020 , \8985 , \9019 );
xor \U$8678 ( \9021 , \7978 , \7980 );
xor \U$8679 ( \9022 , \9021 , \8009 );
and \U$8680 ( \9023 , \8989 , \9022 );
and \U$8681 ( \9024 , \8985 , \8989 );
or \U$8682 ( \9025 , \9020 , \9023 , \9024 );
and \U$8683 ( \9026 , \9017 , \9025 );
and \U$8684 ( \9027 , \9014 , \9016 );
or \U$8685 ( \9028 , \9026 , \9027 );
xor \U$8686 ( \9029 , \8268 , \8270 );
xor \U$8687 ( \9030 , \9029 , \8275 );
and \U$8688 ( \9031 , \8998 , \9030 );
xor \U$8689 ( \9032 , \8268 , \8270 );
xor \U$8690 ( \9033 , \9032 , \8275 );
and \U$8691 ( \9034 , \9000 , \9033 );
and \U$8692 ( \9035 , \8998 , \9000 );
or \U$8693 ( \9036 , \9031 , \9034 , \9035 );
xor \U$8694 ( \9037 , \9028 , \9036 );
xor \U$8695 ( \9038 , \8292 , \8294 );
xor \U$8696 ( \9039 , \9038 , \8297 );
xor \U$8697 ( \9040 , \9037 , \9039 );
and \U$8698 ( \9041 , \9008 , \9040 );
and \U$8699 ( \9042 , \9005 , \9007 );
or \U$8700 ( \9043 , \9041 , \9042 );
xor \U$8701 ( \9044 , \9028 , \9036 );
and \U$8702 ( \9045 , \9044 , \9039 );
and \U$8703 ( \9046 , \9028 , \9036 );
or \U$8704 ( \9047 , \9045 , \9046 );
xor \U$8705 ( \9048 , \8309 , \8315 );
xor \U$8706 ( \9049 , \9047 , \9048 );
xor \U$8707 ( \9050 , \8281 , \8285 );
xor \U$8708 ( \9051 , \9050 , \8300 );
xor \U$8709 ( \9052 , \9049 , \9051 );
and \U$8710 ( \9053 , \9043 , \9052 );
not \U$8711 ( \9054 , \9053 );
xor \U$8712 ( \9055 , \9047 , \9048 );
and \U$8713 ( \9056 , \9055 , \9051 );
and \U$8714 ( \9057 , \9047 , \9048 );
or \U$8715 ( \9058 , \9056 , \9057 );
xor \U$8716 ( \9059 , \8303 , \8316 );
xor \U$8717 ( \9060 , \9059 , \8327 );
xor \U$8718 ( \9061 , \9058 , \9060 );
not \U$8719 ( \9062 , \9061 );
or \U$8720 ( \9063 , \9054 , \9062 );
xor \U$8721 ( \9064 , \9043 , \9052 );
xor \U$8722 ( \9065 , \9005 , \9007 );
xor \U$8723 ( \9066 , \9065 , \9040 );
not \U$8724 ( \9067 , \9066 );
xor \U$8725 ( \9068 , \8949 , \8993 );
xor \U$8726 ( \9069 , \9068 , \9002 );
xor \U$8727 ( \9070 , \9014 , \9016 );
xor \U$8728 ( \9071 , \9070 , \9025 );
and \U$8729 ( \9072 , \9069 , \9071 );
not \U$8730 ( \9073 , \9069 );
not \U$8731 ( \9074 , \9071 );
and \U$8732 ( \9075 , \9073 , \9074 );
xor \U$8733 ( \9076 , \8880 , \8929 );
xor \U$8734 ( \9077 , \9076 , \8944 );
xor \U$8735 ( \9078 , \8635 , \8637 );
xor \U$8736 ( \9079 , \9078 , \8648 );
and \U$8737 ( \9080 , \9077 , \9079 );
xor \U$8738 ( \9081 , \8573 , \8583 );
xor \U$8739 ( \9082 , \9081 , \8596 );
xor \U$8740 ( \9083 , \8563 , \8628 );
xor \U$8741 ( \9084 , \9082 , \9083 );
xor \U$8742 ( \9085 , \8635 , \8637 );
xor \U$8743 ( \9086 , \9085 , \8648 );
and \U$8744 ( \9087 , \9084 , \9086 );
and \U$8745 ( \9088 , \9077 , \9084 );
or \U$8746 ( \9089 , \9080 , \9087 , \9088 );
xor \U$8747 ( \9090 , \8834 , \8836 );
xor \U$8748 ( \9091 , \9090 , \8844 );
not \U$8749 ( \9092 , \9091 );
xor \U$8750 ( \9093 , \8855 , \8862 );
xor \U$8751 ( \9094 , \9093 , \8871 );
not \U$8752 ( \9095 , \9094 );
and \U$8753 ( \9096 , \9092 , \9095 );
and \U$8754 ( \9097 , \9091 , \9094 );
xor \U$8755 ( \9098 , \8809 , \8816 );
xor \U$8756 ( \9099 , \9098 , \8824 );
nor \U$8757 ( \9100 , \9097 , \9099 );
nor \U$8758 ( \9101 , \9096 , \9100 );
not \U$8759 ( \9102 , \9101 );
not \U$8760 ( \9103 , \8798 );
not \U$8761 ( \9104 , \8779 );
or \U$8762 ( \9105 , \9103 , \9104 );
or \U$8763 ( \9106 , \8779 , \8798 );
nand \U$8764 ( \9107 , \9105 , \9106 );
not \U$8765 ( \9108 , \9107 );
not \U$8766 ( \9109 , \8786 );
and \U$8767 ( \9110 , \9108 , \9109 );
and \U$8768 ( \9111 , \9107 , \8786 );
nor \U$8769 ( \9112 , \9110 , \9111 );
not \U$8770 ( \9113 , \9112 );
nand \U$8771 ( \9114 , RI9870ab0_99, RI9871fc8_144);
not \U$8772 ( \9115 , \9114 );
and \U$8773 ( \9116 , \9113 , \9115 );
and \U$8774 ( \9117 , \9112 , \9114 );
not \U$8775 ( \9118 , \8750 );
not \U$8776 ( \9119 , \8769 );
or \U$8777 ( \9120 , \9118 , \9119 );
or \U$8778 ( \9121 , \8750 , \8769 );
nand \U$8779 ( \9122 , \9120 , \9121 );
not \U$8780 ( \9123 , \9122 );
not \U$8781 ( \9124 , \8758 );
and \U$8782 ( \9125 , \9123 , \9124 );
and \U$8783 ( \9126 , \9122 , \8758 );
nor \U$8784 ( \9127 , \9125 , \9126 );
nor \U$8785 ( \9128 , \9117 , \9127 );
nor \U$8786 ( \9129 , \9116 , \9128 );
not \U$8787 ( \9130 , \9129 );
and \U$8788 ( \9131 , \9102 , \9130 );
and \U$8789 ( \9132 , \9101 , \9129 );
xor \U$8790 ( \9133 , \8720 , \8728 );
xor \U$8791 ( \9134 , \9133 , \8736 );
not \U$8792 ( \9135 , \8690 );
xor \U$8793 ( \9136 , \8699 , \8709 );
not \U$8794 ( \9137 , \9136 );
or \U$8795 ( \9138 , \9135 , \9137 );
or \U$8796 ( \9139 , \9136 , \8690 );
nand \U$8797 ( \9140 , \9138 , \9139 );
xor \U$8798 ( \9141 , \9134 , \9140 );
not \U$8799 ( \9142 , \8662 );
xor \U$8800 ( \9143 , \8671 , \8681 );
not \U$8801 ( \9144 , \9143 );
or \U$8802 ( \9145 , \9142 , \9144 );
or \U$8803 ( \9146 , \9143 , \8662 );
nand \U$8804 ( \9147 , \9145 , \9146 );
and \U$8805 ( \9148 , \9141 , \9147 );
and \U$8806 ( \9149 , \9134 , \9140 );
or \U$8807 ( \9150 , \9148 , \9149 );
not \U$8808 ( \9151 , \9150 );
nor \U$8809 ( \9152 , \9132 , \9151 );
nor \U$8810 ( \9153 , \9131 , \9152 );
and \U$8811 ( \9154 , \4203 , RI986e620_21);
and \U$8812 ( \9155 , RI986f7f0_59, \4201 );
nor \U$8813 ( \9156 , \9154 , \9155 );
and \U$8814 ( \9157 , \9156 , \3922 );
not \U$8815 ( \9158 , \9156 );
and \U$8816 ( \9159 , \9158 , \4207 );
nor \U$8817 ( \9160 , \9157 , \9159 );
not \U$8818 ( \9161 , \9160 );
and \U$8819 ( \9162 , \5318 , RI986f8e0_61);
and \U$8820 ( \9163 , RI986f430_51, \5316 );
nor \U$8821 ( \9164 , \9162 , \9163 );
and \U$8822 ( \9165 , \9164 , \5322 );
not \U$8823 ( \9166 , \9164 );
and \U$8824 ( \9167 , \9166 , \5052 );
nor \U$8825 ( \9168 , \9165 , \9167 );
not \U$8826 ( \9169 , \9168 );
and \U$8827 ( \9170 , \9161 , \9169 );
and \U$8828 ( \9171 , \9168 , \9160 );
and \U$8829 ( \9172 , \4710 , RI986f700_57);
and \U$8830 ( \9173 , RI986f9d0_63, \4708 );
nor \U$8831 ( \9174 , \9172 , \9173 );
not \U$8832 ( \9175 , \9174 );
not \U$8833 ( \9176 , \4521 );
and \U$8834 ( \9177 , \9175 , \9176 );
and \U$8835 ( \9178 , \9174 , \4519 );
nor \U$8836 ( \9179 , \9177 , \9178 );
nor \U$8837 ( \9180 , \9171 , \9179 );
nor \U$8838 ( \9181 , \9170 , \9180 );
not \U$8839 ( \9182 , \9181 );
and \U$8840 ( \9183 , \5881 , RI986f340_49);
and \U$8841 ( \9184 , RI986f520_53, \5879 );
nor \U$8842 ( \9185 , \9183 , \9184 );
and \U$8843 ( \9186 , \9185 , \5885 );
not \U$8844 ( \9187 , \9185 );
and \U$8845 ( \9188 , \9187 , \5594 );
nor \U$8846 ( \9189 , \9186 , \9188 );
not \U$8847 ( \9190 , \9189 );
and \U$8848 ( \9191 , \6453 , RI986f610_55);
and \U$8849 ( \9192 , RI986df90_7, \6451 );
nor \U$8850 ( \9193 , \9191 , \9192 );
and \U$8851 ( \9194 , \9193 , \6705 );
not \U$8852 ( \9195 , \9193 );
and \U$8853 ( \9196 , \9195 , \6190 );
nor \U$8854 ( \9197 , \9194 , \9196 );
not \U$8855 ( \9198 , \9197 );
and \U$8856 ( \9199 , \9190 , \9198 );
and \U$8857 ( \9200 , \9197 , \9189 );
and \U$8858 ( \9201 , \7079 , RI986dea0_5);
and \U$8859 ( \9202 , RI986ddb0_3, \7077 );
nor \U$8860 ( \9203 , \9201 , \9202 );
and \U$8861 ( \9204 , \9203 , \6709 );
not \U$8862 ( \9205 , \9203 );
and \U$8863 ( \9206 , \9205 , \6710 );
nor \U$8864 ( \9207 , \9204 , \9206 );
nor \U$8865 ( \9208 , \9200 , \9207 );
nor \U$8866 ( \9209 , \9199 , \9208 );
not \U$8867 ( \9210 , \9209 );
and \U$8868 ( \9211 , \9182 , \9210 );
and \U$8869 ( \9212 , \9181 , \9209 );
and \U$8870 ( \9213 , \7729 , RI986dcc0_1);
and \U$8871 ( \9214 , RI986e170_11, \7727 );
nor \U$8872 ( \9215 , \9213 , \9214 );
and \U$8873 ( \9216 , \9215 , \7733 );
not \U$8874 ( \9217 , \9215 );
and \U$8875 ( \9218 , \9217 , \7480 );
nor \U$8876 ( \9219 , \9216 , \9218 );
not \U$8877 ( \9220 , \9219 );
and \U$8878 ( \9221 , \8486 , RI986e080_9);
and \U$8879 ( \9222 , RI986e260_13, \8484 );
nor \U$8880 ( \9223 , \9221 , \9222 );
and \U$8881 ( \9224 , \9223 , \8051 );
not \U$8882 ( \9225 , \9223 );
and \U$8883 ( \9226 , \9225 , \8050 );
nor \U$8884 ( \9227 , \9224 , \9226 );
not \U$8885 ( \9228 , \9227 );
and \U$8886 ( \9229 , \9220 , \9228 );
and \U$8887 ( \9230 , \9227 , \9219 );
and \U$8888 ( \9231 , RI9872e50_175, RI9872ec8_176);
not \U$8889 ( \9232 , RI9872f40_177);
and \U$8890 ( \9233 , \9232 , RI9872ec8_176);
nor \U$8891 ( \9234 , \9232 , RI9872ec8_176);
or \U$8892 ( \9235 , \9233 , \9234 );
nor \U$8893 ( \9236 , RI9872e50_175, RI9872ec8_176);
nor \U$8894 ( \9237 , \9231 , \9235 , \9236 );
nand \U$8895 ( \9238 , RI986e350_15, \9237 );
and \U$8896 ( \9239 , \9238 , \8836 );
not \U$8897 ( \9240 , \9238 );
not \U$8898 ( \9241 , \8836 );
and \U$8899 ( \9242 , \9240 , \9241 );
nor \U$8900 ( \9243 , \9239 , \9242 );
nor \U$8901 ( \9244 , \9230 , \9243 );
nor \U$8902 ( \9245 , \9229 , \9244 );
nor \U$8903 ( \9246 , \9212 , \9245 );
nor \U$8904 ( \9247 , \9211 , \9246 );
not \U$8905 ( \9248 , \9247 );
not \U$8906 ( \9249 , \1128 );
and \U$8907 ( \9250 , \1293 , RI98715f0_123);
and \U$8908 ( \9251 , RI986ead0_31, \1291 );
nor \U$8909 ( \9252 , \9250 , \9251 );
not \U$8910 ( \9253 , \9252 );
or \U$8911 ( \9254 , \9249 , \9253 );
or \U$8912 ( \9255 , \9252 , \1128 );
nand \U$8913 ( \9256 , \9254 , \9255 );
and \U$8914 ( \9257 , \1329 , RI986e9e0_29);
and \U$8915 ( \9258 , RI986e8f0_27, \1327 );
nor \U$8916 ( \9259 , \9257 , \9258 );
and \U$8917 ( \9260 , \9259 , \1336 );
not \U$8918 ( \9261 , \9259 );
and \U$8919 ( \9262 , \9261 , \1337 );
nor \U$8920 ( \9263 , \9260 , \9262 );
xor \U$8921 ( \9264 , \9256 , \9263 );
and \U$8922 ( \9265 , \776 , RI98717d0_127);
and \U$8923 ( \9266 , RI9871500_121, \774 );
nor \U$8924 ( \9267 , \9265 , \9266 );
and \U$8925 ( \9268 , \9267 , \474 );
not \U$8926 ( \9269 , \9267 );
and \U$8927 ( \9270 , \9269 , \451 );
nor \U$8928 ( \9271 , \9268 , \9270 );
and \U$8929 ( \9272 , \9264 , \9271 );
and \U$8930 ( \9273 , \9256 , \9263 );
nor \U$8931 ( \9274 , \9272 , \9273 );
not \U$8932 ( \9275 , \9274 );
not \U$8933 ( \9276 , \2935 );
and \U$8934 ( \9277 , \3254 , RI986f160_45);
and \U$8935 ( \9278 , RI986e530_19, \3252 );
nor \U$8936 ( \9279 , \9277 , \9278 );
not \U$8937 ( \9280 , \9279 );
or \U$8938 ( \9281 , \9276 , \9280 );
or \U$8939 ( \9282 , \9279 , \2935 );
nand \U$8940 ( \9283 , \9281 , \9282 );
not \U$8941 ( \9284 , \3918 );
and \U$8942 ( \9285 , \3683 , RI986e440_17);
and \U$8943 ( \9286 , RI986e710_23, \3681 );
nor \U$8944 ( \9287 , \9285 , \9286 );
not \U$8945 ( \9288 , \9287 );
or \U$8946 ( \9289 , \9284 , \9288 );
or \U$8947 ( \9290 , \9287 , \3412 );
nand \U$8948 ( \9291 , \9289 , \9290 );
xor \U$8949 ( \9292 , \9283 , \9291 );
and \U$8950 ( \9293 , \2464 , RI986ef80_41);
and \U$8951 ( \9294 , RI986f250_47, \2462 );
nor \U$8952 ( \9295 , \9293 , \9294 );
and \U$8953 ( \9296 , \9295 , \2468 );
not \U$8954 ( \9297 , \9295 );
and \U$8955 ( \9298 , \9297 , \2263 );
nor \U$8956 ( \9299 , \9296 , \9298 );
and \U$8957 ( \9300 , \9292 , \9299 );
and \U$8958 ( \9301 , \9283 , \9291 );
nor \U$8959 ( \9302 , \9300 , \9301 );
not \U$8960 ( \9303 , \9302 );
and \U$8961 ( \9304 , \9275 , \9303 );
and \U$8962 ( \9305 , \9274 , \9302 );
and \U$8963 ( \9306 , \1311 , RI986e800_25);
and \U$8964 ( \9307 , RI986ee90_39, \1309 );
nor \U$8965 ( \9308 , \9306 , \9307 );
and \U$8966 ( \9309 , \9308 , \1315 );
not \U$8967 ( \9310 , \9308 );
and \U$8968 ( \9311 , \9310 , \1458 );
nor \U$8969 ( \9312 , \9309 , \9311 );
not \U$8970 ( \9313 , \9312 );
and \U$8971 ( \9314 , \2042 , RI986eda0_37);
and \U$8972 ( \9315 , RI986ebc0_33, \2040 );
nor \U$8973 ( \9316 , \9314 , \9315 );
not \U$8974 ( \9317 , \9316 );
not \U$8975 ( \9318 , \2034 );
and \U$8976 ( \9319 , \9317 , \9318 );
and \U$8977 ( \9320 , \9316 , \1462 );
nor \U$8978 ( \9321 , \9319 , \9320 );
not \U$8979 ( \9322 , \9321 );
and \U$8980 ( \9323 , \9313 , \9322 );
and \U$8981 ( \9324 , \9321 , \9312 );
and \U$8982 ( \9325 , \2274 , RI986ecb0_35);
and \U$8983 ( \9326 , RI986f070_43, \2272 );
nor \U$8984 ( \9327 , \9325 , \9326 );
and \U$8985 ( \9328 , \9327 , \2031 );
not \U$8986 ( \9329 , \9327 );
and \U$8987 ( \9330 , \9329 , \2030 );
nor \U$8988 ( \9331 , \9328 , \9330 );
nor \U$8989 ( \9332 , \9324 , \9331 );
nor \U$8990 ( \9333 , \9323 , \9332 );
nor \U$8991 ( \9334 , \9305 , \9333 );
nor \U$8992 ( \9335 , \9304 , \9334 );
not \U$8993 ( \9336 , \9335 );
and \U$8994 ( \9337 , \9248 , \9336 );
and \U$8995 ( \9338 , \9247 , \9335 );
and \U$8996 ( \9339 , \438 , RI9871410_119);
and \U$8997 ( \9340 , RI98716e0_125, \436 );
nor \U$8998 ( \9341 , \9339 , \9340 );
and \U$8999 ( \9342 , \9341 , \444 );
not \U$9000 ( \9343 , \9341 );
and \U$9001 ( \9344 , \9343 , \443 );
nor \U$9002 ( \9345 , \9342 , \9344 );
not \U$9003 ( \9346 , \456 );
and \U$9004 ( \9347 , \465 , RI9871140_113);
and \U$9005 ( \9348 , RI9871320_117, \463 );
nor \U$9006 ( \9349 , \9347 , \9348 );
not \U$9007 ( \9350 , \9349 );
or \U$9008 ( \9351 , \9346 , \9350 );
or \U$9009 ( \9352 , \9349 , \454 );
nand \U$9010 ( \9353 , \9351 , \9352 );
xor \U$9011 ( \9354 , \9345 , \9353 );
not \U$9012 ( \9355 , \365 );
and \U$9013 ( \9356 , \376 , RI9870c90_103);
and \U$9014 ( \9357 , RI9871230_115, \374 );
nor \U$9015 ( \9358 , \9356 , \9357 );
not \U$9016 ( \9359 , \9358 );
or \U$9017 ( \9360 , \9355 , \9359 );
or \U$9018 ( \9361 , \9358 , \367 );
nand \U$9019 ( \9362 , \9360 , \9361 );
and \U$9020 ( \9363 , \9354 , \9362 );
and \U$9021 ( \9364 , \9345 , \9353 );
or \U$9022 ( \9365 , \9363 , \9364 );
not \U$9023 ( \9366 , \487 );
and \U$9024 ( \9367 , \395 , RI9870ba0_101);
and \U$9025 ( \9368 , RI9871050_111, \393 );
nor \U$9026 ( \9369 , \9367 , \9368 );
not \U$9027 ( \9370 , \9369 );
or \U$9028 ( \9371 , \9366 , \9370 );
or \U$9029 ( \9372 , \9369 , \487 );
nand \U$9030 ( \9373 , \9371 , \9372 );
not \U$9031 ( \9374 , \361 );
and \U$9032 ( \9375 , \354 , RI98709c0_97);
and \U$9033 ( \9376 , RI9870e70_107, \352 );
nor \U$9034 ( \9377 , \9375 , \9376 );
not \U$9035 ( \9378 , \9377 );
or \U$9036 ( \9379 , \9374 , \9378 );
or \U$9037 ( \9380 , \9377 , \361 );
nand \U$9038 ( \9381 , \9379 , \9380 );
xor \U$9039 ( \9382 , \9373 , \9381 );
and \U$9040 ( \9383 , \416 , RI9870ab0_99);
and \U$9041 ( \9384 , RI9870d80_105, \414 );
nor \U$9042 ( \9385 , \9383 , \9384 );
and \U$9043 ( \9386 , \9385 , \422 );
not \U$9044 ( \9387 , \9385 );
and \U$9045 ( \9388 , \9387 , \421 );
nor \U$9046 ( \9389 , \9386 , \9388 );
and \U$9047 ( \9390 , \9382 , \9389 );
and \U$9048 ( \9391 , \9373 , \9381 );
or \U$9049 ( \9392 , \9390 , \9391 );
xor \U$9050 ( \9393 , \9365 , \9392 );
nand \U$9051 ( \9394 , RI9870f60_109, RI9871fc8_144);
not \U$9052 ( \9395 , \9394 );
and \U$9053 ( \9396 , \9393 , \9395 );
and \U$9054 ( \9397 , \9365 , \9392 );
or \U$9055 ( \9398 , \9396 , \9397 );
not \U$9056 ( \9399 , \9398 );
nor \U$9057 ( \9400 , \9338 , \9399 );
nor \U$9058 ( \9401 , \9337 , \9400 );
xor \U$9059 ( \9402 , \9153 , \9401 );
not \U$9060 ( \9403 , \8882 );
not \U$9061 ( \9404 , \8894 );
or \U$9062 ( \9405 , \9403 , \9404 );
or \U$9063 ( \9406 , \8882 , \8894 );
nand \U$9064 ( \9407 , \9405 , \9406 );
not \U$9065 ( \9408 , \9407 );
not \U$9066 ( \9409 , \8884 );
and \U$9067 ( \9410 , \9408 , \9409 );
and \U$9068 ( \9411 , \9407 , \8884 );
nor \U$9069 ( \9412 , \9410 , \9411 );
not \U$9070 ( \9413 , \9412 );
not \U$9071 ( \9414 , \8898 );
not \U$9072 ( \9415 , \8901 );
and \U$9073 ( \9416 , \9414 , \9415 );
and \U$9074 ( \9417 , \8898 , \8901 );
nor \U$9075 ( \9418 , \9416 , \9417 );
not \U$9076 ( \9419 , \9418 );
and \U$9077 ( \9420 , \9413 , \9419 );
and \U$9078 ( \9421 , \9412 , \9418 );
not \U$9079 ( \9422 , \8925 );
xor \U$9080 ( \9423 , \8913 , \8919 );
not \U$9081 ( \9424 , \9423 );
or \U$9082 ( \9425 , \9422 , \9424 );
or \U$9083 ( \9426 , \9423 , \8925 );
nand \U$9084 ( \9427 , \9425 , \9426 );
not \U$9085 ( \9428 , \9427 );
nor \U$9086 ( \9429 , \9421 , \9428 );
nor \U$9087 ( \9430 , \9420 , \9429 );
and \U$9088 ( \9431 , \9402 , \9430 );
and \U$9089 ( \9432 , \9153 , \9401 );
or \U$9090 ( \9433 , \9431 , \9432 );
xor \U$9091 ( \9434 , \8742 , \8801 );
xor \U$9092 ( \9435 , \9434 , \8877 );
not \U$9093 ( \9436 , \9435 );
not \U$9094 ( \9437 , \8902 );
not \U$9095 ( \9438 , \8896 );
not \U$9096 ( \9439 , \8927 );
or \U$9097 ( \9440 , \9438 , \9439 );
or \U$9098 ( \9441 , \8927 , \8896 );
nand \U$9099 ( \9442 , \9440 , \9441 );
not \U$9100 ( \9443 , \9442 );
or \U$9101 ( \9444 , \9437 , \9443 );
or \U$9102 ( \9445 , \9442 , \8902 );
nand \U$9103 ( \9446 , \9444 , \9445 );
nand \U$9104 ( \9447 , \9436 , \9446 );
xor \U$9105 ( \9448 , \9433 , \9447 );
xor \U$9106 ( \9449 , \8827 , \8847 );
xor \U$9107 ( \9450 , \9449 , \8874 );
not \U$9108 ( \9451 , \9450 );
and \U$9109 ( \9452 , \8771 , \8800 );
nor \U$9110 ( \9453 , \9452 , \8801 );
not \U$9111 ( \9454 , \9453 );
and \U$9112 ( \9455 , \9451 , \9454 );
and \U$9113 ( \9456 , \9450 , \9453 );
xor \U$9114 ( \9457 , \8683 , \8711 );
xor \U$9115 ( \9458 , \9457 , \8739 );
nor \U$9116 ( \9459 , \9456 , \9458 );
nor \U$9117 ( \9460 , \9455 , \9459 );
xor \U$9118 ( \9461 , \8640 , \8642 );
xor \U$9119 ( \9462 , \9461 , \8645 );
and \U$9120 ( \9463 , \9460 , \9462 );
xor \U$9121 ( \9464 , \8565 , \8567 );
xor \U$9122 ( \9465 , \9464 , \8570 );
xor \U$9123 ( \9466 , \8932 , \8939 );
xor \U$9124 ( \9467 , \9465 , \9466 );
xor \U$9125 ( \9468 , \8640 , \8642 );
xor \U$9126 ( \9469 , \9468 , \8645 );
and \U$9127 ( \9470 , \9467 , \9469 );
and \U$9128 ( \9471 , \9460 , \9467 );
or \U$9129 ( \9472 , \9463 , \9470 , \9471 );
and \U$9130 ( \9473 , \9448 , \9472 );
and \U$9131 ( \9474 , \9433 , \9447 );
or \U$9132 ( \9475 , \9473 , \9474 );
xor \U$9133 ( \9476 , \9089 , \9475 );
xnor \U$9134 ( \9477 , \8975 , \8969 );
not \U$9135 ( \9478 , \9477 );
not \U$9136 ( \9479 , \8991 );
and \U$9137 ( \9480 , \9478 , \9479 );
and \U$9138 ( \9481 , \9477 , \8991 );
nor \U$9139 ( \9482 , \9480 , \9481 );
and \U$9140 ( \9483 , \9476 , \9482 );
and \U$9141 ( \9484 , \9089 , \9475 );
or \U$9142 ( \9485 , \9483 , \9484 );
nor \U$9143 ( \9486 , \9075 , \9485 );
nor \U$9144 ( \9487 , \9072 , \9486 );
nor \U$9145 ( \9488 , \9067 , \9487 );
and \U$9146 ( \9489 , \9064 , \9488 );
xor \U$9147 ( \9490 , \9488 , \9064 );
and \U$9148 ( \9491 , \8486 , RI986dcc0_1);
and \U$9149 ( \9492 , RI986e170_11, \8484 );
nor \U$9150 ( \9493 , \9491 , \9492 );
and \U$9151 ( \9494 , \9493 , \8050 );
not \U$9152 ( \9495 , \9493 );
and \U$9153 ( \9496 , \9495 , \8051 );
nor \U$9154 ( \9497 , \9494 , \9496 );
and \U$9155 ( \9498 , RI9872f40_177, RI9872fb8_178);
not \U$9156 ( \9499 , RI9872fb8_178);
nor \U$9157 ( \9500 , \9499 , RI9873030_179);
not \U$9158 ( \9501 , RI9873030_179);
nor \U$9159 ( \9502 , \9501 , RI9872fb8_178);
or \U$9160 ( \9503 , \9500 , \9502 );
nor \U$9161 ( \9504 , RI9872f40_177, RI9872fb8_178);
nor \U$9162 ( \9505 , \9498 , \9503 , \9504 );
nand \U$9163 ( \9506 , RI986e350_15, \9505 );
not \U$9164 ( \9507 , RI9873030_179);
not \U$9165 ( \9508 , RI9872fb8_178);
or \U$9166 ( \9509 , \9507 , \9508 );
nand \U$9167 ( \9510 , \9509 , RI9872f40_177);
and \U$9168 ( \9511 , \9506 , \9510 );
not \U$9169 ( \9512 , \9506 );
not \U$9170 ( \9513 , \9510 );
and \U$9171 ( \9514 , \9512 , \9513 );
nor \U$9172 ( \9515 , \9511 , \9514 );
xor \U$9173 ( \9516 , \9497 , \9515 );
and \U$9174 ( \9517 , \9237 , RI986e080_9);
and \U$9175 ( \9518 , RI986e260_13, \9235 );
nor \U$9176 ( \9519 , \9517 , \9518 );
and \U$9177 ( \9520 , \9519 , \9241 );
not \U$9178 ( \9521 , \9519 );
and \U$9179 ( \9522 , \9521 , \8836 );
nor \U$9180 ( \9523 , \9520 , \9522 );
xor \U$9181 ( \9524 , \9516 , \9523 );
and \U$9182 ( \9525 , \7729 , RI986dea0_5);
and \U$9183 ( \9526 , RI986ddb0_3, \7727 );
nor \U$9184 ( \9527 , \9525 , \9526 );
and \U$9185 ( \9528 , \9527 , \7480 );
not \U$9186 ( \9529 , \9527 );
and \U$9187 ( \9530 , \9529 , \7733 );
nor \U$9188 ( \9531 , \9528 , \9530 );
and \U$9189 ( \9532 , \6453 , RI986f340_49);
and \U$9190 ( \9533 , RI986f520_53, \6451 );
nor \U$9191 ( \9534 , \9532 , \9533 );
and \U$9192 ( \9535 , \9534 , \6190 );
not \U$9193 ( \9536 , \9534 );
and \U$9194 ( \9537 , \9536 , \6705 );
nor \U$9195 ( \9538 , \9535 , \9537 );
xor \U$9196 ( \9539 , \9531 , \9538 );
and \U$9197 ( \9540 , \7079 , RI986f610_55);
and \U$9198 ( \9541 , RI986df90_7, \7077 );
nor \U$9199 ( \9542 , \9540 , \9541 );
and \U$9200 ( \9543 , \9542 , \6710 );
not \U$9201 ( \9544 , \9542 );
and \U$9202 ( \9545 , \9544 , \6709 );
nor \U$9203 ( \9546 , \9543 , \9545 );
xor \U$9204 ( \9547 , \9539 , \9546 );
and \U$9205 ( \9548 , \9524 , \9547 );
and \U$9206 ( \9549 , \5318 , RI986f700_57);
and \U$9207 ( \9550 , RI986f9d0_63, \5316 );
nor \U$9208 ( \9551 , \9549 , \9550 );
and \U$9209 ( \9552 , \9551 , \5052 );
not \U$9210 ( \9553 , \9551 );
and \U$9211 ( \9554 , \9553 , \5322 );
nor \U$9212 ( \9555 , \9552 , \9554 );
not \U$9213 ( \9556 , \4519 );
and \U$9214 ( \9557 , \4710 , RI986e620_21);
and \U$9215 ( \9558 , RI986f7f0_59, \4708 );
nor \U$9216 ( \9559 , \9557 , \9558 );
not \U$9217 ( \9560 , \9559 );
or \U$9218 ( \9561 , \9556 , \9560 );
or \U$9219 ( \9562 , \9559 , \4521 );
nand \U$9220 ( \9563 , \9561 , \9562 );
xor \U$9221 ( \9564 , \9555 , \9563 );
and \U$9222 ( \9565 , \5881 , RI986f8e0_61);
and \U$9223 ( \9566 , RI986f430_51, \5879 );
nor \U$9224 ( \9567 , \9565 , \9566 );
and \U$9225 ( \9568 , \9567 , \5594 );
not \U$9226 ( \9569 , \9567 );
and \U$9227 ( \9570 , \9569 , \5885 );
nor \U$9228 ( \9571 , \9568 , \9570 );
xor \U$9229 ( \9572 , \9564 , \9571 );
xor \U$9230 ( \9573 , \9531 , \9538 );
xor \U$9231 ( \9574 , \9573 , \9546 );
and \U$9232 ( \9575 , \9572 , \9574 );
and \U$9233 ( \9576 , \9524 , \9572 );
or \U$9234 ( \9577 , \9548 , \9575 , \9576 );
not \U$9235 ( \9578 , \454 );
and \U$9236 ( \9579 , \465 , RI9870c90_103);
and \U$9237 ( \9580 , RI9871230_115, \463 );
nor \U$9238 ( \9581 , \9579 , \9580 );
not \U$9239 ( \9582 , \9581 );
or \U$9240 ( \9583 , \9578 , \9582 );
or \U$9241 ( \9584 , \9581 , \454 );
nand \U$9242 ( \9585 , \9583 , \9584 );
and \U$9243 ( \9586 , \776 , RI9871410_119);
and \U$9244 ( \9587 , RI98716e0_125, \774 );
nor \U$9245 ( \9588 , \9586 , \9587 );
and \U$9246 ( \9589 , \9588 , \474 );
not \U$9247 ( \9590 , \9588 );
and \U$9248 ( \9591 , \9590 , \451 );
nor \U$9249 ( \9592 , \9589 , \9591 );
xor \U$9250 ( \9593 , \9585 , \9592 );
and \U$9251 ( \9594 , \438 , RI9871140_113);
and \U$9252 ( \9595 , RI9871320_117, \436 );
nor \U$9253 ( \9596 , \9594 , \9595 );
and \U$9254 ( \9597 , \9596 , \444 );
not \U$9255 ( \9598 , \9596 );
and \U$9256 ( \9599 , \9598 , \443 );
nor \U$9257 ( \9600 , \9597 , \9599 );
xor \U$9258 ( \9601 , \9593 , \9600 );
and \U$9259 ( \9602 , \416 , RI9870150_79);
and \U$9260 ( \9603 , RI9870f60_109, \414 );
nor \U$9261 ( \9604 , \9602 , \9603 );
and \U$9262 ( \9605 , \9604 , \421 );
not \U$9263 ( \9606 , \9604 );
and \U$9264 ( \9607 , \9606 , \422 );
nor \U$9265 ( \9608 , \9605 , \9607 );
nand \U$9266 ( \9609 , RI9870060_77, RI9871fc8_144);
or \U$9267 ( \9610 , \9608 , \9609 );
nand \U$9268 ( \9611 , \9609 , \9608 );
nand \U$9269 ( \9612 , \9610 , \9611 );
xor \U$9270 ( \9613 , \9601 , \9612 );
not \U$9271 ( \9614 , \361 );
and \U$9272 ( \9615 , \354 , RI9870ab0_99);
and \U$9273 ( \9616 , RI9870d80_105, \352 );
nor \U$9274 ( \9617 , \9615 , \9616 );
not \U$9275 ( \9618 , \9617 );
or \U$9276 ( \9619 , \9614 , \9618 );
or \U$9277 ( \9620 , \9617 , \345 );
nand \U$9278 ( \9621 , \9619 , \9620 );
not \U$9279 ( \9622 , \367 );
and \U$9280 ( \9623 , \376 , RI9870ba0_101);
and \U$9281 ( \9624 , RI9871050_111, \374 );
nor \U$9282 ( \9625 , \9623 , \9624 );
not \U$9283 ( \9626 , \9625 );
or \U$9284 ( \9627 , \9622 , \9626 );
or \U$9285 ( \9628 , \9625 , \367 );
nand \U$9286 ( \9629 , \9627 , \9628 );
xor \U$9287 ( \9630 , \9621 , \9629 );
not \U$9288 ( \9631 , \487 );
and \U$9289 ( \9632 , \395 , RI98709c0_97);
and \U$9290 ( \9633 , RI9870e70_107, \393 );
nor \U$9291 ( \9634 , \9632 , \9633 );
not \U$9292 ( \9635 , \9634 );
or \U$9293 ( \9636 , \9631 , \9635 );
or \U$9294 ( \9637 , \9634 , \487 );
nand \U$9295 ( \9638 , \9636 , \9637 );
xor \U$9296 ( \9639 , \9630 , \9638 );
and \U$9297 ( \9640 , \9613 , \9639 );
and \U$9298 ( \9641 , \9601 , \9612 );
or \U$9299 ( \9642 , \9640 , \9641 );
xor \U$9300 ( \9643 , \9577 , \9642 );
and \U$9301 ( \9644 , \2274 , RI986eda0_37);
and \U$9302 ( \9645 , RI986ebc0_33, \2272 );
nor \U$9303 ( \9646 , \9644 , \9645 );
and \U$9304 ( \9647 , \9646 , \2030 );
not \U$9305 ( \9648 , \9646 );
and \U$9306 ( \9649 , \9648 , \2031 );
nor \U$9307 ( \9650 , \9647 , \9649 );
not \U$9308 ( \9651 , \2034 );
and \U$9309 ( \9652 , \2042 , RI986e800_25);
and \U$9310 ( \9653 , RI986ee90_39, \2040 );
nor \U$9311 ( \9654 , \9652 , \9653 );
not \U$9312 ( \9655 , \9654 );
or \U$9313 ( \9656 , \9651 , \9655 );
or \U$9314 ( \9657 , \9654 , \1462 );
nand \U$9315 ( \9658 , \9656 , \9657 );
xor \U$9316 ( \9659 , \9650 , \9658 );
and \U$9317 ( \9660 , \2464 , RI986ecb0_35);
and \U$9318 ( \9661 , RI986f070_43, \2462 );
nor \U$9319 ( \9662 , \9660 , \9661 );
and \U$9320 ( \9663 , \9662 , \2468 );
not \U$9321 ( \9664 , \9662 );
and \U$9322 ( \9665 , \9664 , \2263 );
nor \U$9323 ( \9666 , \9663 , \9665 );
xor \U$9324 ( \9667 , \9659 , \9666 );
and \U$9325 ( \9668 , \1329 , RI98715f0_123);
and \U$9326 ( \9669 , RI986ead0_31, \1327 );
nor \U$9327 ( \9670 , \9668 , \9669 );
and \U$9328 ( \9671 , \9670 , \1336 );
not \U$9329 ( \9672 , \9670 );
and \U$9330 ( \9673 , \9672 , \1337 );
nor \U$9331 ( \9674 , \9671 , \9673 );
not \U$9332 ( \9675 , \1128 );
and \U$9333 ( \9676 , \1293 , RI98717d0_127);
and \U$9334 ( \9677 , RI9871500_121, \1291 );
nor \U$9335 ( \9678 , \9676 , \9677 );
not \U$9336 ( \9679 , \9678 );
or \U$9337 ( \9680 , \9675 , \9679 );
or \U$9338 ( \9681 , \9678 , \1128 );
nand \U$9339 ( \9682 , \9680 , \9681 );
xor \U$9340 ( \9683 , \9674 , \9682 );
and \U$9341 ( \9684 , \1311 , RI986e9e0_29);
and \U$9342 ( \9685 , RI986e8f0_27, \1309 );
nor \U$9343 ( \9686 , \9684 , \9685 );
and \U$9344 ( \9687 , \9686 , \1458 );
not \U$9345 ( \9688 , \9686 );
and \U$9346 ( \9689 , \9688 , \1315 );
nor \U$9347 ( \9690 , \9687 , \9689 );
xor \U$9348 ( \9691 , \9683 , \9690 );
and \U$9349 ( \9692 , \9667 , \9691 );
and \U$9350 ( \9693 , \4203 , RI986e440_17);
and \U$9351 ( \9694 , RI986e710_23, \4201 );
nor \U$9352 ( \9695 , \9693 , \9694 );
and \U$9353 ( \9696 , \9695 , \4207 );
not \U$9354 ( \9697 , \9695 );
and \U$9355 ( \9698 , \9697 , \3922 );
nor \U$9356 ( \9699 , \9696 , \9698 );
not \U$9357 ( \9700 , \2935 );
and \U$9358 ( \9701 , \3254 , RI986ef80_41);
and \U$9359 ( \9702 , RI986f250_47, \3252 );
nor \U$9360 ( \9703 , \9701 , \9702 );
not \U$9361 ( \9704 , \9703 );
or \U$9362 ( \9705 , \9700 , \9704 );
or \U$9363 ( \9706 , \9703 , \2935 );
nand \U$9364 ( \9707 , \9705 , \9706 );
xor \U$9365 ( \9708 , \9699 , \9707 );
not \U$9366 ( \9709 , \3918 );
and \U$9367 ( \9710 , \3683 , RI986f160_45);
and \U$9368 ( \9711 , RI986e530_19, \3681 );
nor \U$9369 ( \9712 , \9710 , \9711 );
not \U$9370 ( \9713 , \9712 );
or \U$9371 ( \9714 , \9709 , \9713 );
or \U$9372 ( \9715 , \9712 , \3412 );
nand \U$9373 ( \9716 , \9714 , \9715 );
xor \U$9374 ( \9717 , \9708 , \9716 );
xor \U$9375 ( \9718 , \9674 , \9682 );
xor \U$9376 ( \9719 , \9718 , \9690 );
and \U$9377 ( \9720 , \9717 , \9719 );
and \U$9378 ( \9721 , \9667 , \9717 );
or \U$9379 ( \9722 , \9692 , \9720 , \9721 );
and \U$9380 ( \9723 , \9643 , \9722 );
and \U$9381 ( \9724 , \9577 , \9642 );
or \U$9382 ( \9725 , \9723 , \9724 );
not \U$9383 ( \9726 , \386 );
and \U$9384 ( \9727 , \395 , RI9870d80_105);
and \U$9385 ( \9728 , RI98709c0_97, \393 );
nor \U$9386 ( \9729 , \9727 , \9728 );
not \U$9387 ( \9730 , \9729 );
or \U$9388 ( \9731 , \9726 , \9730 );
or \U$9389 ( \9732 , \9729 , \386 );
nand \U$9390 ( \9733 , \9731 , \9732 );
not \U$9391 ( \9734 , \456 );
and \U$9392 ( \9735 , \465 , RI9871050_111);
and \U$9393 ( \9736 , RI9870c90_103, \463 );
nor \U$9394 ( \9737 , \9735 , \9736 );
not \U$9395 ( \9738 , \9737 );
or \U$9396 ( \9739 , \9734 , \9738 );
or \U$9397 ( \9740 , \9737 , \454 );
nand \U$9398 ( \9741 , \9739 , \9740 );
xor \U$9399 ( \9742 , \9733 , \9741 );
not \U$9400 ( \9743 , \367 );
and \U$9401 ( \9744 , \376 , RI9870e70_107);
and \U$9402 ( \9745 , RI9870ba0_101, \374 );
nor \U$9403 ( \9746 , \9744 , \9745 );
not \U$9404 ( \9747 , \9746 );
or \U$9405 ( \9748 , \9743 , \9747 );
or \U$9406 ( \9749 , \9746 , \367 );
nand \U$9407 ( \9750 , \9748 , \9749 );
and \U$9408 ( \9751 , \9742 , \9750 );
and \U$9409 ( \9752 , \9733 , \9741 );
or \U$9410 ( \9753 , \9751 , \9752 );
not \U$9411 ( \9754 , \361 );
and \U$9412 ( \9755 , \354 , RI9870f60_109);
and \U$9413 ( \9756 , RI9870ab0_99, \352 );
nor \U$9414 ( \9757 , \9755 , \9756 );
not \U$9415 ( \9758 , \9757 );
or \U$9416 ( \9759 , \9754 , \9758 );
or \U$9417 ( \9760 , \9757 , \361 );
nand \U$9418 ( \9761 , \9759 , \9760 );
not \U$9419 ( \9762 , RI986fe80_73);
nor \U$9420 ( \9763 , \9762 , \407 );
xor \U$9421 ( \9764 , \9761 , \9763 );
and \U$9422 ( \9765 , \416 , RI9870060_77);
and \U$9423 ( \9766 , RI9870150_79, \414 );
nor \U$9424 ( \9767 , \9765 , \9766 );
and \U$9425 ( \9768 , \9767 , \422 );
not \U$9426 ( \9769 , \9767 );
and \U$9427 ( \9770 , \9769 , \421 );
nor \U$9428 ( \9771 , \9768 , \9770 );
and \U$9429 ( \9772 , \9764 , \9771 );
and \U$9430 ( \9773 , \9761 , \9763 );
or \U$9431 ( \9774 , \9772 , \9773 );
xor \U$9432 ( \9775 , \9753 , \9774 );
and \U$9433 ( \9776 , \438 , RI9871230_115);
and \U$9434 ( \9777 , RI9871140_113, \436 );
nor \U$9435 ( \9778 , \9776 , \9777 );
and \U$9436 ( \9779 , \9778 , \444 );
not \U$9437 ( \9780 , \9778 );
and \U$9438 ( \9781 , \9780 , \443 );
nor \U$9439 ( \9782 , \9779 , \9781 );
and \U$9440 ( \9783 , \776 , RI9871320_117);
and \U$9441 ( \9784 , RI9871410_119, \774 );
nor \U$9442 ( \9785 , \9783 , \9784 );
and \U$9443 ( \9786 , \9785 , \474 );
not \U$9444 ( \9787 , \9785 );
and \U$9445 ( \9788 , \9787 , \451 );
nor \U$9446 ( \9789 , \9786 , \9788 );
xor \U$9447 ( \9790 , \9782 , \9789 );
not \U$9448 ( \9791 , \1128 );
and \U$9449 ( \9792 , \1293 , RI98716e0_125);
and \U$9450 ( \9793 , RI98717d0_127, \1291 );
nor \U$9451 ( \9794 , \9792 , \9793 );
not \U$9452 ( \9795 , \9794 );
or \U$9453 ( \9796 , \9791 , \9795 );
or \U$9454 ( \9797 , \9794 , \1301 );
nand \U$9455 ( \9798 , \9796 , \9797 );
and \U$9456 ( \9799 , \9790 , \9798 );
and \U$9457 ( \9800 , \9782 , \9789 );
or \U$9458 ( \9801 , \9799 , \9800 );
and \U$9459 ( \9802 , \9775 , \9801 );
and \U$9460 ( \9803 , \9753 , \9774 );
or \U$9461 ( \9804 , \9802 , \9803 );
and \U$9462 ( \9805 , \5318 , RI986f7f0_59);
and \U$9463 ( \9806 , RI986f700_57, \5316 );
nor \U$9464 ( \9807 , \9805 , \9806 );
and \U$9465 ( \9808 , \9807 , \5052 );
not \U$9466 ( \9809 , \9807 );
and \U$9467 ( \9810 , \9809 , \5322 );
nor \U$9468 ( \9811 , \9808 , \9810 );
and \U$9469 ( \9812 , \5881 , RI986f9d0_63);
and \U$9470 ( \9813 , RI986f8e0_61, \5879 );
nor \U$9471 ( \9814 , \9812 , \9813 );
and \U$9472 ( \9815 , \9814 , \5594 );
not \U$9473 ( \9816 , \9814 );
and \U$9474 ( \9817 , \9816 , \5885 );
nor \U$9475 ( \9818 , \9815 , \9817 );
xor \U$9476 ( \9819 , \9811 , \9818 );
and \U$9477 ( \9820 , \6453 , RI986f430_51);
and \U$9478 ( \9821 , RI986f340_49, \6451 );
nor \U$9479 ( \9822 , \9820 , \9821 );
and \U$9480 ( \9823 , \9822 , \6190 );
not \U$9481 ( \9824 , \9822 );
and \U$9482 ( \9825 , \9824 , \6180 );
nor \U$9483 ( \9826 , \9823 , \9825 );
and \U$9484 ( \9827 , \9819 , \9826 );
and \U$9485 ( \9828 , \9811 , \9818 );
or \U$9486 ( \9829 , \9827 , \9828 );
and \U$9487 ( \9830 , \9237 , RI986e170_11);
and \U$9488 ( \9831 , RI986e080_9, \9235 );
nor \U$9489 ( \9832 , \9830 , \9831 );
and \U$9490 ( \9833 , \9832 , \9241 );
not \U$9491 ( \9834 , \9832 );
and \U$9492 ( \9835 , \9834 , \8836 );
nor \U$9493 ( \9836 , \9833 , \9835 );
not \U$9494 ( \9837 , RI98730a8_180);
not \U$9495 ( \9838 , RI9873120_181);
or \U$9496 ( \9839 , \9837 , \9838 );
nand \U$9497 ( \9840 , \9839 , RI9873030_179);
xor \U$9498 ( \9841 , \9836 , \9840 );
and \U$9499 ( \9842 , \9505 , RI986e260_13);
and \U$9500 ( \9843 , RI986e350_15, \9503 );
nor \U$9501 ( \9844 , \9842 , \9843 );
and \U$9502 ( \9845 , \9844 , \9510 );
not \U$9503 ( \9846 , \9844 );
and \U$9504 ( \9847 , \9846 , \9513 );
nor \U$9505 ( \9848 , \9845 , \9847 );
and \U$9506 ( \9849 , \9841 , \9848 );
and \U$9507 ( \9850 , \9836 , \9840 );
or \U$9508 ( \9851 , \9849 , \9850 );
xor \U$9509 ( \9852 , \9829 , \9851 );
and \U$9510 ( \9853 , \7079 , RI986f520_53);
and \U$9511 ( \9854 , RI986f610_55, \7077 );
nor \U$9512 ( \9855 , \9853 , \9854 );
and \U$9513 ( \9856 , \9855 , \6710 );
not \U$9514 ( \9857 , \9855 );
and \U$9515 ( \9858 , \9857 , \6709 );
nor \U$9516 ( \9859 , \9856 , \9858 );
and \U$9517 ( \9860 , \7729 , RI986df90_7);
and \U$9518 ( \9861 , RI986dea0_5, \7727 );
nor \U$9519 ( \9862 , \9860 , \9861 );
and \U$9520 ( \9863 , \9862 , \7480 );
not \U$9521 ( \9864 , \9862 );
and \U$9522 ( \9865 , \9864 , \7733 );
nor \U$9523 ( \9866 , \9863 , \9865 );
xor \U$9524 ( \9867 , \9859 , \9866 );
and \U$9525 ( \9868 , \8486 , RI986ddb0_3);
and \U$9526 ( \9869 , RI986dcc0_1, \8484 );
nor \U$9527 ( \9870 , \9868 , \9869 );
and \U$9528 ( \9871 , \9870 , \8050 );
not \U$9529 ( \9872 , \9870 );
and \U$9530 ( \9873 , \9872 , \8051 );
nor \U$9531 ( \9874 , \9871 , \9873 );
and \U$9532 ( \9875 , \9867 , \9874 );
and \U$9533 ( \9876 , \9859 , \9866 );
or \U$9534 ( \9877 , \9875 , \9876 );
and \U$9535 ( \9878 , \9852 , \9877 );
and \U$9536 ( \9879 , \9829 , \9851 );
or \U$9537 ( \9880 , \9878 , \9879 );
xor \U$9538 ( \9881 , \9804 , \9880 );
and \U$9539 ( \9882 , \4203 , RI986e530_19);
and \U$9540 ( \9883 , RI986e440_17, \4201 );
nor \U$9541 ( \9884 , \9882 , \9883 );
and \U$9542 ( \9885 , \9884 , \4207 );
not \U$9543 ( \9886 , \9884 );
and \U$9544 ( \9887 , \9886 , \3923 );
nor \U$9545 ( \9888 , \9885 , \9887 );
not \U$9546 ( \9889 , \3918 );
and \U$9547 ( \9890 , \3683 , RI986f250_47);
and \U$9548 ( \9891 , RI986f160_45, \3681 );
nor \U$9549 ( \9892 , \9890 , \9891 );
not \U$9550 ( \9893 , \9892 );
or \U$9551 ( \9894 , \9889 , \9893 );
or \U$9552 ( \9895 , \9892 , \3412 );
nand \U$9553 ( \9896 , \9894 , \9895 );
xor \U$9554 ( \9897 , \9888 , \9896 );
not \U$9555 ( \9898 , \4521 );
and \U$9556 ( \9899 , \4710 , RI986e710_23);
and \U$9557 ( \9900 , RI986e620_21, \4708 );
nor \U$9558 ( \9901 , \9899 , \9900 );
not \U$9559 ( \9902 , \9901 );
or \U$9560 ( \9903 , \9898 , \9902 );
or \U$9561 ( \9904 , \9901 , \4519 );
nand \U$9562 ( \9905 , \9903 , \9904 );
and \U$9563 ( \9906 , \9897 , \9905 );
and \U$9564 ( \9907 , \9888 , \9896 );
or \U$9565 ( \9908 , \9906 , \9907 );
not \U$9566 ( \9909 , \3406 );
and \U$9567 ( \9910 , \3254 , RI986f070_43);
and \U$9568 ( \9911 , RI986ef80_41, \3252 );
nor \U$9569 ( \9912 , \9910 , \9911 );
not \U$9570 ( \9913 , \9912 );
or \U$9571 ( \9914 , \9909 , \9913 );
or \U$9572 ( \9915 , \9912 , \3406 );
nand \U$9573 ( \9916 , \9914 , \9915 );
and \U$9574 ( \9917 , \2274 , RI986ee90_39);
and \U$9575 ( \9918 , RI986eda0_37, \2272 );
nor \U$9576 ( \9919 , \9917 , \9918 );
and \U$9577 ( \9920 , \9919 , \2030 );
not \U$9578 ( \9921 , \9919 );
and \U$9579 ( \9922 , \9921 , \2031 );
nor \U$9580 ( \9923 , \9920 , \9922 );
xor \U$9581 ( \9924 , \9916 , \9923 );
and \U$9582 ( \9925 , \2464 , RI986ebc0_33);
and \U$9583 ( \9926 , RI986ecb0_35, \2462 );
nor \U$9584 ( \9927 , \9925 , \9926 );
and \U$9585 ( \9928 , \9927 , \2468 );
not \U$9586 ( \9929 , \9927 );
and \U$9587 ( \9930 , \9929 , \2263 );
nor \U$9588 ( \9931 , \9928 , \9930 );
and \U$9589 ( \9932 , \9924 , \9931 );
and \U$9590 ( \9933 , \9916 , \9923 );
or \U$9591 ( \9934 , \9932 , \9933 );
xor \U$9592 ( \9935 , \9908 , \9934 );
and \U$9593 ( \9936 , \1311 , RI986ead0_31);
and \U$9594 ( \9937 , RI986e9e0_29, \1309 );
nor \U$9595 ( \9938 , \9936 , \9937 );
and \U$9596 ( \9939 , \9938 , \1458 );
not \U$9597 ( \9940 , \9938 );
and \U$9598 ( \9941 , \9940 , \1315 );
nor \U$9599 ( \9942 , \9939 , \9941 );
and \U$9600 ( \9943 , \1329 , RI9871500_121);
and \U$9601 ( \9944 , RI98715f0_123, \1327 );
nor \U$9602 ( \9945 , \9943 , \9944 );
and \U$9603 ( \9946 , \9945 , \1336 );
not \U$9604 ( \9947 , \9945 );
and \U$9605 ( \9948 , \9947 , \1337 );
nor \U$9606 ( \9949 , \9946 , \9948 );
xor \U$9607 ( \9950 , \9942 , \9949 );
not \U$9608 ( \9951 , \2034 );
and \U$9609 ( \9952 , \2042 , RI986e8f0_27);
and \U$9610 ( \9953 , RI986e800_25, \2040 );
nor \U$9611 ( \9954 , \9952 , \9953 );
not \U$9612 ( \9955 , \9954 );
or \U$9613 ( \9956 , \9951 , \9955 );
or \U$9614 ( \9957 , \9954 , \1462 );
nand \U$9615 ( \9958 , \9956 , \9957 );
and \U$9616 ( \9959 , \9950 , \9958 );
and \U$9617 ( \9960 , \9942 , \9949 );
or \U$9618 ( \9961 , \9959 , \9960 );
and \U$9619 ( \9962 , \9935 , \9961 );
and \U$9620 ( \9963 , \9908 , \9934 );
or \U$9621 ( \9964 , \9962 , \9963 );
and \U$9622 ( \9965 , \9881 , \9964 );
and \U$9623 ( \9966 , \9804 , \9880 );
or \U$9624 ( \9967 , \9965 , \9966 );
xor \U$9625 ( \9968 , \9725 , \9967 );
and \U$9626 ( \9969 , \776 , RI98716e0_125);
and \U$9627 ( \9970 , RI98717d0_127, \774 );
nor \U$9628 ( \9971 , \9969 , \9970 );
and \U$9629 ( \9972 , \9971 , \474 );
not \U$9630 ( \9973 , \9971 );
and \U$9631 ( \9974 , \9973 , \451 );
nor \U$9632 ( \9975 , \9972 , \9974 );
and \U$9633 ( \9976 , \438 , RI9871320_117);
and \U$9634 ( \9977 , RI9871410_119, \436 );
nor \U$9635 ( \9978 , \9976 , \9977 );
and \U$9636 ( \9979 , \9978 , \444 );
not \U$9637 ( \9980 , \9978 );
and \U$9638 ( \9981 , \9980 , \443 );
nor \U$9639 ( \9982 , \9979 , \9981 );
xor \U$9640 ( \9983 , \9975 , \9982 );
not \U$9641 ( \9984 , \454 );
and \U$9642 ( \9985 , \465 , RI9871230_115);
and \U$9643 ( \9986 , RI9871140_113, \463 );
nor \U$9644 ( \9987 , \9985 , \9986 );
not \U$9645 ( \9988 , \9987 );
or \U$9646 ( \9989 , \9984 , \9988 );
or \U$9647 ( \9990 , \9987 , \456 );
nand \U$9648 ( \9991 , \9989 , \9990 );
xor \U$9649 ( \9992 , \9983 , \9991 );
not \U$9650 ( \9993 , RI9870150_79);
nor \U$9651 ( \9994 , \9993 , \407 );
and \U$9652 ( \9995 , \416 , RI9870f60_109);
and \U$9653 ( \9996 , RI9870ab0_99, \414 );
nor \U$9654 ( \9997 , \9995 , \9996 );
and \U$9655 ( \9998 , \9997 , \422 );
not \U$9656 ( \9999 , \9997 );
and \U$9657 ( \10000 , \9999 , \421 );
nor \U$9658 ( \10001 , \9998 , \10000 );
xor \U$9659 ( \10002 , \9994 , \10001 );
not \U$9660 ( \10003 , \367 );
and \U$9661 ( \10004 , \376 , RI9871050_111);
and \U$9662 ( \10005 , RI9870c90_103, \374 );
nor \U$9663 ( \10006 , \10004 , \10005 );
not \U$9664 ( \10007 , \10006 );
or \U$9665 ( \10008 , \10003 , \10007 );
or \U$9666 ( \10009 , \10006 , \367 );
nand \U$9667 ( \10010 , \10008 , \10009 );
not \U$9668 ( \10011 , \487 );
and \U$9669 ( \10012 , \395 , RI9870e70_107);
and \U$9670 ( \10013 , RI9870ba0_101, \393 );
nor \U$9671 ( \10014 , \10012 , \10013 );
not \U$9672 ( \10015 , \10014 );
or \U$9673 ( \10016 , \10011 , \10015 );
or \U$9674 ( \10017 , \10014 , \386 );
nand \U$9675 ( \10018 , \10016 , \10017 );
xor \U$9676 ( \10019 , \10010 , \10018 );
not \U$9677 ( \10020 , \345 );
and \U$9678 ( \10021 , \354 , RI9870d80_105);
and \U$9679 ( \10022 , RI98709c0_97, \352 );
nor \U$9680 ( \10023 , \10021 , \10022 );
not \U$9681 ( \10024 , \10023 );
or \U$9682 ( \10025 , \10020 , \10024 );
or \U$9683 ( \10026 , \10023 , \345 );
nand \U$9684 ( \10027 , \10025 , \10026 );
xor \U$9685 ( \10028 , \10019 , \10027 );
xor \U$9686 ( \10029 , \10002 , \10028 );
xor \U$9687 ( \10030 , \9992 , \10029 );
and \U$9688 ( \10031 , \9237 , RI986e260_13);
and \U$9689 ( \10032 , RI986e350_15, \9235 );
nor \U$9690 ( \10033 , \10031 , \10032 );
and \U$9691 ( \10034 , \10033 , \9241 );
not \U$9692 ( \10035 , \10033 );
and \U$9693 ( \10036 , \10035 , \8836 );
nor \U$9694 ( \10037 , \10034 , \10036 );
xor \U$9695 ( \10038 , \10037 , \9510 );
and \U$9696 ( \10039 , \8486 , RI986e170_11);
and \U$9697 ( \10040 , RI986e080_9, \8484 );
nor \U$9698 ( \10041 , \10039 , \10040 );
and \U$9699 ( \10042 , \10041 , \8050 );
not \U$9700 ( \10043 , \10041 );
and \U$9701 ( \10044 , \10043 , \8051 );
nor \U$9702 ( \10045 , \10042 , \10044 );
xor \U$9703 ( \10046 , \10038 , \10045 );
not \U$9704 ( \10047 , \4521 );
and \U$9705 ( \10048 , \4710 , RI986f7f0_59);
and \U$9706 ( \10049 , RI986f700_57, \4708 );
nor \U$9707 ( \10050 , \10048 , \10049 );
not \U$9708 ( \10051 , \10050 );
or \U$9709 ( \10052 , \10047 , \10051 );
or \U$9710 ( \10053 , \10050 , \4519 );
nand \U$9711 ( \10054 , \10052 , \10053 );
and \U$9712 ( \10055 , \5318 , RI986f9d0_63);
and \U$9713 ( \10056 , RI986f8e0_61, \5316 );
nor \U$9714 ( \10057 , \10055 , \10056 );
and \U$9715 ( \10058 , \10057 , \5052 );
not \U$9716 ( \10059 , \10057 );
and \U$9717 ( \10060 , \10059 , \5322 );
nor \U$9718 ( \10061 , \10058 , \10060 );
xor \U$9719 ( \10062 , \10054 , \10061 );
and \U$9720 ( \10063 , \5881 , RI986f430_51);
and \U$9721 ( \10064 , RI986f340_49, \5879 );
nor \U$9722 ( \10065 , \10063 , \10064 );
and \U$9723 ( \10066 , \10065 , \5594 );
not \U$9724 ( \10067 , \10065 );
and \U$9725 ( \10068 , \10067 , \5885 );
nor \U$9726 ( \10069 , \10066 , \10068 );
xor \U$9727 ( \10070 , \10062 , \10069 );
xor \U$9728 ( \10071 , \10046 , \10070 );
and \U$9729 ( \10072 , \7079 , RI986df90_7);
and \U$9730 ( \10073 , RI986dea0_5, \7077 );
nor \U$9731 ( \10074 , \10072 , \10073 );
and \U$9732 ( \10075 , \10074 , \6710 );
not \U$9733 ( \10076 , \10074 );
and \U$9734 ( \10077 , \10076 , \6709 );
nor \U$9735 ( \10078 , \10075 , \10077 );
and \U$9736 ( \10079 , \6453 , RI986f520_53);
and \U$9737 ( \10080 , RI986f610_55, \6451 );
nor \U$9738 ( \10081 , \10079 , \10080 );
and \U$9739 ( \10082 , \10081 , \6190 );
not \U$9740 ( \10083 , \10081 );
and \U$9741 ( \10084 , \10083 , \6180 );
nor \U$9742 ( \10085 , \10082 , \10084 );
xor \U$9743 ( \10086 , \10078 , \10085 );
and \U$9744 ( \10087 , \7729 , RI986ddb0_3);
and \U$9745 ( \10088 , RI986dcc0_1, \7727 );
nor \U$9746 ( \10089 , \10087 , \10088 );
and \U$9747 ( \10090 , \10089 , \7480 );
not \U$9748 ( \10091 , \10089 );
and \U$9749 ( \10092 , \10091 , \7733 );
nor \U$9750 ( \10093 , \10090 , \10092 );
xor \U$9751 ( \10094 , \10086 , \10093 );
xor \U$9752 ( \10095 , \10071 , \10094 );
and \U$9753 ( \10096 , \10030 , \10095 );
not \U$9754 ( \10097 , \1128 );
and \U$9755 ( \10098 , \1293 , RI9871500_121);
and \U$9756 ( \10099 , RI98715f0_123, \1291 );
nor \U$9757 ( \10100 , \10098 , \10099 );
not \U$9758 ( \10101 , \10100 );
or \U$9759 ( \10102 , \10097 , \10101 );
or \U$9760 ( \10103 , \10100 , \1128 );
nand \U$9761 ( \10104 , \10102 , \10103 );
and \U$9762 ( \10105 , \1329 , RI986ead0_31);
and \U$9763 ( \10106 , RI986e9e0_29, \1327 );
nor \U$9764 ( \10107 , \10105 , \10106 );
and \U$9765 ( \10108 , \10107 , \1336 );
not \U$9766 ( \10109 , \10107 );
and \U$9767 ( \10110 , \10109 , \1337 );
nor \U$9768 ( \10111 , \10108 , \10110 );
xor \U$9769 ( \10112 , \10104 , \10111 );
and \U$9770 ( \10113 , \1311 , RI986e8f0_27);
and \U$9771 ( \10114 , RI986e800_25, \1309 );
nor \U$9772 ( \10115 , \10113 , \10114 );
and \U$9773 ( \10116 , \10115 , \1458 );
not \U$9774 ( \10117 , \10115 );
and \U$9775 ( \10118 , \10117 , \1315 );
nor \U$9776 ( \10119 , \10116 , \10118 );
xor \U$9777 ( \10120 , \10112 , \10119 );
not \U$9778 ( \10121 , \1462 );
and \U$9779 ( \10122 , \2042 , RI986ee90_39);
and \U$9780 ( \10123 , RI986eda0_37, \2040 );
nor \U$9781 ( \10124 , \10122 , \10123 );
not \U$9782 ( \10125 , \10124 );
or \U$9783 ( \10126 , \10121 , \10125 );
or \U$9784 ( \10127 , \10124 , \2034 );
nand \U$9785 ( \10128 , \10126 , \10127 );
and \U$9786 ( \10129 , \2274 , RI986ebc0_33);
and \U$9787 ( \10130 , RI986ecb0_35, \2272 );
nor \U$9788 ( \10131 , \10129 , \10130 );
and \U$9789 ( \10132 , \10131 , \2030 );
not \U$9790 ( \10133 , \10131 );
and \U$9791 ( \10134 , \10133 , \2031 );
nor \U$9792 ( \10135 , \10132 , \10134 );
xor \U$9793 ( \10136 , \10128 , \10135 );
and \U$9794 ( \10137 , \2464 , RI986f070_43);
and \U$9795 ( \10138 , RI986ef80_41, \2462 );
nor \U$9796 ( \10139 , \10137 , \10138 );
and \U$9797 ( \10140 , \10139 , \2468 );
not \U$9798 ( \10141 , \10139 );
and \U$9799 ( \10142 , \10141 , \2263 );
nor \U$9800 ( \10143 , \10140 , \10142 );
xor \U$9801 ( \10144 , \10136 , \10143 );
not \U$9802 ( \10145 , \2935 );
and \U$9803 ( \10146 , \3254 , RI986f250_47);
and \U$9804 ( \10147 , RI986f160_45, \3252 );
nor \U$9805 ( \10148 , \10146 , \10147 );
not \U$9806 ( \10149 , \10148 );
or \U$9807 ( \10150 , \10145 , \10149 );
or \U$9808 ( \10151 , \10148 , \3406 );
nand \U$9809 ( \10152 , \10150 , \10151 );
not \U$9810 ( \10153 , \3918 );
and \U$9811 ( \10154 , \3683 , RI986e530_19);
and \U$9812 ( \10155 , RI986e440_17, \3681 );
nor \U$9813 ( \10156 , \10154 , \10155 );
not \U$9814 ( \10157 , \10156 );
or \U$9815 ( \10158 , \10153 , \10157 );
or \U$9816 ( \10159 , \10156 , \3412 );
nand \U$9817 ( \10160 , \10158 , \10159 );
xor \U$9818 ( \10161 , \10152 , \10160 );
and \U$9819 ( \10162 , \4203 , RI986e710_23);
and \U$9820 ( \10163 , RI986e620_21, \4201 );
nor \U$9821 ( \10164 , \10162 , \10163 );
and \U$9822 ( \10165 , \10164 , \4207 );
not \U$9823 ( \10166 , \10164 );
and \U$9824 ( \10167 , \10166 , \3922 );
nor \U$9825 ( \10168 , \10165 , \10167 );
xor \U$9826 ( \10169 , \10161 , \10168 );
xor \U$9827 ( \10170 , \10144 , \10169 );
xor \U$9828 ( \10171 , \10120 , \10170 );
xor \U$9829 ( \10172 , \10046 , \10070 );
xor \U$9830 ( \10173 , \10172 , \10094 );
and \U$9831 ( \10174 , \10171 , \10173 );
and \U$9832 ( \10175 , \10030 , \10171 );
or \U$9833 ( \10176 , \10096 , \10174 , \10175 );
and \U$9834 ( \10177 , \9968 , \10176 );
and \U$9835 ( \10178 , \9725 , \9967 );
or \U$9836 ( \10179 , \10177 , \10178 );
xor \U$9837 ( \10180 , \9650 , \9658 );
and \U$9838 ( \10181 , \10180 , \9666 );
and \U$9839 ( \10182 , \9650 , \9658 );
or \U$9840 ( \10183 , \10181 , \10182 );
xor \U$9841 ( \10184 , \9674 , \9682 );
and \U$9842 ( \10185 , \10184 , \9690 );
and \U$9843 ( \10186 , \9674 , \9682 );
or \U$9844 ( \10187 , \10185 , \10186 );
xor \U$9845 ( \10188 , \10183 , \10187 );
xor \U$9846 ( \10189 , \9699 , \9707 );
and \U$9847 ( \10190 , \10189 , \9716 );
and \U$9848 ( \10191 , \9699 , \9707 );
or \U$9849 ( \10192 , \10190 , \10191 );
and \U$9850 ( \10193 , \10188 , \10192 );
and \U$9851 ( \10194 , \10183 , \10187 );
or \U$9852 ( \10195 , \10193 , \10194 );
xor \U$9853 ( \10196 , \9621 , \9629 );
and \U$9854 ( \10197 , \10196 , \9638 );
and \U$9855 ( \10198 , \9621 , \9629 );
or \U$9856 ( \10199 , \10197 , \10198 );
xor \U$9857 ( \10200 , \10199 , \9611 );
xor \U$9858 ( \10201 , \9585 , \9592 );
and \U$9859 ( \10202 , \10201 , \9600 );
and \U$9860 ( \10203 , \9585 , \9592 );
or \U$9861 ( \10204 , \10202 , \10203 );
and \U$9862 ( \10205 , \10200 , \10204 );
and \U$9863 ( \10206 , \10199 , \9611 );
or \U$9864 ( \10207 , \10205 , \10206 );
xor \U$9865 ( \10208 , \10195 , \10207 );
xor \U$9866 ( \10209 , \9531 , \9538 );
and \U$9867 ( \10210 , \10209 , \9546 );
and \U$9868 ( \10211 , \9531 , \9538 );
or \U$9869 ( \10212 , \10210 , \10211 );
xor \U$9870 ( \10213 , \9497 , \9515 );
and \U$9871 ( \10214 , \10213 , \9523 );
and \U$9872 ( \10215 , \9497 , \9515 );
or \U$9873 ( \10216 , \10214 , \10215 );
xor \U$9874 ( \10217 , \10212 , \10216 );
xor \U$9875 ( \10218 , \9555 , \9563 );
and \U$9876 ( \10219 , \10218 , \9571 );
and \U$9877 ( \10220 , \9555 , \9563 );
or \U$9878 ( \10221 , \10219 , \10220 );
and \U$9879 ( \10222 , \10217 , \10221 );
and \U$9880 ( \10223 , \10212 , \10216 );
or \U$9881 ( \10224 , \10222 , \10223 );
xor \U$9882 ( \10225 , \10208 , \10224 );
xor \U$9883 ( \10226 , \10046 , \10070 );
and \U$9884 ( \10227 , \10226 , \10094 );
and \U$9885 ( \10228 , \10046 , \10070 );
or \U$9886 ( \10229 , \10227 , \10228 );
xor \U$9887 ( \10230 , \9975 , \9982 );
xor \U$9888 ( \10231 , \10230 , \9991 );
and \U$9889 ( \10232 , \10002 , \10231 );
xor \U$9890 ( \10233 , \9975 , \9982 );
xor \U$9891 ( \10234 , \10233 , \9991 );
and \U$9892 ( \10235 , \10028 , \10234 );
and \U$9893 ( \10236 , \10002 , \10028 );
or \U$9894 ( \10237 , \10232 , \10235 , \10236 );
xor \U$9895 ( \10238 , \10229 , \10237 );
xor \U$9896 ( \10239 , \10104 , \10111 );
xor \U$9897 ( \10240 , \10239 , \10119 );
and \U$9898 ( \10241 , \10144 , \10240 );
xor \U$9899 ( \10242 , \10104 , \10111 );
xor \U$9900 ( \10243 , \10242 , \10119 );
and \U$9901 ( \10244 , \10169 , \10243 );
and \U$9902 ( \10245 , \10144 , \10169 );
or \U$9903 ( \10246 , \10241 , \10244 , \10245 );
xor \U$9904 ( \10247 , \10238 , \10246 );
and \U$9905 ( \10248 , \10225 , \10247 );
xor \U$9906 ( \10249 , \10179 , \10248 );
xor \U$9907 ( \10250 , \10199 , \9611 );
xor \U$9908 ( \10251 , \10250 , \10204 );
xor \U$9909 ( \10252 , \10212 , \10216 );
xor \U$9910 ( \10253 , \10252 , \10221 );
xor \U$9911 ( \10254 , \10251 , \10253 );
xor \U$9912 ( \10255 , \10183 , \10187 );
xor \U$9913 ( \10256 , \10255 , \10192 );
and \U$9914 ( \10257 , \10254 , \10256 );
and \U$9915 ( \10258 , \10251 , \10253 );
or \U$9916 ( \10259 , \10257 , \10258 );
xor \U$9917 ( \10260 , \10010 , \10018 );
and \U$9918 ( \10261 , \10260 , \10027 );
and \U$9919 ( \10262 , \10010 , \10018 );
or \U$9920 ( \10263 , \10261 , \10262 );
and \U$9921 ( \10264 , \9994 , \10001 );
xor \U$9922 ( \10265 , \10263 , \10264 );
xor \U$9923 ( \10266 , \9975 , \9982 );
and \U$9924 ( \10267 , \10266 , \9991 );
and \U$9925 ( \10268 , \9975 , \9982 );
or \U$9926 ( \10269 , \10267 , \10268 );
xor \U$9927 ( \10270 , \10265 , \10269 );
xor \U$9928 ( \10271 , \10152 , \10160 );
and \U$9929 ( \10272 , \10271 , \10168 );
and \U$9930 ( \10273 , \10152 , \10160 );
or \U$9931 ( \10274 , \10272 , \10273 );
xor \U$9932 ( \10275 , \10128 , \10135 );
and \U$9933 ( \10276 , \10275 , \10143 );
and \U$9934 ( \10277 , \10128 , \10135 );
or \U$9935 ( \10278 , \10276 , \10277 );
xor \U$9936 ( \10279 , \10274 , \10278 );
xor \U$9937 ( \10280 , \10104 , \10111 );
and \U$9938 ( \10281 , \10280 , \10119 );
and \U$9939 ( \10282 , \10104 , \10111 );
or \U$9940 ( \10283 , \10281 , \10282 );
xor \U$9941 ( \10284 , \10279 , \10283 );
xor \U$9942 ( \10285 , \10270 , \10284 );
xor \U$9943 ( \10286 , \10054 , \10061 );
and \U$9944 ( \10287 , \10286 , \10069 );
and \U$9945 ( \10288 , \10054 , \10061 );
or \U$9946 ( \10289 , \10287 , \10288 );
xor \U$9947 ( \10290 , \10037 , \9510 );
and \U$9948 ( \10291 , \10290 , \10045 );
and \U$9949 ( \10292 , \10037 , \9510 );
or \U$9950 ( \10293 , \10291 , \10292 );
xor \U$9951 ( \10294 , \10289 , \10293 );
xor \U$9952 ( \10295 , \10078 , \10085 );
and \U$9953 ( \10296 , \10295 , \10093 );
and \U$9954 ( \10297 , \10078 , \10085 );
or \U$9955 ( \10298 , \10296 , \10297 );
xor \U$9956 ( \10299 , \10294 , \10298 );
xor \U$9957 ( \10300 , \10285 , \10299 );
and \U$9958 ( \10301 , \10259 , \10300 );
not \U$9959 ( \10302 , \9219 );
xor \U$9960 ( \10303 , \9243 , \9227 );
not \U$9961 ( \10304 , \10303 );
or \U$9962 ( \10305 , \10302 , \10304 );
or \U$9963 ( \10306 , \10303 , \9219 );
nand \U$9964 ( \10307 , \10305 , \10306 );
not \U$9965 ( \10308 , \9160 );
xor \U$9966 ( \10309 , \9179 , \9168 );
not \U$9967 ( \10310 , \10309 );
or \U$9968 ( \10311 , \10308 , \10310 );
or \U$9969 ( \10312 , \10309 , \9160 );
nand \U$9970 ( \10313 , \10311 , \10312 );
xor \U$9971 ( \10314 , \10307 , \10313 );
not \U$9972 ( \10315 , \9189 );
xor \U$9973 ( \10316 , \9197 , \9207 );
not \U$9974 ( \10317 , \10316 );
or \U$9975 ( \10318 , \10315 , \10317 );
or \U$9976 ( \10319 , \10316 , \9189 );
nand \U$9977 ( \10320 , \10318 , \10319 );
xor \U$9978 ( \10321 , \10314 , \10320 );
xor \U$9979 ( \10322 , \9283 , \9291 );
xor \U$9980 ( \10323 , \10322 , \9299 );
xor \U$9981 ( \10324 , \9256 , \9263 );
xor \U$9982 ( \10325 , \10324 , \9271 );
xor \U$9983 ( \10326 , \10323 , \10325 );
not \U$9984 ( \10327 , \9312 );
xor \U$9985 ( \10328 , \9321 , \9331 );
not \U$9986 ( \10329 , \10328 );
or \U$9987 ( \10330 , \10327 , \10329 );
or \U$9988 ( \10331 , \10328 , \9312 );
nand \U$9989 ( \10332 , \10330 , \10331 );
xor \U$9990 ( \10333 , \10326 , \10332 );
xor \U$9991 ( \10334 , \9373 , \9381 );
xor \U$9992 ( \10335 , \10334 , \9389 );
xor \U$9993 ( \10336 , \9345 , \9353 );
xor \U$9994 ( \10337 , \10336 , \9362 );
xor \U$9995 ( \10338 , \9394 , \10337 );
xor \U$9996 ( \10339 , \10335 , \10338 );
xor \U$9997 ( \10340 , \10333 , \10339 );
xor \U$9998 ( \10341 , \10321 , \10340 );
xor \U$9999 ( \10342 , \10270 , \10284 );
xor \U$10000 ( \10343 , \10342 , \10299 );
and \U$10001 ( \10344 , \10341 , \10343 );
and \U$10002 ( \10345 , \10259 , \10341 );
or \U$10003 ( \10346 , \10301 , \10344 , \10345 );
xor \U$10004 ( \10347 , \10249 , \10346 );
xor \U$10005 ( \10348 , \9916 , \9923 );
xor \U$10006 ( \10349 , \10348 , \9931 );
xor \U$10007 ( \10350 , \9942 , \9949 );
xor \U$10008 ( \10351 , \10350 , \9958 );
and \U$10009 ( \10352 , \10349 , \10351 );
xor \U$10010 ( \10353 , \9888 , \9896 );
xor \U$10011 ( \10354 , \10353 , \9905 );
xor \U$10012 ( \10355 , \9942 , \9949 );
xor \U$10013 ( \10356 , \10355 , \9958 );
and \U$10014 ( \10357 , \10354 , \10356 );
and \U$10015 ( \10358 , \10349 , \10354 );
or \U$10016 ( \10359 , \10352 , \10357 , \10358 );
xor \U$10017 ( \10360 , \9761 , \9763 );
xor \U$10018 ( \10361 , \10360 , \9771 );
xor \U$10019 ( \10362 , \9733 , \9741 );
xor \U$10020 ( \10363 , \10362 , \9750 );
xor \U$10021 ( \10364 , \10361 , \10363 );
xor \U$10022 ( \10365 , \9782 , \9789 );
xor \U$10023 ( \10366 , \10365 , \9798 );
and \U$10024 ( \10367 , \10364 , \10366 );
and \U$10025 ( \10368 , \10361 , \10363 );
or \U$10026 ( \10369 , \10367 , \10368 );
xor \U$10027 ( \10370 , \10359 , \10369 );
xor \U$10028 ( \10371 , \9811 , \9818 );
xor \U$10029 ( \10372 , \10371 , \9826 );
xor \U$10030 ( \10373 , \9836 , \9840 );
xor \U$10031 ( \10374 , \10373 , \9848 );
and \U$10032 ( \10375 , \10372 , \10374 );
xor \U$10033 ( \10376 , \9859 , \9866 );
xor \U$10034 ( \10377 , \10376 , \9874 );
xor \U$10035 ( \10378 , \9836 , \9840 );
xor \U$10036 ( \10379 , \10378 , \9848 );
and \U$10037 ( \10380 , \10377 , \10379 );
and \U$10038 ( \10381 , \10372 , \10377 );
or \U$10039 ( \10382 , \10375 , \10380 , \10381 );
and \U$10040 ( \10383 , \10370 , \10382 );
and \U$10041 ( \10384 , \10359 , \10369 );
or \U$10042 ( \10385 , \10383 , \10384 );
and \U$10043 ( \10386 , \5318 , RI986e620_21);
and \U$10044 ( \10387 , RI986f7f0_59, \5316 );
nor \U$10045 ( \10388 , \10386 , \10387 );
and \U$10046 ( \10389 , \10388 , \5052 );
not \U$10047 ( \10390 , \10388 );
and \U$10048 ( \10391 , \10390 , \5322 );
nor \U$10049 ( \10392 , \10389 , \10391 );
and \U$10050 ( \10393 , \5881 , RI986f700_57);
and \U$10051 ( \10394 , RI986f9d0_63, \5879 );
nor \U$10052 ( \10395 , \10393 , \10394 );
and \U$10053 ( \10396 , \10395 , \5594 );
not \U$10054 ( \10397 , \10395 );
and \U$10055 ( \10398 , \10397 , \5885 );
nor \U$10056 ( \10399 , \10396 , \10398 );
xor \U$10057 ( \10400 , \10392 , \10399 );
and \U$10058 ( \10401 , \6453 , RI986f8e0_61);
and \U$10059 ( \10402 , RI986f430_51, \6451 );
nor \U$10060 ( \10403 , \10401 , \10402 );
and \U$10061 ( \10404 , \10403 , \6190 );
not \U$10062 ( \10405 , \10403 );
and \U$10063 ( \10406 , \10405 , \6705 );
nor \U$10064 ( \10407 , \10404 , \10406 );
and \U$10065 ( \10408 , \10400 , \10407 );
and \U$10066 ( \10409 , \10392 , \10399 );
or \U$10067 ( \10410 , \10408 , \10409 );
and \U$10068 ( \10411 , \9237 , RI986dcc0_1);
and \U$10069 ( \10412 , RI986e170_11, \9235 );
nor \U$10070 ( \10413 , \10411 , \10412 );
and \U$10071 ( \10414 , \10413 , \9241 );
not \U$10072 ( \10415 , \10413 );
and \U$10073 ( \10416 , \10415 , \8836 );
nor \U$10074 ( \10417 , \10414 , \10416 );
and \U$10075 ( \10418 , RI9873030_179, RI9873120_181);
not \U$10076 ( \10419 , RI98730a8_180);
and \U$10077 ( \10420 , \10419 , RI9873120_181);
nor \U$10078 ( \10421 , \10419 , RI9873120_181);
or \U$10079 ( \10422 , \10420 , \10421 );
nor \U$10080 ( \10423 , RI9873030_179, RI9873120_181);
nor \U$10081 ( \10424 , \10418 , \10422 , \10423 );
nand \U$10082 ( \10425 , RI986e350_15, \10424 );
and \U$10083 ( \10426 , \10425 , \9840 );
not \U$10084 ( \10427 , \10425 );
not \U$10085 ( \10428 , \9840 );
and \U$10086 ( \10429 , \10427 , \10428 );
nor \U$10087 ( \10430 , \10426 , \10429 );
xor \U$10088 ( \10431 , \10417 , \10430 );
and \U$10089 ( \10432 , \9505 , RI986e080_9);
and \U$10090 ( \10433 , RI986e260_13, \9503 );
nor \U$10091 ( \10434 , \10432 , \10433 );
and \U$10092 ( \10435 , \10434 , \9510 );
not \U$10093 ( \10436 , \10434 );
and \U$10094 ( \10437 , \10436 , \9513 );
nor \U$10095 ( \10438 , \10435 , \10437 );
and \U$10096 ( \10439 , \10431 , \10438 );
and \U$10097 ( \10440 , \10417 , \10430 );
or \U$10098 ( \10441 , \10439 , \10440 );
xor \U$10099 ( \10442 , \10410 , \10441 );
and \U$10100 ( \10443 , \8486 , RI986dea0_5);
and \U$10101 ( \10444 , RI986ddb0_3, \8484 );
nor \U$10102 ( \10445 , \10443 , \10444 );
and \U$10103 ( \10446 , \10445 , \8050 );
not \U$10104 ( \10447 , \10445 );
and \U$10105 ( \10448 , \10447 , \8051 );
nor \U$10106 ( \10449 , \10446 , \10448 );
and \U$10107 ( \10450 , \7079 , RI986f340_49);
and \U$10108 ( \10451 , RI986f520_53, \7077 );
nor \U$10109 ( \10452 , \10450 , \10451 );
and \U$10110 ( \10453 , \10452 , \6710 );
not \U$10111 ( \10454 , \10452 );
and \U$10112 ( \10455 , \10454 , \6709 );
nor \U$10113 ( \10456 , \10453 , \10455 );
xor \U$10114 ( \10457 , \10449 , \10456 );
and \U$10115 ( \10458 , \7729 , RI986f610_55);
and \U$10116 ( \10459 , RI986df90_7, \7727 );
nor \U$10117 ( \10460 , \10458 , \10459 );
and \U$10118 ( \10461 , \10460 , \7480 );
not \U$10119 ( \10462 , \10460 );
and \U$10120 ( \10463 , \10462 , \7733 );
nor \U$10121 ( \10464 , \10461 , \10463 );
and \U$10122 ( \10465 , \10457 , \10464 );
and \U$10123 ( \10466 , \10449 , \10456 );
or \U$10124 ( \10467 , \10465 , \10466 );
and \U$10125 ( \10468 , \10442 , \10467 );
and \U$10126 ( \10469 , \10410 , \10441 );
or \U$10127 ( \10470 , \10468 , \10469 );
and \U$10128 ( \10471 , \376 , RI98709c0_97);
and \U$10129 ( \10472 , RI9870e70_107, \374 );
nor \U$10130 ( \10473 , \10471 , \10472 );
not \U$10131 ( \10474 , \10473 );
not \U$10132 ( \10475 , \367 );
and \U$10133 ( \10476 , \10474 , \10475 );
and \U$10134 ( \10477 , \10473 , \365 );
nor \U$10135 ( \10478 , \10476 , \10477 );
and \U$10136 ( \10479 , \395 , RI9870ab0_99);
and \U$10137 ( \10480 , RI9870d80_105, \393 );
nor \U$10138 ( \10481 , \10479 , \10480 );
not \U$10139 ( \10482 , \10481 );
not \U$10140 ( \10483 , \487 );
and \U$10141 ( \10484 , \10482 , \10483 );
and \U$10142 ( \10485 , \10481 , \386 );
nor \U$10143 ( \10486 , \10484 , \10485 );
or \U$10144 ( \10487 , \10478 , \10486 );
not \U$10145 ( \10488 , \10486 );
not \U$10146 ( \10489 , \10478 );
or \U$10147 ( \10490 , \10488 , \10489 );
not \U$10148 ( \10491 , \454 );
and \U$10149 ( \10492 , \465 , RI9870ba0_101);
and \U$10150 ( \10493 , RI9871050_111, \463 );
nor \U$10151 ( \10494 , \10492 , \10493 );
not \U$10152 ( \10495 , \10494 );
or \U$10153 ( \10496 , \10491 , \10495 );
or \U$10154 ( \10497 , \10494 , \454 );
nand \U$10155 ( \10498 , \10496 , \10497 );
nand \U$10156 ( \10499 , \10490 , \10498 );
nand \U$10157 ( \10500 , \10487 , \10499 );
and \U$10158 ( \10501 , \416 , RI986fe80_73);
and \U$10159 ( \10502 , RI9870060_77, \414 );
nor \U$10160 ( \10503 , \10501 , \10502 );
and \U$10161 ( \10504 , \10503 , \421 );
not \U$10162 ( \10505 , \10503 );
and \U$10163 ( \10506 , \10505 , \422 );
nor \U$10164 ( \10507 , \10504 , \10506 );
nand \U$10165 ( \10508 , RI986ff70_75, RI9871fc8_144);
or \U$10166 ( \10509 , \10507 , \10508 );
not \U$10167 ( \10510 , \10508 );
not \U$10168 ( \10511 , \10507 );
or \U$10169 ( \10512 , \10510 , \10511 );
not \U$10170 ( \10513 , \345 );
and \U$10171 ( \10514 , \354 , RI9870150_79);
and \U$10172 ( \10515 , RI9870f60_109, \352 );
nor \U$10173 ( \10516 , \10514 , \10515 );
not \U$10174 ( \10517 , \10516 );
or \U$10175 ( \10518 , \10513 , \10517 );
or \U$10176 ( \10519 , \10516 , \361 );
nand \U$10177 ( \10520 , \10518 , \10519 );
nand \U$10178 ( \10521 , \10512 , \10520 );
nand \U$10179 ( \10522 , \10509 , \10521 );
xor \U$10180 ( \10523 , \10500 , \10522 );
and \U$10181 ( \10524 , \776 , RI9871140_113);
and \U$10182 ( \10525 , RI9871320_117, \774 );
nor \U$10183 ( \10526 , \10524 , \10525 );
and \U$10184 ( \10527 , \10526 , \474 );
not \U$10185 ( \10528 , \10526 );
and \U$10186 ( \10529 , \10528 , \451 );
nor \U$10187 ( \10530 , \10527 , \10529 );
and \U$10188 ( \10531 , \438 , RI9870c90_103);
and \U$10189 ( \10532 , RI9871230_115, \436 );
nor \U$10190 ( \10533 , \10531 , \10532 );
and \U$10191 ( \10534 , \10533 , \444 );
not \U$10192 ( \10535 , \10533 );
and \U$10193 ( \10536 , \10535 , \443 );
nor \U$10194 ( \10537 , \10534 , \10536 );
xor \U$10195 ( \10538 , \10530 , \10537 );
not \U$10196 ( \10539 , \1301 );
and \U$10197 ( \10540 , \1293 , RI9871410_119);
and \U$10198 ( \10541 , RI98716e0_125, \1291 );
nor \U$10199 ( \10542 , \10540 , \10541 );
not \U$10200 ( \10543 , \10542 );
or \U$10201 ( \10544 , \10539 , \10543 );
or \U$10202 ( \10545 , \10542 , \1301 );
nand \U$10203 ( \10546 , \10544 , \10545 );
and \U$10204 ( \10547 , \10538 , \10546 );
and \U$10205 ( \10548 , \10530 , \10537 );
or \U$10206 ( \10549 , \10547 , \10548 );
and \U$10207 ( \10550 , \10523 , \10549 );
and \U$10208 ( \10551 , \10500 , \10522 );
or \U$10209 ( \10552 , \10550 , \10551 );
xor \U$10210 ( \10553 , \10470 , \10552 );
not \U$10211 ( \10554 , \3412 );
and \U$10212 ( \10555 , \3683 , RI986ef80_41);
and \U$10213 ( \10556 , RI986f250_47, \3681 );
nor \U$10214 ( \10557 , \10555 , \10556 );
not \U$10215 ( \10558 , \10557 );
or \U$10216 ( \10559 , \10554 , \10558 );
or \U$10217 ( \10560 , \10557 , \3918 );
nand \U$10218 ( \10561 , \10559 , \10560 );
and \U$10219 ( \10562 , \4203 , RI986f160_45);
and \U$10220 ( \10563 , RI986e530_19, \4201 );
nor \U$10221 ( \10564 , \10562 , \10563 );
and \U$10222 ( \10565 , \10564 , \4207 );
not \U$10223 ( \10566 , \10564 );
and \U$10224 ( \10567 , \10566 , \3923 );
nor \U$10225 ( \10568 , \10565 , \10567 );
xor \U$10226 ( \10569 , \10561 , \10568 );
not \U$10227 ( \10570 , \4521 );
and \U$10228 ( \10571 , \4710 , RI986e440_17);
and \U$10229 ( \10572 , RI986e710_23, \4708 );
nor \U$10230 ( \10573 , \10571 , \10572 );
not \U$10231 ( \10574 , \10573 );
or \U$10232 ( \10575 , \10570 , \10574 );
or \U$10233 ( \10576 , \10573 , \4519 );
nand \U$10234 ( \10577 , \10575 , \10576 );
and \U$10235 ( \10578 , \10569 , \10577 );
and \U$10236 ( \10579 , \10561 , \10568 );
or \U$10237 ( \10580 , \10578 , \10579 );
and \U$10238 ( \10581 , \2464 , RI986eda0_37);
and \U$10239 ( \10582 , RI986ebc0_33, \2462 );
nor \U$10240 ( \10583 , \10581 , \10582 );
and \U$10241 ( \10584 , \10583 , \2468 );
not \U$10242 ( \10585 , \10583 );
and \U$10243 ( \10586 , \10585 , \2263 );
nor \U$10244 ( \10587 , \10584 , \10586 );
and \U$10245 ( \10588 , \2274 , RI986e800_25);
and \U$10246 ( \10589 , RI986ee90_39, \2272 );
nor \U$10247 ( \10590 , \10588 , \10589 );
and \U$10248 ( \10591 , \10590 , \2030 );
not \U$10249 ( \10592 , \10590 );
and \U$10250 ( \10593 , \10592 , \2031 );
nor \U$10251 ( \10594 , \10591 , \10593 );
xor \U$10252 ( \10595 , \10587 , \10594 );
not \U$10253 ( \10596 , \2935 );
and \U$10254 ( \10597 , \3254 , RI986ecb0_35);
and \U$10255 ( \10598 , RI986f070_43, \3252 );
nor \U$10256 ( \10599 , \10597 , \10598 );
not \U$10257 ( \10600 , \10599 );
or \U$10258 ( \10601 , \10596 , \10600 );
or \U$10259 ( \10602 , \10599 , \2935 );
nand \U$10260 ( \10603 , \10601 , \10602 );
and \U$10261 ( \10604 , \10595 , \10603 );
and \U$10262 ( \10605 , \10587 , \10594 );
or \U$10263 ( \10606 , \10604 , \10605 );
xor \U$10264 ( \10607 , \10580 , \10606 );
and \U$10265 ( \10608 , \1311 , RI98715f0_123);
and \U$10266 ( \10609 , RI986ead0_31, \1309 );
nor \U$10267 ( \10610 , \10608 , \10609 );
and \U$10268 ( \10611 , \10610 , \1458 );
not \U$10269 ( \10612 , \10610 );
and \U$10270 ( \10613 , \10612 , \1318 );
nor \U$10271 ( \10614 , \10611 , \10613 );
and \U$10272 ( \10615 , \1329 , RI98717d0_127);
and \U$10273 ( \10616 , RI9871500_121, \1327 );
nor \U$10274 ( \10617 , \10615 , \10616 );
and \U$10275 ( \10618 , \10617 , \1336 );
not \U$10276 ( \10619 , \10617 );
and \U$10277 ( \10620 , \10619 , \1337 );
nor \U$10278 ( \10621 , \10618 , \10620 );
xor \U$10279 ( \10622 , \10614 , \10621 );
not \U$10280 ( \10623 , \2034 );
and \U$10281 ( \10624 , \2042 , RI986e9e0_29);
and \U$10282 ( \10625 , RI986e8f0_27, \2040 );
nor \U$10283 ( \10626 , \10624 , \10625 );
not \U$10284 ( \10627 , \10626 );
or \U$10285 ( \10628 , \10623 , \10627 );
or \U$10286 ( \10629 , \10626 , \2034 );
nand \U$10287 ( \10630 , \10628 , \10629 );
and \U$10288 ( \10631 , \10622 , \10630 );
and \U$10289 ( \10632 , \10614 , \10621 );
or \U$10290 ( \10633 , \10631 , \10632 );
and \U$10291 ( \10634 , \10607 , \10633 );
and \U$10292 ( \10635 , \10580 , \10606 );
or \U$10293 ( \10636 , \10634 , \10635 );
and \U$10294 ( \10637 , \10553 , \10636 );
and \U$10295 ( \10638 , \10470 , \10552 );
or \U$10296 ( \10639 , \10637 , \10638 );
xor \U$10297 ( \10640 , \10385 , \10639 );
xor \U$10298 ( \10641 , \9531 , \9538 );
xor \U$10299 ( \10642 , \10641 , \9546 );
xor \U$10300 ( \10643 , \9524 , \9572 );
xor \U$10301 ( \10644 , \10642 , \10643 );
xor \U$10302 ( \10645 , \9601 , \9612 );
xor \U$10303 ( \10646 , \10645 , \9639 );
and \U$10304 ( \10647 , \10644 , \10646 );
xor \U$10305 ( \10648 , \9674 , \9682 );
xor \U$10306 ( \10649 , \10648 , \9690 );
xor \U$10307 ( \10650 , \9667 , \9717 );
xor \U$10308 ( \10651 , \10649 , \10650 );
xor \U$10309 ( \10652 , \9601 , \9612 );
xor \U$10310 ( \10653 , \10652 , \9639 );
and \U$10311 ( \10654 , \10651 , \10653 );
and \U$10312 ( \10655 , \10644 , \10651 );
or \U$10313 ( \10656 , \10647 , \10654 , \10655 );
and \U$10314 ( \10657 , \10640 , \10656 );
and \U$10315 ( \10658 , \10385 , \10639 );
or \U$10316 ( \10659 , \10657 , \10658 );
xor \U$10317 ( \10660 , \9804 , \9880 );
xor \U$10318 ( \10661 , \10660 , \9964 );
xor \U$10319 ( \10662 , \9577 , \9642 );
xor \U$10320 ( \10663 , \10662 , \9722 );
and \U$10321 ( \10664 , \10661 , \10663 );
xor \U$10322 ( \10665 , \10659 , \10664 );
xor \U$10323 ( \10666 , \9829 , \9851 );
xor \U$10324 ( \10667 , \10666 , \9877 );
xor \U$10325 ( \10668 , \9908 , \9934 );
xor \U$10326 ( \10669 , \10668 , \9961 );
xor \U$10327 ( \10670 , \10667 , \10669 );
xor \U$10328 ( \10671 , \9753 , \9774 );
xor \U$10329 ( \10672 , \10671 , \9801 );
and \U$10330 ( \10673 , \10670 , \10672 );
and \U$10331 ( \10674 , \10667 , \10669 );
or \U$10332 ( \10675 , \10673 , \10674 );
xor \U$10333 ( \10676 , \10251 , \10253 );
xor \U$10334 ( \10677 , \10676 , \10256 );
and \U$10335 ( \10678 , \10675 , \10677 );
xor \U$10336 ( \10679 , \10046 , \10070 );
xor \U$10337 ( \10680 , \10679 , \10094 );
xor \U$10338 ( \10681 , \10030 , \10171 );
xor \U$10339 ( \10682 , \10680 , \10681 );
xor \U$10340 ( \10683 , \10251 , \10253 );
xor \U$10341 ( \10684 , \10683 , \10256 );
and \U$10342 ( \10685 , \10682 , \10684 );
and \U$10343 ( \10686 , \10675 , \10682 );
or \U$10344 ( \10687 , \10678 , \10685 , \10686 );
and \U$10345 ( \10688 , \10665 , \10687 );
and \U$10346 ( \10689 , \10659 , \10664 );
or \U$10347 ( \10690 , \10688 , \10689 );
xor \U$10348 ( \10691 , \10225 , \10247 );
xor \U$10349 ( \10692 , \9725 , \9967 );
xor \U$10350 ( \10693 , \10692 , \10176 );
and \U$10351 ( \10694 , \10691 , \10693 );
xor \U$10352 ( \10695 , \10270 , \10284 );
xor \U$10353 ( \10696 , \10695 , \10299 );
xor \U$10354 ( \10697 , \10259 , \10341 );
xor \U$10355 ( \10698 , \10696 , \10697 );
xor \U$10356 ( \10699 , \9725 , \9967 );
xor \U$10357 ( \10700 , \10699 , \10176 );
and \U$10358 ( \10701 , \10698 , \10700 );
and \U$10359 ( \10702 , \10691 , \10698 );
or \U$10360 ( \10703 , \10694 , \10701 , \10702 );
xor \U$10361 ( \10704 , \10690 , \10703 );
xor \U$10362 ( \10705 , \10229 , \10237 );
and \U$10363 ( \10706 , \10705 , \10246 );
and \U$10364 ( \10707 , \10229 , \10237 );
or \U$10365 ( \10708 , \10706 , \10707 );
xor \U$10366 ( \10709 , \10195 , \10207 );
and \U$10367 ( \10710 , \10709 , \10224 );
and \U$10368 ( \10711 , \10195 , \10207 );
or \U$10369 ( \10712 , \10710 , \10711 );
xor \U$10370 ( \10713 , \10708 , \10712 );
xor \U$10371 ( \10714 , \10307 , \10313 );
xor \U$10372 ( \10715 , \10714 , \10320 );
and \U$10373 ( \10716 , \10333 , \10715 );
xor \U$10374 ( \10717 , \10307 , \10313 );
xor \U$10375 ( \10718 , \10717 , \10320 );
and \U$10376 ( \10719 , \10339 , \10718 );
and \U$10377 ( \10720 , \10333 , \10339 );
or \U$10378 ( \10721 , \10716 , \10719 , \10720 );
xor \U$10379 ( \10722 , \10713 , \10721 );
xor \U$10380 ( \10723 , \10289 , \10293 );
and \U$10381 ( \10724 , \10723 , \10298 );
and \U$10382 ( \10725 , \10289 , \10293 );
or \U$10383 ( \10726 , \10724 , \10725 );
xor \U$10384 ( \10727 , \10263 , \10264 );
and \U$10385 ( \10728 , \10727 , \10269 );
and \U$10386 ( \10729 , \10263 , \10264 );
or \U$10387 ( \10730 , \10728 , \10729 );
xor \U$10388 ( \10731 , \10726 , \10730 );
xor \U$10389 ( \10732 , \10274 , \10278 );
and \U$10390 ( \10733 , \10732 , \10283 );
and \U$10391 ( \10734 , \10274 , \10278 );
or \U$10392 ( \10735 , \10733 , \10734 );
xor \U$10393 ( \10736 , \10731 , \10735 );
xor \U$10394 ( \10737 , \10307 , \10313 );
and \U$10395 ( \10738 , \10737 , \10320 );
and \U$10396 ( \10739 , \10307 , \10313 );
or \U$10397 ( \10740 , \10738 , \10739 );
xor \U$10398 ( \10741 , \9373 , \9381 );
xor \U$10399 ( \10742 , \10741 , \9389 );
and \U$10400 ( \10743 , \9394 , \10742 );
xor \U$10401 ( \10744 , \9373 , \9381 );
xor \U$10402 ( \10745 , \10744 , \9389 );
and \U$10403 ( \10746 , \10337 , \10745 );
and \U$10404 ( \10747 , \9394 , \10337 );
or \U$10405 ( \10748 , \10743 , \10746 , \10747 );
xor \U$10406 ( \10749 , \10740 , \10748 );
xor \U$10407 ( \10750 , \10323 , \10325 );
and \U$10408 ( \10751 , \10750 , \10332 );
and \U$10409 ( \10752 , \10323 , \10325 );
or \U$10410 ( \10753 , \10751 , \10752 );
xor \U$10411 ( \10754 , \10749 , \10753 );
xor \U$10412 ( \10755 , \10736 , \10754 );
not \U$10413 ( \10756 , \9181 );
xor \U$10414 ( \10757 , \9245 , \9209 );
not \U$10415 ( \10758 , \10757 );
or \U$10416 ( \10759 , \10756 , \10758 );
or \U$10417 ( \10760 , \10757 , \9181 );
nand \U$10418 ( \10761 , \10759 , \10760 );
not \U$10419 ( \10762 , \9274 );
xor \U$10420 ( \10763 , \9333 , \9302 );
not \U$10421 ( \10764 , \10763 );
or \U$10422 ( \10765 , \10762 , \10764 );
or \U$10423 ( \10766 , \10763 , \9274 );
nand \U$10424 ( \10767 , \10765 , \10766 );
xor \U$10425 ( \10768 , \10761 , \10767 );
xor \U$10426 ( \10769 , \9365 , \9392 );
not \U$10427 ( \10770 , \9394 );
xor \U$10428 ( \10771 , \10769 , \10770 );
xor \U$10429 ( \10772 , \10768 , \10771 );
xor \U$10430 ( \10773 , \10270 , \10284 );
and \U$10431 ( \10774 , \10773 , \10299 );
and \U$10432 ( \10775 , \10270 , \10284 );
or \U$10433 ( \10776 , \10774 , \10775 );
not \U$10434 ( \10777 , \9112 );
xor \U$10435 ( \10778 , \9114 , \9127 );
not \U$10436 ( \10779 , \10778 );
or \U$10437 ( \10780 , \10777 , \10779 );
or \U$10438 ( \10781 , \10778 , \9112 );
nand \U$10439 ( \10782 , \10780 , \10781 );
not \U$10440 ( \10783 , \9094 );
xor \U$10441 ( \10784 , \9091 , \9099 );
not \U$10442 ( \10785 , \10784 );
or \U$10443 ( \10786 , \10783 , \10785 );
or \U$10444 ( \10787 , \10784 , \9094 );
nand \U$10445 ( \10788 , \10786 , \10787 );
xor \U$10446 ( \10789 , \10782 , \10788 );
xor \U$10447 ( \10790 , \9134 , \9140 );
xor \U$10448 ( \10791 , \10790 , \9147 );
xor \U$10449 ( \10792 , \10789 , \10791 );
xor \U$10450 ( \10793 , \10776 , \10792 );
xor \U$10451 ( \10794 , \10772 , \10793 );
xor \U$10452 ( \10795 , \10755 , \10794 );
xor \U$10453 ( \10796 , \10722 , \10795 );
xor \U$10454 ( \10797 , \10704 , \10796 );
and \U$10455 ( \10798 , \10347 , \10797 );
xor \U$10456 ( \10799 , \10392 , \10399 );
xor \U$10457 ( \10800 , \10799 , \10407 );
xor \U$10458 ( \10801 , \10561 , \10568 );
xor \U$10459 ( \10802 , \10801 , \10577 );
xor \U$10460 ( \10803 , \10800 , \10802 );
xor \U$10461 ( \10804 , \10449 , \10456 );
xor \U$10462 ( \10805 , \10804 , \10464 );
and \U$10463 ( \10806 , \10803 , \10805 );
and \U$10464 ( \10807 , \10800 , \10802 );
or \U$10465 ( \10808 , \10806 , \10807 );
not \U$10466 ( \10809 , \10507 );
not \U$10467 ( \10810 , \10520 );
or \U$10468 ( \10811 , \10809 , \10810 );
or \U$10469 ( \10812 , \10507 , \10520 );
nand \U$10470 ( \10813 , \10811 , \10812 );
not \U$10471 ( \10814 , \10813 );
not \U$10472 ( \10815 , \10508 );
and \U$10473 ( \10816 , \10814 , \10815 );
and \U$10474 ( \10817 , \10813 , \10508 );
nor \U$10475 ( \10818 , \10816 , \10817 );
not \U$10476 ( \10819 , \10478 );
not \U$10477 ( \10820 , \10498 );
or \U$10478 ( \10821 , \10819 , \10820 );
or \U$10479 ( \10822 , \10478 , \10498 );
nand \U$10480 ( \10823 , \10821 , \10822 );
not \U$10481 ( \10824 , \10823 );
not \U$10482 ( \10825 , \10486 );
and \U$10483 ( \10826 , \10824 , \10825 );
and \U$10484 ( \10827 , \10823 , \10486 );
nor \U$10485 ( \10828 , \10826 , \10827 );
nand \U$10486 ( \10829 , \10818 , \10828 );
xor \U$10487 ( \10830 , \10808 , \10829 );
xor \U$10488 ( \10831 , \10530 , \10537 );
xor \U$10489 ( \10832 , \10831 , \10546 );
xor \U$10490 ( \10833 , \10587 , \10594 );
xor \U$10491 ( \10834 , \10833 , \10603 );
and \U$10492 ( \10835 , \10832 , \10834 );
xor \U$10493 ( \10836 , \10614 , \10621 );
xor \U$10494 ( \10837 , \10836 , \10630 );
xor \U$10495 ( \10838 , \10587 , \10594 );
xor \U$10496 ( \10839 , \10838 , \10603 );
and \U$10497 ( \10840 , \10837 , \10839 );
and \U$10498 ( \10841 , \10832 , \10837 );
or \U$10499 ( \10842 , \10835 , \10840 , \10841 );
and \U$10500 ( \10843 , \10830 , \10842 );
and \U$10501 ( \10844 , \10808 , \10829 );
or \U$10502 ( \10845 , \10843 , \10844 );
not \U$10503 ( \10846 , \454 );
and \U$10504 ( \10847 , \465 , RI9870e70_107);
and \U$10505 ( \10848 , RI9870ba0_101, \463 );
nor \U$10506 ( \10849 , \10847 , \10848 );
not \U$10507 ( \10850 , \10849 );
or \U$10508 ( \10851 , \10846 , \10850 );
or \U$10509 ( \10852 , \10849 , \454 );
nand \U$10510 ( \10853 , \10851 , \10852 );
and \U$10511 ( \10854 , \438 , RI9871050_111);
and \U$10512 ( \10855 , RI9870c90_103, \436 );
nor \U$10513 ( \10856 , \10854 , \10855 );
and \U$10514 ( \10857 , \10856 , \444 );
not \U$10515 ( \10858 , \10856 );
and \U$10516 ( \10859 , \10858 , \443 );
nor \U$10517 ( \10860 , \10857 , \10859 );
xor \U$10518 ( \10861 , \10853 , \10860 );
not \U$10519 ( \10862 , \365 );
and \U$10520 ( \10863 , \376 , RI9870d80_105);
and \U$10521 ( \10864 , RI98709c0_97, \374 );
nor \U$10522 ( \10865 , \10863 , \10864 );
not \U$10523 ( \10866 , \10865 );
or \U$10524 ( \10867 , \10862 , \10866 );
or \U$10525 ( \10868 , \10865 , \365 );
nand \U$10526 ( \10869 , \10867 , \10868 );
and \U$10527 ( \10870 , \10861 , \10869 );
and \U$10528 ( \10871 , \10853 , \10860 );
or \U$10529 ( \10872 , \10870 , \10871 );
and \U$10530 ( \10873 , \416 , RI986ff70_75);
and \U$10531 ( \10874 , RI986fe80_73, \414 );
nor \U$10532 ( \10875 , \10873 , \10874 );
and \U$10533 ( \10876 , \10875 , \422 );
not \U$10534 ( \10877 , \10875 );
and \U$10535 ( \10878 , \10877 , \421 );
nor \U$10536 ( \10879 , \10876 , \10878 );
not \U$10537 ( \10880 , \386 );
and \U$10538 ( \10881 , \395 , RI9870f60_109);
and \U$10539 ( \10882 , RI9870ab0_99, \393 );
nor \U$10540 ( \10883 , \10881 , \10882 );
not \U$10541 ( \10884 , \10883 );
or \U$10542 ( \10885 , \10880 , \10884 );
or \U$10543 ( \10886 , \10883 , \487 );
nand \U$10544 ( \10887 , \10885 , \10886 );
xor \U$10545 ( \10888 , \10879 , \10887 );
not \U$10546 ( \10889 , \345 );
and \U$10547 ( \10890 , \354 , RI9870060_77);
and \U$10548 ( \10891 , RI9870150_79, \352 );
nor \U$10549 ( \10892 , \10890 , \10891 );
not \U$10550 ( \10893 , \10892 );
or \U$10551 ( \10894 , \10889 , \10893 );
or \U$10552 ( \10895 , \10892 , \345 );
nand \U$10553 ( \10896 , \10894 , \10895 );
and \U$10554 ( \10897 , \10888 , \10896 );
and \U$10555 ( \10898 , \10879 , \10887 );
or \U$10556 ( \10899 , \10897 , \10898 );
xor \U$10557 ( \10900 , \10872 , \10899 );
not \U$10558 ( \10901 , \1128 );
and \U$10559 ( \10902 , \1293 , RI9871320_117);
and \U$10560 ( \10903 , RI9871410_119, \1291 );
nor \U$10561 ( \10904 , \10902 , \10903 );
not \U$10562 ( \10905 , \10904 );
or \U$10563 ( \10906 , \10901 , \10905 );
or \U$10564 ( \10907 , \10904 , \1301 );
nand \U$10565 ( \10908 , \10906 , \10907 );
and \U$10566 ( \10909 , \776 , RI9871230_115);
and \U$10567 ( \10910 , RI9871140_113, \774 );
nor \U$10568 ( \10911 , \10909 , \10910 );
and \U$10569 ( \10912 , \10911 , \474 );
not \U$10570 ( \10913 , \10911 );
and \U$10571 ( \10914 , \10913 , \451 );
nor \U$10572 ( \10915 , \10912 , \10914 );
xor \U$10573 ( \10916 , \10908 , \10915 );
and \U$10574 ( \10917 , \1329 , RI98716e0_125);
and \U$10575 ( \10918 , RI98717d0_127, \1327 );
nor \U$10576 ( \10919 , \10917 , \10918 );
and \U$10577 ( \10920 , \10919 , \1336 );
not \U$10578 ( \10921 , \10919 );
and \U$10579 ( \10922 , \10921 , \1337 );
nor \U$10580 ( \10923 , \10920 , \10922 );
and \U$10581 ( \10924 , \10916 , \10923 );
and \U$10582 ( \10925 , \10908 , \10915 );
or \U$10583 ( \10926 , \10924 , \10925 );
and \U$10584 ( \10927 , \10900 , \10926 );
and \U$10585 ( \10928 , \10872 , \10899 );
or \U$10586 ( \10929 , \10927 , \10928 );
and \U$10587 ( \10930 , \7729 , RI986f520_53);
and \U$10588 ( \10931 , RI986f610_55, \7727 );
nor \U$10589 ( \10932 , \10930 , \10931 );
and \U$10590 ( \10933 , \10932 , \7480 );
not \U$10591 ( \10934 , \10932 );
and \U$10592 ( \10935 , \10934 , \7733 );
nor \U$10593 ( \10936 , \10933 , \10935 );
and \U$10594 ( \10937 , \8486 , RI986df90_7);
and \U$10595 ( \10938 , RI986dea0_5, \8484 );
nor \U$10596 ( \10939 , \10937 , \10938 );
and \U$10597 ( \10940 , \10939 , \8050 );
not \U$10598 ( \10941 , \10939 );
and \U$10599 ( \10942 , \10941 , \8051 );
nor \U$10600 ( \10943 , \10940 , \10942 );
xor \U$10601 ( \10944 , \10936 , \10943 );
and \U$10602 ( \10945 , \9237 , RI986ddb0_3);
and \U$10603 ( \10946 , RI986dcc0_1, \9235 );
nor \U$10604 ( \10947 , \10945 , \10946 );
and \U$10605 ( \10948 , \10947 , \9241 );
not \U$10606 ( \10949 , \10947 );
and \U$10607 ( \10950 , \10949 , \8836 );
nor \U$10608 ( \10951 , \10948 , \10950 );
and \U$10609 ( \10952 , \10944 , \10951 );
and \U$10610 ( \10953 , \10936 , \10943 );
or \U$10611 ( \10954 , \10952 , \10953 );
and \U$10612 ( \10955 , \9505 , RI986e170_11);
and \U$10613 ( \10956 , RI986e080_9, \9503 );
nor \U$10614 ( \10957 , \10955 , \10956 );
and \U$10615 ( \10958 , \10957 , \9510 );
not \U$10616 ( \10959 , \10957 );
and \U$10617 ( \10960 , \10959 , \9513 );
nor \U$10618 ( \10961 , \10958 , \10960 );
not \U$10619 ( \10962 , RI9873210_183);
not \U$10620 ( \10963 , RI9873198_182);
or \U$10621 ( \10964 , \10962 , \10963 );
nand \U$10622 ( \10965 , \10964 , RI98730a8_180);
xor \U$10623 ( \10966 , \10961 , \10965 );
and \U$10624 ( \10967 , \10424 , RI986e260_13);
and \U$10625 ( \10968 , RI986e350_15, \10422 );
nor \U$10626 ( \10969 , \10967 , \10968 );
and \U$10627 ( \10970 , \10969 , \9840 );
not \U$10628 ( \10971 , \10969 );
and \U$10629 ( \10972 , \10971 , \10428 );
nor \U$10630 ( \10973 , \10970 , \10972 );
and \U$10631 ( \10974 , \10966 , \10973 );
and \U$10632 ( \10975 , \10961 , \10965 );
or \U$10633 ( \10976 , \10974 , \10975 );
xor \U$10634 ( \10977 , \10954 , \10976 );
and \U$10635 ( \10978 , \7079 , RI986f430_51);
and \U$10636 ( \10979 , RI986f340_49, \7077 );
nor \U$10637 ( \10980 , \10978 , \10979 );
and \U$10638 ( \10981 , \10980 , \6710 );
not \U$10639 ( \10982 , \10980 );
and \U$10640 ( \10983 , \10982 , \6709 );
nor \U$10641 ( \10984 , \10981 , \10983 );
and \U$10642 ( \10985 , \5881 , RI986f7f0_59);
and \U$10643 ( \10986 , RI986f700_57, \5879 );
nor \U$10644 ( \10987 , \10985 , \10986 );
and \U$10645 ( \10988 , \10987 , \5594 );
not \U$10646 ( \10989 , \10987 );
and \U$10647 ( \10990 , \10989 , \5885 );
nor \U$10648 ( \10991 , \10988 , \10990 );
xor \U$10649 ( \10992 , \10984 , \10991 );
and \U$10650 ( \10993 , \6453 , RI986f9d0_63);
and \U$10651 ( \10994 , RI986f8e0_61, \6451 );
nor \U$10652 ( \10995 , \10993 , \10994 );
and \U$10653 ( \10996 , \10995 , \6190 );
not \U$10654 ( \10997 , \10995 );
and \U$10655 ( \10998 , \10997 , \6705 );
nor \U$10656 ( \10999 , \10996 , \10998 );
and \U$10657 ( \11000 , \10992 , \10999 );
and \U$10658 ( \11001 , \10984 , \10991 );
or \U$10659 ( \11002 , \11000 , \11001 );
and \U$10660 ( \11003 , \10977 , \11002 );
and \U$10661 ( \11004 , \10954 , \10976 );
or \U$10662 ( \11005 , \11003 , \11004 );
xor \U$10663 ( \11006 , \10929 , \11005 );
and \U$10664 ( \11007 , \4203 , RI986f250_47);
and \U$10665 ( \11008 , RI986f160_45, \4201 );
nor \U$10666 ( \11009 , \11007 , \11008 );
and \U$10667 ( \11010 , \11009 , \4207 );
not \U$10668 ( \11011 , \11009 );
and \U$10669 ( \11012 , \11011 , \3922 );
nor \U$10670 ( \11013 , \11010 , \11012 );
not \U$10671 ( \11014 , \4521 );
and \U$10672 ( \11015 , \4710 , RI986e530_19);
and \U$10673 ( \11016 , RI986e440_17, \4708 );
nor \U$10674 ( \11017 , \11015 , \11016 );
not \U$10675 ( \11018 , \11017 );
or \U$10676 ( \11019 , \11014 , \11018 );
or \U$10677 ( \11020 , \11017 , \4519 );
nand \U$10678 ( \11021 , \11019 , \11020 );
xor \U$10679 ( \11022 , \11013 , \11021 );
and \U$10680 ( \11023 , \5318 , RI986e710_23);
and \U$10681 ( \11024 , RI986e620_21, \5316 );
nor \U$10682 ( \11025 , \11023 , \11024 );
and \U$10683 ( \11026 , \11025 , \5052 );
not \U$10684 ( \11027 , \11025 );
and \U$10685 ( \11028 , \11027 , \5322 );
nor \U$10686 ( \11029 , \11026 , \11028 );
and \U$10687 ( \11030 , \11022 , \11029 );
and \U$10688 ( \11031 , \11013 , \11021 );
or \U$10689 ( \11032 , \11030 , \11031 );
not \U$10690 ( \11033 , \2935 );
and \U$10691 ( \11034 , \3254 , RI986ebc0_33);
and \U$10692 ( \11035 , RI986ecb0_35, \3252 );
nor \U$10693 ( \11036 , \11034 , \11035 );
not \U$10694 ( \11037 , \11036 );
or \U$10695 ( \11038 , \11033 , \11037 );
or \U$10696 ( \11039 , \11036 , \3406 );
nand \U$10697 ( \11040 , \11038 , \11039 );
and \U$10698 ( \11041 , \2464 , RI986ee90_39);
and \U$10699 ( \11042 , RI986eda0_37, \2462 );
nor \U$10700 ( \11043 , \11041 , \11042 );
and \U$10701 ( \11044 , \11043 , \2468 );
not \U$10702 ( \11045 , \11043 );
and \U$10703 ( \11046 , \11045 , \2263 );
nor \U$10704 ( \11047 , \11044 , \11046 );
xor \U$10705 ( \11048 , \11040 , \11047 );
not \U$10706 ( \11049 , \3412 );
and \U$10707 ( \11050 , \3683 , RI986f070_43);
and \U$10708 ( \11051 , RI986ef80_41, \3681 );
nor \U$10709 ( \11052 , \11050 , \11051 );
not \U$10710 ( \11053 , \11052 );
or \U$10711 ( \11054 , \11049 , \11053 );
or \U$10712 ( \11055 , \11052 , \3918 );
nand \U$10713 ( \11056 , \11054 , \11055 );
and \U$10714 ( \11057 , \11048 , \11056 );
and \U$10715 ( \11058 , \11040 , \11047 );
or \U$10716 ( \11059 , \11057 , \11058 );
xor \U$10717 ( \11060 , \11032 , \11059 );
and \U$10718 ( \11061 , \1311 , RI9871500_121);
and \U$10719 ( \11062 , RI98715f0_123, \1309 );
nor \U$10720 ( \11063 , \11061 , \11062 );
and \U$10721 ( \11064 , \11063 , \1458 );
not \U$10722 ( \11065 , \11063 );
and \U$10723 ( \11066 , \11065 , \1318 );
nor \U$10724 ( \11067 , \11064 , \11066 );
not \U$10725 ( \11068 , \2034 );
and \U$10726 ( \11069 , \2042 , RI986ead0_31);
and \U$10727 ( \11070 , RI986e9e0_29, \2040 );
nor \U$10728 ( \11071 , \11069 , \11070 );
not \U$10729 ( \11072 , \11071 );
or \U$10730 ( \11073 , \11068 , \11072 );
or \U$10731 ( \11074 , \11071 , \1462 );
nand \U$10732 ( \11075 , \11073 , \11074 );
xor \U$10733 ( \11076 , \11067 , \11075 );
and \U$10734 ( \11077 , \2274 , RI986e8f0_27);
and \U$10735 ( \11078 , RI986e800_25, \2272 );
nor \U$10736 ( \11079 , \11077 , \11078 );
and \U$10737 ( \11080 , \11079 , \2030 );
not \U$10738 ( \11081 , \11079 );
and \U$10739 ( \11082 , \11081 , \2031 );
nor \U$10740 ( \11083 , \11080 , \11082 );
and \U$10741 ( \11084 , \11076 , \11083 );
and \U$10742 ( \11085 , \11067 , \11075 );
or \U$10743 ( \11086 , \11084 , \11085 );
and \U$10744 ( \11087 , \11060 , \11086 );
and \U$10745 ( \11088 , \11032 , \11059 );
or \U$10746 ( \11089 , \11087 , \11088 );
and \U$10747 ( \11090 , \11006 , \11089 );
and \U$10748 ( \11091 , \10929 , \11005 );
or \U$10749 ( \11092 , \11090 , \11091 );
xor \U$10750 ( \11093 , \10845 , \11092 );
xor \U$10751 ( \11094 , \9836 , \9840 );
xor \U$10752 ( \11095 , \11094 , \9848 );
xor \U$10753 ( \11096 , \10372 , \10377 );
xor \U$10754 ( \11097 , \11095 , \11096 );
xor \U$10755 ( \11098 , \10361 , \10363 );
xor \U$10756 ( \11099 , \11098 , \10366 );
and \U$10757 ( \11100 , \11097 , \11099 );
xor \U$10758 ( \11101 , \9942 , \9949 );
xor \U$10759 ( \11102 , \11101 , \9958 );
xor \U$10760 ( \11103 , \10349 , \10354 );
xor \U$10761 ( \11104 , \11102 , \11103 );
xor \U$10762 ( \11105 , \10361 , \10363 );
xor \U$10763 ( \11106 , \11105 , \10366 );
and \U$10764 ( \11107 , \11104 , \11106 );
and \U$10765 ( \11108 , \11097 , \11104 );
or \U$10766 ( \11109 , \11100 , \11107 , \11108 );
and \U$10767 ( \11110 , \11093 , \11109 );
and \U$10768 ( \11111 , \10845 , \11092 );
or \U$10769 ( \11112 , \11110 , \11111 );
xor \U$10770 ( \11113 , \10470 , \10552 );
xor \U$10771 ( \11114 , \11113 , \10636 );
xor \U$10772 ( \11115 , \10359 , \10369 );
xor \U$10773 ( \11116 , \11115 , \10382 );
and \U$10774 ( \11117 , \11114 , \11116 );
xor \U$10775 ( \11118 , \11112 , \11117 );
xor \U$10776 ( \11119 , \10410 , \10441 );
xor \U$10777 ( \11120 , \11119 , \10467 );
xor \U$10778 ( \11121 , \10580 , \10606 );
xor \U$10779 ( \11122 , \11121 , \10633 );
xor \U$10780 ( \11123 , \11120 , \11122 );
xor \U$10781 ( \11124 , \10500 , \10522 );
xor \U$10782 ( \11125 , \11124 , \10549 );
and \U$10783 ( \11126 , \11123 , \11125 );
and \U$10784 ( \11127 , \11120 , \11122 );
or \U$10785 ( \11128 , \11126 , \11127 );
xor \U$10786 ( \11129 , \10667 , \10669 );
xor \U$10787 ( \11130 , \11129 , \10672 );
and \U$10788 ( \11131 , \11128 , \11130 );
xor \U$10789 ( \11132 , \9601 , \9612 );
xor \U$10790 ( \11133 , \11132 , \9639 );
xor \U$10791 ( \11134 , \10644 , \10651 );
xor \U$10792 ( \11135 , \11133 , \11134 );
xor \U$10793 ( \11136 , \10667 , \10669 );
xor \U$10794 ( \11137 , \11136 , \10672 );
and \U$10795 ( \11138 , \11135 , \11137 );
and \U$10796 ( \11139 , \11128 , \11135 );
or \U$10797 ( \11140 , \11131 , \11138 , \11139 );
and \U$10798 ( \11141 , \11118 , \11140 );
and \U$10799 ( \11142 , \11112 , \11117 );
or \U$10800 ( \11143 , \11141 , \11142 );
xor \U$10801 ( \11144 , \10661 , \10663 );
xor \U$10802 ( \11145 , \10385 , \10639 );
xor \U$10803 ( \11146 , \11145 , \10656 );
and \U$10804 ( \11147 , \11144 , \11146 );
xor \U$10805 ( \11148 , \10251 , \10253 );
xor \U$10806 ( \11149 , \11148 , \10256 );
xor \U$10807 ( \11150 , \10675 , \10682 );
xor \U$10808 ( \11151 , \11149 , \11150 );
xor \U$10809 ( \11152 , \10385 , \10639 );
xor \U$10810 ( \11153 , \11152 , \10656 );
and \U$10811 ( \11154 , \11151 , \11153 );
and \U$10812 ( \11155 , \11144 , \11151 );
or \U$10813 ( \11156 , \11147 , \11154 , \11155 );
xor \U$10814 ( \11157 , \11143 , \11156 );
xor \U$10815 ( \11158 , \9725 , \9967 );
xor \U$10816 ( \11159 , \11158 , \10176 );
xor \U$10817 ( \11160 , \10691 , \10698 );
xor \U$10818 ( \11161 , \11159 , \11160 );
and \U$10819 ( \11162 , \11157 , \11161 );
and \U$10820 ( \11163 , \11143 , \11156 );
or \U$10821 ( \11164 , \11162 , \11163 );
xor \U$10822 ( \11165 , \10690 , \10703 );
xor \U$10823 ( \11166 , \11165 , \10796 );
and \U$10824 ( \11167 , \11164 , \11166 );
and \U$10825 ( \11168 , \10347 , \11164 );
or \U$10826 ( \11169 , \10798 , \11167 , \11168 );
xor \U$10827 ( \11170 , \10690 , \10703 );
and \U$10828 ( \11171 , \11170 , \10796 );
and \U$10829 ( \11172 , \10690 , \10703 );
or \U$10830 ( \11173 , \11171 , \11172 );
xor \U$10831 ( \11174 , \10708 , \10712 );
and \U$10832 ( \11175 , \11174 , \10721 );
and \U$10833 ( \11176 , \10708 , \10712 );
or \U$10834 ( \11177 , \11175 , \11176 );
and \U$10835 ( \11178 , \10736 , \10754 );
xor \U$10836 ( \11179 , \11177 , \11178 );
xor \U$10837 ( \11180 , \10761 , \10767 );
xor \U$10838 ( \11181 , \11180 , \10771 );
and \U$10839 ( \11182 , \10776 , \11181 );
xor \U$10840 ( \11183 , \10761 , \10767 );
xor \U$10841 ( \11184 , \11183 , \10771 );
and \U$10842 ( \11185 , \10792 , \11184 );
and \U$10843 ( \11186 , \10776 , \10792 );
or \U$10844 ( \11187 , \11182 , \11185 , \11186 );
xor \U$10845 ( \11188 , \11179 , \11187 );
xor \U$10846 ( \11189 , \11173 , \11188 );
xor \U$10847 ( \11190 , \10179 , \10248 );
and \U$10848 ( \11191 , \11190 , \10346 );
and \U$10849 ( \11192 , \10179 , \10248 );
or \U$10850 ( \11193 , \11191 , \11192 );
xor \U$10851 ( \11194 , \10708 , \10712 );
xor \U$10852 ( \11195 , \11194 , \10721 );
and \U$10853 ( \11196 , \10755 , \11195 );
xor \U$10854 ( \11197 , \10708 , \10712 );
xor \U$10855 ( \11198 , \11197 , \10721 );
and \U$10856 ( \11199 , \10794 , \11198 );
and \U$10857 ( \11200 , \10755 , \10794 );
or \U$10858 ( \11201 , \11196 , \11199 , \11200 );
xor \U$10859 ( \11202 , \11193 , \11201 );
xor \U$10860 ( \11203 , \10740 , \10748 );
and \U$10861 ( \11204 , \11203 , \10753 );
and \U$10862 ( \11205 , \10740 , \10748 );
or \U$10863 ( \11206 , \11204 , \11205 );
xor \U$10864 ( \11207 , \10726 , \10730 );
and \U$10865 ( \11208 , \11207 , \10735 );
and \U$10866 ( \11209 , \10726 , \10730 );
or \U$10867 ( \11210 , \11208 , \11209 );
xor \U$10868 ( \11211 , \11206 , \11210 );
xor \U$10869 ( \11212 , \10782 , \10788 );
and \U$10870 ( \11213 , \11212 , \10791 );
and \U$10871 ( \11214 , \10782 , \10788 );
or \U$10872 ( \11215 , \11213 , \11214 );
xor \U$10873 ( \11216 , \11211 , \11215 );
not \U$10874 ( \11217 , \9247 );
xor \U$10875 ( \11218 , \9399 , \9335 );
not \U$10876 ( \11219 , \11218 );
or \U$10877 ( \11220 , \11217 , \11219 );
or \U$10878 ( \11221 , \11218 , \9247 );
nand \U$10879 ( \11222 , \11220 , \11221 );
not \U$10880 ( \11223 , \9129 );
not \U$10881 ( \11224 , \9150 );
not \U$10882 ( \11225 , \9101 );
or \U$10883 ( \11226 , \11224 , \11225 );
or \U$10884 ( \11227 , \9101 , \9150 );
nand \U$10885 ( \11228 , \11226 , \11227 );
not \U$10886 ( \11229 , \11228 );
or \U$10887 ( \11230 , \11223 , \11229 );
or \U$10888 ( \11231 , \11228 , \9129 );
nand \U$10889 ( \11232 , \11230 , \11231 );
xor \U$10890 ( \11233 , \11222 , \11232 );
not \U$10891 ( \11234 , \9453 );
xor \U$10892 ( \11235 , \9450 , \9458 );
not \U$10893 ( \11236 , \11235 );
or \U$10894 ( \11237 , \11234 , \11236 );
or \U$10895 ( \11238 , \11235 , \9453 );
nand \U$10896 ( \11239 , \11237 , \11238 );
xor \U$10897 ( \11240 , \10761 , \10767 );
and \U$10898 ( \11241 , \11240 , \10771 );
and \U$10899 ( \11242 , \10761 , \10767 );
or \U$10900 ( \11243 , \11241 , \11242 );
xor \U$10901 ( \11244 , \11239 , \11243 );
not \U$10902 ( \11245 , \9418 );
not \U$10903 ( \11246 , \9412 );
not \U$10904 ( \11247 , \9427 );
or \U$10905 ( \11248 , \11246 , \11247 );
or \U$10906 ( \11249 , \9427 , \9412 );
nand \U$10907 ( \11250 , \11248 , \11249 );
not \U$10908 ( \11251 , \11250 );
or \U$10909 ( \11252 , \11245 , \11251 );
or \U$10910 ( \11253 , \11250 , \9418 );
nand \U$10911 ( \11254 , \11252 , \11253 );
xor \U$10912 ( \11255 , \11244 , \11254 );
xor \U$10913 ( \11256 , \11233 , \11255 );
xor \U$10914 ( \11257 , \11216 , \11256 );
xor \U$10915 ( \11258 , \11202 , \11257 );
xor \U$10916 ( \11259 , \11189 , \11258 );
and \U$10917 ( \11260 , \11169 , \11259 );
not \U$10918 ( \11261 , \11260 );
xor \U$10919 ( \11262 , \11173 , \11188 );
and \U$10920 ( \11263 , \11262 , \11258 );
and \U$10921 ( \11264 , \11173 , \11188 );
or \U$10922 ( \11265 , \11263 , \11264 );
xor \U$10923 ( \11266 , \11193 , \11201 );
and \U$10924 ( \11267 , \11266 , \11257 );
and \U$10925 ( \11268 , \11193 , \11201 );
or \U$10926 ( \11269 , \11267 , \11268 );
and \U$10927 ( \11270 , \11222 , \11232 );
xor \U$10928 ( \11271 , \11206 , \11210 );
and \U$10929 ( \11272 , \11271 , \11215 );
and \U$10930 ( \11273 , \11206 , \11210 );
or \U$10931 ( \11274 , \11272 , \11273 );
xor \U$10932 ( \11275 , \11270 , \11274 );
xor \U$10933 ( \11276 , \11239 , \11243 );
and \U$10934 ( \11277 , \11276 , \11254 );
and \U$10935 ( \11278 , \11239 , \11243 );
or \U$10936 ( \11279 , \11277 , \11278 );
xor \U$10937 ( \11280 , \11275 , \11279 );
xor \U$10938 ( \11281 , \11269 , \11280 );
xor \U$10939 ( \11282 , \9153 , \9401 );
xor \U$10940 ( \11283 , \11282 , \9430 );
not \U$10941 ( \11284 , \9446 );
not \U$10942 ( \11285 , \9435 );
and \U$10943 ( \11286 , \11284 , \11285 );
and \U$10944 ( \11287 , \9446 , \9435 );
nor \U$10945 ( \11288 , \11286 , \11287 );
xor \U$10946 ( \11289 , \8640 , \8642 );
xor \U$10947 ( \11290 , \11289 , \8645 );
xor \U$10948 ( \11291 , \9460 , \9467 );
xor \U$10949 ( \11292 , \11290 , \11291 );
xor \U$10950 ( \11293 , \11288 , \11292 );
xor \U$10951 ( \11294 , \11283 , \11293 );
not \U$10952 ( \11295 , \11294 );
xor \U$10953 ( \11296 , \11206 , \11210 );
xor \U$10954 ( \11297 , \11296 , \11215 );
and \U$10955 ( \11298 , \11233 , \11297 );
xor \U$10956 ( \11299 , \11206 , \11210 );
xor \U$10957 ( \11300 , \11299 , \11215 );
and \U$10958 ( \11301 , \11255 , \11300 );
and \U$10959 ( \11302 , \11233 , \11255 );
or \U$10960 ( \11303 , \11298 , \11301 , \11302 );
xor \U$10961 ( \11304 , \11177 , \11178 );
and \U$10962 ( \11305 , \11304 , \11187 );
and \U$10963 ( \11306 , \11177 , \11178 );
or \U$10964 ( \11307 , \11305 , \11306 );
xor \U$10965 ( \11308 , \11303 , \11307 );
not \U$10966 ( \11309 , \11308 );
or \U$10967 ( \11310 , \11295 , \11309 );
or \U$10968 ( \11311 , \11308 , \11294 );
nand \U$10969 ( \11312 , \11310 , \11311 );
xor \U$10970 ( \11313 , \11281 , \11312 );
xor \U$10971 ( \11314 , \11265 , \11313 );
not \U$10972 ( \11315 , \11314 );
or \U$10973 ( \11316 , \11261 , \11315 );
and \U$10974 ( \11317 , \4203 , RI986ef80_41);
and \U$10975 ( \11318 , RI986f250_47, \4201 );
nor \U$10976 ( \11319 , \11317 , \11318 );
and \U$10977 ( \11320 , \11319 , \4207 );
not \U$10978 ( \11321 , \11319 );
and \U$10979 ( \11322 , \11321 , \3922 );
nor \U$10980 ( \11323 , \11320 , \11322 );
not \U$10981 ( \11324 , \4519 );
and \U$10982 ( \11325 , \4710 , RI986f160_45);
and \U$10983 ( \11326 , RI986e530_19, \4708 );
nor \U$10984 ( \11327 , \11325 , \11326 );
not \U$10985 ( \11328 , \11327 );
or \U$10986 ( \11329 , \11324 , \11328 );
or \U$10987 ( \11330 , \11327 , \4519 );
nand \U$10988 ( \11331 , \11329 , \11330 );
xor \U$10989 ( \11332 , \11323 , \11331 );
and \U$10990 ( \11333 , \5318 , RI986e440_17);
and \U$10991 ( \11334 , RI986e710_23, \5316 );
nor \U$10992 ( \11335 , \11333 , \11334 );
and \U$10993 ( \11336 , \11335 , \5052 );
not \U$10994 ( \11337 , \11335 );
and \U$10995 ( \11338 , \11337 , \5322 );
nor \U$10996 ( \11339 , \11336 , \11338 );
and \U$10997 ( \11340 , \11332 , \11339 );
and \U$10998 ( \11341 , \11323 , \11331 );
or \U$10999 ( \11342 , \11340 , \11341 );
and \U$11000 ( \11343 , \2274 , RI986e9e0_29);
and \U$11001 ( \11344 , RI986e8f0_27, \2272 );
nor \U$11002 ( \11345 , \11343 , \11344 );
and \U$11003 ( \11346 , \11345 , \2030 );
not \U$11004 ( \11347 , \11345 );
and \U$11005 ( \11348 , \11347 , \2031 );
nor \U$11006 ( \11349 , \11346 , \11348 );
and \U$11007 ( \11350 , \1311 , RI98717d0_127);
and \U$11008 ( \11351 , RI9871500_121, \1309 );
nor \U$11009 ( \11352 , \11350 , \11351 );
and \U$11010 ( \11353 , \11352 , \1458 );
not \U$11011 ( \11354 , \11352 );
and \U$11012 ( \11355 , \11354 , \1318 );
nor \U$11013 ( \11356 , \11353 , \11355 );
xor \U$11014 ( \11357 , \11349 , \11356 );
not \U$11015 ( \11358 , \2034 );
and \U$11016 ( \11359 , \2042 , RI98715f0_123);
and \U$11017 ( \11360 , RI986ead0_31, \2040 );
nor \U$11018 ( \11361 , \11359 , \11360 );
not \U$11019 ( \11362 , \11361 );
or \U$11020 ( \11363 , \11358 , \11362 );
or \U$11021 ( \11364 , \11361 , \1462 );
nand \U$11022 ( \11365 , \11363 , \11364 );
and \U$11023 ( \11366 , \11357 , \11365 );
and \U$11024 ( \11367 , \11349 , \11356 );
or \U$11025 ( \11368 , \11366 , \11367 );
xor \U$11026 ( \11369 , \11342 , \11368 );
not \U$11027 ( \11370 , \3412 );
and \U$11028 ( \11371 , \3683 , RI986ecb0_35);
and \U$11029 ( \11372 , RI986f070_43, \3681 );
nor \U$11030 ( \11373 , \11371 , \11372 );
not \U$11031 ( \11374 , \11373 );
or \U$11032 ( \11375 , \11370 , \11374 );
or \U$11033 ( \11376 , \11373 , \3918 );
nand \U$11034 ( \11377 , \11375 , \11376 );
and \U$11035 ( \11378 , \2464 , RI986e800_25);
and \U$11036 ( \11379 , RI986ee90_39, \2462 );
nor \U$11037 ( \11380 , \11378 , \11379 );
and \U$11038 ( \11381 , \11380 , \2468 );
not \U$11039 ( \11382 , \11380 );
and \U$11040 ( \11383 , \11382 , \2263 );
nor \U$11041 ( \11384 , \11381 , \11383 );
xor \U$11042 ( \11385 , \11377 , \11384 );
not \U$11043 ( \11386 , \3406 );
and \U$11044 ( \11387 , \3254 , RI986eda0_37);
and \U$11045 ( \11388 , RI986ebc0_33, \3252 );
nor \U$11046 ( \11389 , \11387 , \11388 );
not \U$11047 ( \11390 , \11389 );
or \U$11048 ( \11391 , \11386 , \11390 );
or \U$11049 ( \11392 , \11389 , \2935 );
nand \U$11050 ( \11393 , \11391 , \11392 );
and \U$11051 ( \11394 , \11385 , \11393 );
and \U$11052 ( \11395 , \11377 , \11384 );
or \U$11053 ( \11396 , \11394 , \11395 );
xor \U$11054 ( \11397 , \11369 , \11396 );
not \U$11055 ( \11398 , \367 );
and \U$11056 ( \11399 , \376 , RI9870ab0_99);
and \U$11057 ( \11400 , RI9870d80_105, \374 );
nor \U$11058 ( \11401 , \11399 , \11400 );
not \U$11059 ( \11402 , \11401 );
or \U$11060 ( \11403 , \11398 , \11402 );
or \U$11061 ( \11404 , \11401 , \365 );
nand \U$11062 ( \11405 , \11403 , \11404 );
and \U$11063 ( \11406 , \438 , RI9870ba0_101);
and \U$11064 ( \11407 , RI9871050_111, \436 );
nor \U$11065 ( \11408 , \11406 , \11407 );
and \U$11066 ( \11409 , \11408 , \444 );
not \U$11067 ( \11410 , \11408 );
and \U$11068 ( \11411 , \11410 , \443 );
nor \U$11069 ( \11412 , \11409 , \11411 );
xor \U$11070 ( \11413 , \11405 , \11412 );
not \U$11071 ( \11414 , \456 );
and \U$11072 ( \11415 , \465 , RI98709c0_97);
and \U$11073 ( \11416 , RI9870e70_107, \463 );
nor \U$11074 ( \11417 , \11415 , \11416 );
not \U$11075 ( \11418 , \11417 );
or \U$11076 ( \11419 , \11414 , \11418 );
or \U$11077 ( \11420 , \11417 , \456 );
nand \U$11078 ( \11421 , \11419 , \11420 );
and \U$11079 ( \11422 , \11413 , \11421 );
and \U$11080 ( \11423 , \11405 , \11412 );
or \U$11081 ( \11424 , \11422 , \11423 );
and \U$11082 ( \11425 , \354 , RI986fe80_73);
and \U$11083 ( \11426 , RI9870060_77, \352 );
nor \U$11084 ( \11427 , \11425 , \11426 );
not \U$11085 ( \11428 , \11427 );
not \U$11086 ( \11429 , \345 );
and \U$11087 ( \11430 , \11428 , \11429 );
and \U$11088 ( \11431 , \11427 , \361 );
nor \U$11089 ( \11432 , \11430 , \11431 );
and \U$11090 ( \11433 , \416 , RI986fca0_69);
and \U$11091 ( \11434 , RI986ff70_75, \414 );
nor \U$11092 ( \11435 , \11433 , \11434 );
and \U$11093 ( \11436 , \11435 , \421 );
not \U$11094 ( \11437 , \11435 );
and \U$11095 ( \11438 , \11437 , \422 );
nor \U$11096 ( \11439 , \11436 , \11438 );
or \U$11097 ( \11440 , \11432 , \11439 );
not \U$11098 ( \11441 , \11439 );
not \U$11099 ( \11442 , \11432 );
or \U$11100 ( \11443 , \11441 , \11442 );
not \U$11101 ( \11444 , \386 );
and \U$11102 ( \11445 , \395 , RI9870150_79);
and \U$11103 ( \11446 , RI9870f60_109, \393 );
nor \U$11104 ( \11447 , \11445 , \11446 );
not \U$11105 ( \11448 , \11447 );
or \U$11106 ( \11449 , \11444 , \11448 );
or \U$11107 ( \11450 , \11447 , \386 );
nand \U$11108 ( \11451 , \11449 , \11450 );
nand \U$11109 ( \11452 , \11443 , \11451 );
nand \U$11110 ( \11453 , \11440 , \11452 );
xor \U$11111 ( \11454 , \11424 , \11453 );
and \U$11112 ( \11455 , \1329 , RI9871410_119);
and \U$11113 ( \11456 , RI98716e0_125, \1327 );
nor \U$11114 ( \11457 , \11455 , \11456 );
and \U$11115 ( \11458 , \11457 , \1336 );
not \U$11116 ( \11459 , \11457 );
and \U$11117 ( \11460 , \11459 , \1337 );
nor \U$11118 ( \11461 , \11458 , \11460 );
and \U$11119 ( \11462 , \776 , RI9870c90_103);
and \U$11120 ( \11463 , RI9871230_115, \774 );
nor \U$11121 ( \11464 , \11462 , \11463 );
and \U$11122 ( \11465 , \11464 , \474 );
not \U$11123 ( \11466 , \11464 );
and \U$11124 ( \11467 , \11466 , \451 );
nor \U$11125 ( \11468 , \11465 , \11467 );
xor \U$11126 ( \11469 , \11461 , \11468 );
not \U$11127 ( \11470 , \1301 );
and \U$11128 ( \11471 , \1293 , RI9871140_113);
and \U$11129 ( \11472 , RI9871320_117, \1291 );
nor \U$11130 ( \11473 , \11471 , \11472 );
not \U$11131 ( \11474 , \11473 );
or \U$11132 ( \11475 , \11470 , \11474 );
or \U$11133 ( \11476 , \11473 , \1128 );
nand \U$11134 ( \11477 , \11475 , \11476 );
and \U$11135 ( \11478 , \11469 , \11477 );
and \U$11136 ( \11479 , \11461 , \11468 );
or \U$11137 ( \11480 , \11478 , \11479 );
xor \U$11138 ( \11481 , \11454 , \11480 );
and \U$11139 ( \11482 , \11397 , \11481 );
xor \U$11140 ( \11483 , \10853 , \10860 );
xor \U$11141 ( \11484 , \11483 , \10869 );
not \U$11142 ( \11485 , RI986fca0_69);
nor \U$11143 ( \11486 , \11485 , \407 );
xor \U$11144 ( \11487 , \10879 , \10887 );
xor \U$11145 ( \11488 , \11487 , \10896 );
xor \U$11146 ( \11489 , \11486 , \11488 );
xor \U$11147 ( \11490 , \11484 , \11489 );
xor \U$11148 ( \11491 , \11424 , \11453 );
xor \U$11149 ( \11492 , \11491 , \11480 );
and \U$11150 ( \11493 , \11490 , \11492 );
and \U$11151 ( \11494 , \11397 , \11490 );
or \U$11152 ( \11495 , \11482 , \11493 , \11494 );
xor \U$11153 ( \11496 , \10954 , \10976 );
xor \U$11154 ( \11497 , \11496 , \11002 );
xor \U$11155 ( \11498 , \11495 , \11497 );
xor \U$11156 ( \11499 , \10872 , \10899 );
xor \U$11157 ( \11500 , \11499 , \10926 );
or \U$11158 ( \11501 , \10818 , \10828 );
nand \U$11159 ( \11502 , \11501 , \10829 );
xor \U$11160 ( \11503 , \11032 , \11059 );
xor \U$11161 ( \11504 , \11503 , \11086 );
xor \U$11162 ( \11505 , \11502 , \11504 );
xor \U$11163 ( \11506 , \11500 , \11505 );
and \U$11164 ( \11507 , \11498 , \11506 );
and \U$11165 ( \11508 , \11495 , \11497 );
or \U$11166 ( \11509 , \11507 , \11508 );
xor \U$11167 ( \11510 , \11377 , \11384 );
xor \U$11168 ( \11511 , \11510 , \11393 );
xor \U$11169 ( \11512 , \11323 , \11331 );
xor \U$11170 ( \11513 , \11512 , \11339 );
and \U$11171 ( \11514 , \11511 , \11513 );
and \U$11172 ( \11515 , \7079 , RI986f8e0_61);
and \U$11173 ( \11516 , RI986f430_51, \7077 );
nor \U$11174 ( \11517 , \11515 , \11516 );
and \U$11175 ( \11518 , \11517 , \6710 );
not \U$11176 ( \11519 , \11517 );
and \U$11177 ( \11520 , \11519 , \6709 );
nor \U$11178 ( \11521 , \11518 , \11520 );
and \U$11179 ( \11522 , \5881 , RI986e620_21);
and \U$11180 ( \11523 , RI986f7f0_59, \5879 );
nor \U$11181 ( \11524 , \11522 , \11523 );
and \U$11182 ( \11525 , \11524 , \5594 );
not \U$11183 ( \11526 , \11524 );
and \U$11184 ( \11527 , \11526 , \5885 );
nor \U$11185 ( \11528 , \11525 , \11527 );
xor \U$11186 ( \11529 , \11521 , \11528 );
and \U$11187 ( \11530 , \6453 , RI986f700_57);
and \U$11188 ( \11531 , RI986f9d0_63, \6451 );
nor \U$11189 ( \11532 , \11530 , \11531 );
and \U$11190 ( \11533 , \11532 , \6190 );
not \U$11191 ( \11534 , \11532 );
and \U$11192 ( \11535 , \11534 , \6705 );
nor \U$11193 ( \11536 , \11533 , \11535 );
xor \U$11194 ( \11537 , \11529 , \11536 );
xor \U$11195 ( \11538 , \11323 , \11331 );
xor \U$11196 ( \11539 , \11538 , \11339 );
and \U$11197 ( \11540 , \11537 , \11539 );
and \U$11198 ( \11541 , \11511 , \11537 );
or \U$11199 ( \11542 , \11514 , \11540 , \11541 );
nand \U$11200 ( \11543 , RI986fd90_71, RI9871fc8_144);
not \U$11201 ( \11544 , \11432 );
not \U$11202 ( \11545 , \11451 );
or \U$11203 ( \11546 , \11544 , \11545 );
or \U$11204 ( \11547 , \11432 , \11451 );
nand \U$11205 ( \11548 , \11546 , \11547 );
not \U$11206 ( \11549 , \11548 );
not \U$11207 ( \11550 , \11439 );
and \U$11208 ( \11551 , \11549 , \11550 );
and \U$11209 ( \11552 , \11548 , \11439 );
nor \U$11210 ( \11553 , \11551 , \11552 );
nand \U$11211 ( \11554 , \11543 , \11553 );
xor \U$11212 ( \11555 , \11542 , \11554 );
xor \U$11213 ( \11556 , \11461 , \11468 );
xor \U$11214 ( \11557 , \11556 , \11477 );
xor \U$11215 ( \11558 , \11405 , \11412 );
xor \U$11216 ( \11559 , \11558 , \11421 );
xor \U$11217 ( \11560 , \11557 , \11559 );
xor \U$11218 ( \11561 , \11349 , \11356 );
xor \U$11219 ( \11562 , \11561 , \11365 );
and \U$11220 ( \11563 , \11560 , \11562 );
and \U$11221 ( \11564 , \11557 , \11559 );
or \U$11222 ( \11565 , \11563 , \11564 );
and \U$11223 ( \11566 , \11555 , \11565 );
and \U$11224 ( \11567 , \11542 , \11554 );
or \U$11225 ( \11568 , \11566 , \11567 );
not \U$11226 ( \11569 , \456 );
and \U$11227 ( \11570 , \465 , RI9870d80_105);
and \U$11228 ( \11571 , RI98709c0_97, \463 );
nor \U$11229 ( \11572 , \11570 , \11571 );
not \U$11230 ( \11573 , \11572 );
or \U$11231 ( \11574 , \11569 , \11573 );
or \U$11232 ( \11575 , \11572 , \454 );
nand \U$11233 ( \11576 , \11574 , \11575 );
and \U$11234 ( \11577 , \776 , RI9871050_111);
and \U$11235 ( \11578 , RI9870c90_103, \774 );
nor \U$11236 ( \11579 , \11577 , \11578 );
and \U$11237 ( \11580 , \11579 , \474 );
not \U$11238 ( \11581 , \11579 );
and \U$11239 ( \11582 , \11581 , \451 );
nor \U$11240 ( \11583 , \11580 , \11582 );
xor \U$11241 ( \11584 , \11576 , \11583 );
and \U$11242 ( \11585 , \438 , RI9870e70_107);
and \U$11243 ( \11586 , RI9870ba0_101, \436 );
nor \U$11244 ( \11587 , \11585 , \11586 );
and \U$11245 ( \11588 , \11587 , \444 );
not \U$11246 ( \11589 , \11587 );
and \U$11247 ( \11590 , \11589 , \443 );
nor \U$11248 ( \11591 , \11588 , \11590 );
and \U$11249 ( \11592 , \11584 , \11591 );
and \U$11250 ( \11593 , \11576 , \11583 );
or \U$11251 ( \11594 , \11592 , \11593 );
not \U$11252 ( \11595 , \365 );
and \U$11253 ( \11596 , \376 , RI9870f60_109);
and \U$11254 ( \11597 , RI9870ab0_99, \374 );
nor \U$11255 ( \11598 , \11596 , \11597 );
not \U$11256 ( \11599 , \11598 );
or \U$11257 ( \11600 , \11595 , \11599 );
or \U$11258 ( \11601 , \11598 , \365 );
nand \U$11259 ( \11602 , \11600 , \11601 );
not \U$11260 ( \11603 , \487 );
and \U$11261 ( \11604 , \395 , RI9870060_77);
and \U$11262 ( \11605 , RI9870150_79, \393 );
nor \U$11263 ( \11606 , \11604 , \11605 );
not \U$11264 ( \11607 , \11606 );
or \U$11265 ( \11608 , \11603 , \11607 );
or \U$11266 ( \11609 , \11606 , \487 );
nand \U$11267 ( \11610 , \11608 , \11609 );
xor \U$11268 ( \11611 , \11602 , \11610 );
not \U$11269 ( \11612 , \361 );
and \U$11270 ( \11613 , \354 , RI986ff70_75);
and \U$11271 ( \11614 , RI986fe80_73, \352 );
nor \U$11272 ( \11615 , \11613 , \11614 );
not \U$11273 ( \11616 , \11615 );
or \U$11274 ( \11617 , \11612 , \11616 );
or \U$11275 ( \11618 , \11615 , \361 );
nand \U$11276 ( \11619 , \11617 , \11618 );
and \U$11277 ( \11620 , \11611 , \11619 );
and \U$11278 ( \11621 , \11602 , \11610 );
or \U$11279 ( \11622 , \11620 , \11621 );
xor \U$11280 ( \11623 , \11594 , \11622 );
and \U$11281 ( \11624 , \1311 , RI98716e0_125);
and \U$11282 ( \11625 , RI98717d0_127, \1309 );
nor \U$11283 ( \11626 , \11624 , \11625 );
and \U$11284 ( \11627 , \11626 , \1458 );
not \U$11285 ( \11628 , \11626 );
and \U$11286 ( \11629 , \11628 , \1318 );
nor \U$11287 ( \11630 , \11627 , \11629 );
not \U$11288 ( \11631 , \1128 );
and \U$11289 ( \11632 , \1293 , RI9871230_115);
and \U$11290 ( \11633 , RI9871140_113, \1291 );
nor \U$11291 ( \11634 , \11632 , \11633 );
not \U$11292 ( \11635 , \11634 );
or \U$11293 ( \11636 , \11631 , \11635 );
or \U$11294 ( \11637 , \11634 , \1128 );
nand \U$11295 ( \11638 , \11636 , \11637 );
xor \U$11296 ( \11639 , \11630 , \11638 );
and \U$11297 ( \11640 , \1329 , RI9871320_117);
and \U$11298 ( \11641 , RI9871410_119, \1327 );
nor \U$11299 ( \11642 , \11640 , \11641 );
and \U$11300 ( \11643 , \11642 , \1336 );
not \U$11301 ( \11644 , \11642 );
and \U$11302 ( \11645 , \11644 , \1337 );
nor \U$11303 ( \11646 , \11643 , \11645 );
and \U$11304 ( \11647 , \11639 , \11646 );
and \U$11305 ( \11648 , \11630 , \11638 );
or \U$11306 ( \11649 , \11647 , \11648 );
and \U$11307 ( \11650 , \11623 , \11649 );
and \U$11308 ( \11651 , \11594 , \11622 );
or \U$11309 ( \11652 , \11650 , \11651 );
and \U$11310 ( \11653 , \7079 , RI986f9d0_63);
and \U$11311 ( \11654 , RI986f8e0_61, \7077 );
nor \U$11312 ( \11655 , \11653 , \11654 );
and \U$11313 ( \11656 , \11655 , \6710 );
not \U$11314 ( \11657 , \11655 );
and \U$11315 ( \11658 , \11657 , \6709 );
nor \U$11316 ( \11659 , \11656 , \11658 );
and \U$11317 ( \11660 , \6453 , RI986f7f0_59);
and \U$11318 ( \11661 , RI986f700_57, \6451 );
nor \U$11319 ( \11662 , \11660 , \11661 );
and \U$11320 ( \11663 , \11662 , \6190 );
not \U$11321 ( \11664 , \11662 );
and \U$11322 ( \11665 , \11664 , \6180 );
nor \U$11323 ( \11666 , \11663 , \11665 );
xor \U$11324 ( \11667 , \11659 , \11666 );
and \U$11325 ( \11668 , \7729 , RI986f430_51);
and \U$11326 ( \11669 , RI986f340_49, \7727 );
nor \U$11327 ( \11670 , \11668 , \11669 );
and \U$11328 ( \11671 , \11670 , \7480 );
not \U$11329 ( \11672 , \11670 );
and \U$11330 ( \11673 , \11672 , \7733 );
nor \U$11331 ( \11674 , \11671 , \11673 );
and \U$11332 ( \11675 , \11667 , \11674 );
and \U$11333 ( \11676 , \11659 , \11666 );
or \U$11334 ( \11677 , \11675 , \11676 );
and \U$11335 ( \11678 , \10424 , RI986e170_11);
and \U$11336 ( \11679 , RI986e080_9, \10422 );
nor \U$11337 ( \11680 , \11678 , \11679 );
and \U$11338 ( \11681 , \11680 , \9840 );
not \U$11339 ( \11682 , \11680 );
and \U$11340 ( \11683 , \11682 , \10428 );
nor \U$11341 ( \11684 , \11681 , \11683 );
nand \U$11342 ( \11685 , RI9873288_184, RI9873300_185);
and \U$11343 ( \11686 , \11685 , RI9873210_183);
not \U$11344 ( \11687 , \11686 );
xor \U$11345 ( \11688 , \11684 , \11687 );
and \U$11346 ( \11689 , RI98730a8_180, RI9873198_182);
not \U$11347 ( \11690 , RI9873198_182);
nor \U$11348 ( \11691 , \11690 , RI9873210_183);
not \U$11349 ( \11692 , RI9873210_183);
nor \U$11350 ( \11693 , \11692 , RI9873198_182);
or \U$11351 ( \11694 , \11691 , \11693 );
nor \U$11352 ( \11695 , RI98730a8_180, RI9873198_182);
nor \U$11353 ( \11696 , \11689 , \11694 , \11695 );
and \U$11354 ( \11697 , \11696 , RI986e260_13);
and \U$11355 ( \11698 , RI986e350_15, \11694 );
nor \U$11356 ( \11699 , \11697 , \11698 );
and \U$11357 ( \11700 , \11699 , \10965 );
not \U$11358 ( \11701 , \11699 );
not \U$11359 ( \11702 , \10965 );
and \U$11360 ( \11703 , \11701 , \11702 );
nor \U$11361 ( \11704 , \11700 , \11703 );
and \U$11362 ( \11705 , \11688 , \11704 );
and \U$11363 ( \11706 , \11684 , \11687 );
or \U$11364 ( \11707 , \11705 , \11706 );
xor \U$11365 ( \11708 , \11677 , \11707 );
and \U$11366 ( \11709 , \9237 , RI986df90_7);
and \U$11367 ( \11710 , RI986dea0_5, \9235 );
nor \U$11368 ( \11711 , \11709 , \11710 );
and \U$11369 ( \11712 , \11711 , \9241 );
not \U$11370 ( \11713 , \11711 );
and \U$11371 ( \11714 , \11713 , \8836 );
nor \U$11372 ( \11715 , \11712 , \11714 );
and \U$11373 ( \11716 , \8486 , RI986f520_53);
and \U$11374 ( \11717 , RI986f610_55, \8484 );
nor \U$11375 ( \11718 , \11716 , \11717 );
and \U$11376 ( \11719 , \11718 , \8050 );
not \U$11377 ( \11720 , \11718 );
and \U$11378 ( \11721 , \11720 , \8051 );
nor \U$11379 ( \11722 , \11719 , \11721 );
xor \U$11380 ( \11723 , \11715 , \11722 );
and \U$11381 ( \11724 , \9505 , RI986ddb0_3);
and \U$11382 ( \11725 , RI986dcc0_1, \9503 );
nor \U$11383 ( \11726 , \11724 , \11725 );
and \U$11384 ( \11727 , \11726 , \9510 );
not \U$11385 ( \11728 , \11726 );
and \U$11386 ( \11729 , \11728 , \9513 );
nor \U$11387 ( \11730 , \11727 , \11729 );
and \U$11388 ( \11731 , \11723 , \11730 );
and \U$11389 ( \11732 , \11715 , \11722 );
or \U$11390 ( \11733 , \11731 , \11732 );
and \U$11391 ( \11734 , \11708 , \11733 );
and \U$11392 ( \11735 , \11677 , \11707 );
or \U$11393 ( \11736 , \11734 , \11735 );
xor \U$11394 ( \11737 , \11652 , \11736 );
not \U$11395 ( \11738 , \4519 );
and \U$11396 ( \11739 , \4710 , RI986f250_47);
and \U$11397 ( \11740 , RI986f160_45, \4708 );
nor \U$11398 ( \11741 , \11739 , \11740 );
not \U$11399 ( \11742 , \11741 );
or \U$11400 ( \11743 , \11738 , \11742 );
or \U$11401 ( \11744 , \11741 , \4521 );
nand \U$11402 ( \11745 , \11743 , \11744 );
and \U$11403 ( \11746 , \5318 , RI986e530_19);
and \U$11404 ( \11747 , RI986e440_17, \5316 );
nor \U$11405 ( \11748 , \11746 , \11747 );
and \U$11406 ( \11749 , \11748 , \5052 );
not \U$11407 ( \11750 , \11748 );
and \U$11408 ( \11751 , \11750 , \5322 );
nor \U$11409 ( \11752 , \11749 , \11751 );
xor \U$11410 ( \11753 , \11745 , \11752 );
and \U$11411 ( \11754 , \5881 , RI986e710_23);
and \U$11412 ( \11755 , RI986e620_21, \5879 );
nor \U$11413 ( \11756 , \11754 , \11755 );
and \U$11414 ( \11757 , \11756 , \5594 );
not \U$11415 ( \11758 , \11756 );
and \U$11416 ( \11759 , \11758 , \5885 );
nor \U$11417 ( \11760 , \11757 , \11759 );
and \U$11418 ( \11761 , \11753 , \11760 );
and \U$11419 ( \11762 , \11745 , \11752 );
or \U$11420 ( \11763 , \11761 , \11762 );
and \U$11421 ( \11764 , \2464 , RI986e8f0_27);
and \U$11422 ( \11765 , RI986e800_25, \2462 );
nor \U$11423 ( \11766 , \11764 , \11765 );
and \U$11424 ( \11767 , \11766 , \2468 );
not \U$11425 ( \11768 , \11766 );
and \U$11426 ( \11769 , \11768 , \2263 );
nor \U$11427 ( \11770 , \11767 , \11769 );
not \U$11428 ( \11771 , \2034 );
and \U$11429 ( \11772 , \2042 , RI9871500_121);
and \U$11430 ( \11773 , RI98715f0_123, \2040 );
nor \U$11431 ( \11774 , \11772 , \11773 );
not \U$11432 ( \11775 , \11774 );
or \U$11433 ( \11776 , \11771 , \11775 );
or \U$11434 ( \11777 , \11774 , \1462 );
nand \U$11435 ( \11778 , \11776 , \11777 );
xor \U$11436 ( \11779 , \11770 , \11778 );
and \U$11437 ( \11780 , \2274 , RI986ead0_31);
and \U$11438 ( \11781 , RI986e9e0_29, \2272 );
nor \U$11439 ( \11782 , \11780 , \11781 );
and \U$11440 ( \11783 , \11782 , \2030 );
not \U$11441 ( \11784 , \11782 );
and \U$11442 ( \11785 , \11784 , \2031 );
nor \U$11443 ( \11786 , \11783 , \11785 );
and \U$11444 ( \11787 , \11779 , \11786 );
and \U$11445 ( \11788 , \11770 , \11778 );
or \U$11446 ( \11789 , \11787 , \11788 );
xor \U$11447 ( \11790 , \11763 , \11789 );
not \U$11448 ( \11791 , \3918 );
and \U$11449 ( \11792 , \3683 , RI986ebc0_33);
and \U$11450 ( \11793 , RI986ecb0_35, \3681 );
nor \U$11451 ( \11794 , \11792 , \11793 );
not \U$11452 ( \11795 , \11794 );
or \U$11453 ( \11796 , \11791 , \11795 );
or \U$11454 ( \11797 , \11794 , \3412 );
nand \U$11455 ( \11798 , \11796 , \11797 );
not \U$11456 ( \11799 , \2935 );
and \U$11457 ( \11800 , \3254 , RI986ee90_39);
and \U$11458 ( \11801 , RI986eda0_37, \3252 );
nor \U$11459 ( \11802 , \11800 , \11801 );
not \U$11460 ( \11803 , \11802 );
or \U$11461 ( \11804 , \11799 , \11803 );
or \U$11462 ( \11805 , \11802 , \2935 );
nand \U$11463 ( \11806 , \11804 , \11805 );
xor \U$11464 ( \11807 , \11798 , \11806 );
and \U$11465 ( \11808 , \4203 , RI986f070_43);
and \U$11466 ( \11809 , RI986ef80_41, \4201 );
nor \U$11467 ( \11810 , \11808 , \11809 );
and \U$11468 ( \11811 , \11810 , \4207 );
not \U$11469 ( \11812 , \11810 );
and \U$11470 ( \11813 , \11812 , \3922 );
nor \U$11471 ( \11814 , \11811 , \11813 );
and \U$11472 ( \11815 , \11807 , \11814 );
and \U$11473 ( \11816 , \11798 , \11806 );
or \U$11474 ( \11817 , \11815 , \11816 );
and \U$11475 ( \11818 , \11790 , \11817 );
and \U$11476 ( \11819 , \11763 , \11789 );
or \U$11477 ( \11820 , \11818 , \11819 );
and \U$11478 ( \11821 , \11737 , \11820 );
and \U$11479 ( \11822 , \11652 , \11736 );
or \U$11480 ( \11823 , \11821 , \11822 );
xor \U$11481 ( \11824 , \11568 , \11823 );
xor \U$11482 ( \11825 , \10961 , \10965 );
xor \U$11483 ( \11826 , \11825 , \10973 );
xor \U$11484 ( \11827 , \10936 , \10943 );
xor \U$11485 ( \11828 , \11827 , \10951 );
xor \U$11486 ( \11829 , \11013 , \11021 );
xor \U$11487 ( \11830 , \11829 , \11029 );
xor \U$11488 ( \11831 , \11828 , \11830 );
xor \U$11489 ( \11832 , \10984 , \10991 );
xor \U$11490 ( \11833 , \11832 , \10999 );
xor \U$11491 ( \11834 , \11831 , \11833 );
and \U$11492 ( \11835 , \11826 , \11834 );
xor \U$11493 ( \11836 , \10908 , \10915 );
xor \U$11494 ( \11837 , \11836 , \10923 );
xor \U$11495 ( \11838 , \11067 , \11075 );
xor \U$11496 ( \11839 , \11838 , \11083 );
xor \U$11497 ( \11840 , \11040 , \11047 );
xor \U$11498 ( \11841 , \11840 , \11056 );
xor \U$11499 ( \11842 , \11839 , \11841 );
xor \U$11500 ( \11843 , \11837 , \11842 );
xor \U$11501 ( \11844 , \11828 , \11830 );
xor \U$11502 ( \11845 , \11844 , \11833 );
and \U$11503 ( \11846 , \11843 , \11845 );
and \U$11504 ( \11847 , \11826 , \11843 );
or \U$11505 ( \11848 , \11835 , \11846 , \11847 );
and \U$11506 ( \11849 , \11824 , \11848 );
and \U$11507 ( \11850 , \11568 , \11823 );
or \U$11508 ( \11851 , \11849 , \11850 );
xor \U$11509 ( \11852 , \11509 , \11851 );
xor \U$11510 ( \11853 , \11424 , \11453 );
and \U$11511 ( \11854 , \11853 , \11480 );
and \U$11512 ( \11855 , \11424 , \11453 );
or \U$11513 ( \11856 , \11854 , \11855 );
and \U$11514 ( \11857 , \9237 , RI986dea0_5);
and \U$11515 ( \11858 , RI986ddb0_3, \9235 );
nor \U$11516 ( \11859 , \11857 , \11858 );
and \U$11517 ( \11860 , \11859 , \9241 );
not \U$11518 ( \11861 , \11859 );
and \U$11519 ( \11862 , \11861 , \8836 );
nor \U$11520 ( \11863 , \11860 , \11862 );
and \U$11521 ( \11864 , \7729 , RI986f340_49);
and \U$11522 ( \11865 , RI986f520_53, \7727 );
nor \U$11523 ( \11866 , \11864 , \11865 );
and \U$11524 ( \11867 , \11866 , \7480 );
not \U$11525 ( \11868 , \11866 );
and \U$11526 ( \11869 , \11868 , \7733 );
nor \U$11527 ( \11870 , \11867 , \11869 );
xor \U$11528 ( \11871 , \11863 , \11870 );
and \U$11529 ( \11872 , \8486 , RI986f610_55);
and \U$11530 ( \11873 , RI986df90_7, \8484 );
nor \U$11531 ( \11874 , \11872 , \11873 );
and \U$11532 ( \11875 , \11874 , \8050 );
not \U$11533 ( \11876 , \11874 );
and \U$11534 ( \11877 , \11876 , \8051 );
nor \U$11535 ( \11878 , \11875 , \11877 );
and \U$11536 ( \11879 , \11871 , \11878 );
and \U$11537 ( \11880 , \11863 , \11870 );
or \U$11538 ( \11881 , \11879 , \11880 );
xor \U$11539 ( \11882 , \11521 , \11528 );
and \U$11540 ( \11883 , \11882 , \11536 );
and \U$11541 ( \11884 , \11521 , \11528 );
or \U$11542 ( \11885 , \11883 , \11884 );
xor \U$11543 ( \11886 , \11881 , \11885 );
and \U$11544 ( \11887 , \9505 , RI986dcc0_1);
and \U$11545 ( \11888 , RI986e170_11, \9503 );
nor \U$11546 ( \11889 , \11887 , \11888 );
and \U$11547 ( \11890 , \11889 , \9510 );
not \U$11548 ( \11891 , \11889 );
and \U$11549 ( \11892 , \11891 , \9513 );
nor \U$11550 ( \11893 , \11890 , \11892 );
nand \U$11551 ( \11894 , RI986e350_15, \11696 );
and \U$11552 ( \11895 , \11894 , \10965 );
not \U$11553 ( \11896 , \11894 );
and \U$11554 ( \11897 , \11896 , \11702 );
nor \U$11555 ( \11898 , \11895 , \11897 );
xor \U$11556 ( \11899 , \11893 , \11898 );
and \U$11557 ( \11900 , \10424 , RI986e080_9);
and \U$11558 ( \11901 , RI986e260_13, \10422 );
nor \U$11559 ( \11902 , \11900 , \11901 );
and \U$11560 ( \11903 , \11902 , \9840 );
not \U$11561 ( \11904 , \11902 );
and \U$11562 ( \11905 , \11904 , \10428 );
nor \U$11563 ( \11906 , \11903 , \11905 );
and \U$11564 ( \11907 , \11899 , \11906 );
and \U$11565 ( \11908 , \11893 , \11898 );
or \U$11566 ( \11909 , \11907 , \11908 );
and \U$11567 ( \11910 , \11886 , \11909 );
and \U$11568 ( \11911 , \11881 , \11885 );
or \U$11569 ( \11912 , \11910 , \11911 );
xor \U$11570 ( \11913 , \11856 , \11912 );
xor \U$11571 ( \11914 , \11342 , \11368 );
and \U$11572 ( \11915 , \11914 , \11396 );
and \U$11573 ( \11916 , \11342 , \11368 );
or \U$11574 ( \11917 , \11915 , \11916 );
xor \U$11575 ( \11918 , \11913 , \11917 );
xor \U$11576 ( \11919 , \10908 , \10915 );
xor \U$11577 ( \11920 , \11919 , \10923 );
and \U$11578 ( \11921 , \11839 , \11920 );
xor \U$11579 ( \11922 , \10908 , \10915 );
xor \U$11580 ( \11923 , \11922 , \10923 );
and \U$11581 ( \11924 , \11841 , \11923 );
and \U$11582 ( \11925 , \11839 , \11841 );
or \U$11583 ( \11926 , \11921 , \11924 , \11925 );
xor \U$11584 ( \11927 , \10853 , \10860 );
xor \U$11585 ( \11928 , \11927 , \10869 );
and \U$11586 ( \11929 , \11486 , \11928 );
xor \U$11587 ( \11930 , \10853 , \10860 );
xor \U$11588 ( \11931 , \11930 , \10869 );
and \U$11589 ( \11932 , \11488 , \11931 );
and \U$11590 ( \11933 , \11486 , \11488 );
or \U$11591 ( \11934 , \11929 , \11932 , \11933 );
xor \U$11592 ( \11935 , \11926 , \11934 );
xor \U$11593 ( \11936 , \11828 , \11830 );
and \U$11594 ( \11937 , \11936 , \11833 );
and \U$11595 ( \11938 , \11828 , \11830 );
or \U$11596 ( \11939 , \11937 , \11938 );
xor \U$11597 ( \11940 , \11935 , \11939 );
and \U$11598 ( \11941 , \11918 , \11940 );
xor \U$11599 ( \11942 , \10800 , \10802 );
xor \U$11600 ( \11943 , \11942 , \10805 );
xor \U$11601 ( \11944 , \10417 , \10430 );
xor \U$11602 ( \11945 , \11944 , \10438 );
xor \U$11603 ( \11946 , \10587 , \10594 );
xor \U$11604 ( \11947 , \11946 , \10603 );
xor \U$11605 ( \11948 , \10832 , \10837 );
xor \U$11606 ( \11949 , \11947 , \11948 );
xor \U$11607 ( \11950 , \11945 , \11949 );
xor \U$11608 ( \11951 , \11943 , \11950 );
xor \U$11609 ( \11952 , \11926 , \11934 );
xor \U$11610 ( \11953 , \11952 , \11939 );
and \U$11611 ( \11954 , \11951 , \11953 );
and \U$11612 ( \11955 , \11918 , \11951 );
or \U$11613 ( \11956 , \11941 , \11954 , \11955 );
and \U$11614 ( \11957 , \11852 , \11956 );
and \U$11615 ( \11958 , \11509 , \11851 );
or \U$11616 ( \11959 , \11957 , \11958 );
xor \U$11617 ( \11960 , \10929 , \11005 );
xor \U$11618 ( \11961 , \11960 , \11089 );
xor \U$11619 ( \11962 , \10808 , \10829 );
xor \U$11620 ( \11963 , \11962 , \10842 );
xor \U$11621 ( \11964 , \11961 , \11963 );
xor \U$11622 ( \11965 , \11926 , \11934 );
and \U$11623 ( \11966 , \11965 , \11939 );
and \U$11624 ( \11967 , \11926 , \11934 );
or \U$11625 ( \11968 , \11966 , \11967 );
xor \U$11626 ( \11969 , \11856 , \11912 );
and \U$11627 ( \11970 , \11969 , \11917 );
and \U$11628 ( \11971 , \11856 , \11912 );
or \U$11629 ( \11972 , \11970 , \11971 );
xor \U$11630 ( \11973 , \11968 , \11972 );
xor \U$11631 ( \11974 , \10800 , \10802 );
xor \U$11632 ( \11975 , \11974 , \10805 );
and \U$11633 ( \11976 , \11945 , \11975 );
xor \U$11634 ( \11977 , \10800 , \10802 );
xor \U$11635 ( \11978 , \11977 , \10805 );
and \U$11636 ( \11979 , \11949 , \11978 );
and \U$11637 ( \11980 , \11945 , \11949 );
or \U$11638 ( \11981 , \11976 , \11979 , \11980 );
xor \U$11639 ( \11982 , \11973 , \11981 );
and \U$11640 ( \11983 , \11964 , \11982 );
xor \U$11641 ( \11984 , \11120 , \11122 );
xor \U$11642 ( \11985 , \11984 , \11125 );
xor \U$11643 ( \11986 , \10872 , \10899 );
xor \U$11644 ( \11987 , \11986 , \10926 );
and \U$11645 ( \11988 , \11502 , \11987 );
xor \U$11646 ( \11989 , \10872 , \10899 );
xor \U$11647 ( \11990 , \11989 , \10926 );
and \U$11648 ( \11991 , \11504 , \11990 );
and \U$11649 ( \11992 , \11502 , \11504 );
or \U$11650 ( \11993 , \11988 , \11991 , \11992 );
xor \U$11651 ( \11994 , \10361 , \10363 );
xor \U$11652 ( \11995 , \11994 , \10366 );
xor \U$11653 ( \11996 , \11097 , \11104 );
xor \U$11654 ( \11997 , \11995 , \11996 );
xor \U$11655 ( \11998 , \11993 , \11997 );
xor \U$11656 ( \11999 , \11985 , \11998 );
xor \U$11657 ( \12000 , \11968 , \11972 );
xor \U$11658 ( \12001 , \12000 , \11981 );
and \U$11659 ( \12002 , \11999 , \12001 );
and \U$11660 ( \12003 , \11964 , \11999 );
or \U$11661 ( \12004 , \11983 , \12002 , \12003 );
xor \U$11662 ( \12005 , \11959 , \12004 );
xor \U$11663 ( \12006 , \10845 , \11092 );
xor \U$11664 ( \12007 , \12006 , \11109 );
xor \U$11665 ( \12008 , \11114 , \11116 );
xor \U$11666 ( \12009 , \10667 , \10669 );
xor \U$11667 ( \12010 , \12009 , \10672 );
xor \U$11668 ( \12011 , \11128 , \11135 );
xor \U$11669 ( \12012 , \12010 , \12011 );
xor \U$11670 ( \12013 , \12008 , \12012 );
xor \U$11671 ( \12014 , \12007 , \12013 );
and \U$11672 ( \12015 , \12005 , \12014 );
and \U$11673 ( \12016 , \11959 , \12004 );
or \U$11674 ( \12017 , \12015 , \12016 );
xor \U$11675 ( \12018 , \11112 , \11117 );
xor \U$11676 ( \12019 , \12018 , \11140 );
xor \U$11677 ( \12020 , \12017 , \12019 );
xor \U$11678 ( \12021 , \11968 , \11972 );
and \U$11679 ( \12022 , \12021 , \11981 );
and \U$11680 ( \12023 , \11968 , \11972 );
or \U$11681 ( \12024 , \12022 , \12023 );
and \U$11682 ( \12025 , \11961 , \11963 );
xor \U$11683 ( \12026 , \12024 , \12025 );
xor \U$11684 ( \12027 , \11120 , \11122 );
xor \U$11685 ( \12028 , \12027 , \11125 );
and \U$11686 ( \12029 , \11993 , \12028 );
xor \U$11687 ( \12030 , \11120 , \11122 );
xor \U$11688 ( \12031 , \12030 , \11125 );
and \U$11689 ( \12032 , \11997 , \12031 );
and \U$11690 ( \12033 , \11993 , \11997 );
or \U$11691 ( \12034 , \12029 , \12032 , \12033 );
and \U$11692 ( \12035 , \12026 , \12034 );
and \U$11693 ( \12036 , \12024 , \12025 );
or \U$11694 ( \12037 , \12035 , \12036 );
xor \U$11695 ( \12038 , \10845 , \11092 );
xor \U$11696 ( \12039 , \12038 , \11109 );
and \U$11697 ( \12040 , \12008 , \12039 );
xor \U$11698 ( \12041 , \10845 , \11092 );
xor \U$11699 ( \12042 , \12041 , \11109 );
and \U$11700 ( \12043 , \12012 , \12042 );
and \U$11701 ( \12044 , \12008 , \12012 );
or \U$11702 ( \12045 , \12040 , \12043 , \12044 );
xor \U$11703 ( \12046 , \12037 , \12045 );
xor \U$11704 ( \12047 , \10385 , \10639 );
xor \U$11705 ( \12048 , \12047 , \10656 );
xor \U$11706 ( \12049 , \11144 , \11151 );
xor \U$11707 ( \12050 , \12048 , \12049 );
xor \U$11708 ( \12051 , \12046 , \12050 );
and \U$11709 ( \12052 , \12020 , \12051 );
and \U$11710 ( \12053 , \12017 , \12019 );
or \U$11711 ( \12054 , \12052 , \12053 );
xor \U$11712 ( \12055 , \12037 , \12045 );
and \U$11713 ( \12056 , \12055 , \12050 );
and \U$11714 ( \12057 , \12037 , \12045 );
or \U$11715 ( \12058 , \12056 , \12057 );
xor \U$11716 ( \12059 , \10659 , \10664 );
xor \U$11717 ( \12060 , \12059 , \10687 );
xor \U$11718 ( \12061 , \12058 , \12060 );
xor \U$11719 ( \12062 , \11143 , \11156 );
xor \U$11720 ( \12063 , \12062 , \11161 );
xor \U$11721 ( \12064 , \12061 , \12063 );
and \U$11722 ( \12065 , \12054 , \12064 );
not \U$11723 ( \12066 , \12065 );
xor \U$11724 ( \12067 , \12058 , \12060 );
and \U$11725 ( \12068 , \12067 , \12063 );
and \U$11726 ( \12069 , \12058 , \12060 );
or \U$11727 ( \12070 , \12068 , \12069 );
xor \U$11728 ( \12071 , \10690 , \10703 );
xor \U$11729 ( \12072 , \12071 , \10796 );
xor \U$11730 ( \12073 , \10347 , \11164 );
xor \U$11731 ( \12074 , \12072 , \12073 );
xor \U$11732 ( \12075 , \12070 , \12074 );
not \U$11733 ( \12076 , \12075 );
or \U$11734 ( \12077 , \12066 , \12076 );
xor \U$11735 ( \12078 , \11652 , \11736 );
xor \U$11736 ( \12079 , \12078 , \11820 );
xor \U$11737 ( \12080 , \11677 , \11707 );
xor \U$11738 ( \12081 , \12080 , \11733 );
xor \U$11739 ( \12082 , \11594 , \11622 );
xor \U$11740 ( \12083 , \12082 , \11649 );
xor \U$11741 ( \12084 , \12081 , \12083 );
xor \U$11742 ( \12085 , \11763 , \11789 );
xor \U$11743 ( \12086 , \12085 , \11817 );
and \U$11744 ( \12087 , \12084 , \12086 );
and \U$11745 ( \12088 , \12081 , \12083 );
or \U$11746 ( \12089 , \12087 , \12088 );
xor \U$11747 ( \12090 , \11881 , \11885 );
xor \U$11748 ( \12091 , \12090 , \11909 );
xor \U$11749 ( \12092 , \12089 , \12091 );
or \U$11750 ( \12093 , \11553 , \11543 );
nand \U$11751 ( \12094 , \12093 , \11554 );
xor \U$11752 ( \12095 , \11557 , \11559 );
xor \U$11753 ( \12096 , \12095 , \11562 );
and \U$11754 ( \12097 , \12094 , \12096 );
xor \U$11755 ( \12098 , \11323 , \11331 );
xor \U$11756 ( \12099 , \12098 , \11339 );
xor \U$11757 ( \12100 , \11511 , \11537 );
xor \U$11758 ( \12101 , \12099 , \12100 );
xor \U$11759 ( \12102 , \11557 , \11559 );
xor \U$11760 ( \12103 , \12102 , \11562 );
and \U$11761 ( \12104 , \12101 , \12103 );
and \U$11762 ( \12105 , \12094 , \12101 );
or \U$11763 ( \12106 , \12097 , \12104 , \12105 );
xor \U$11764 ( \12107 , \12092 , \12106 );
and \U$11765 ( \12108 , \12079 , \12107 );
xor \U$11766 ( \12109 , \11542 , \11554 );
xor \U$11767 ( \12110 , \12109 , \11565 );
xor \U$11768 ( \12111 , \11424 , \11453 );
xor \U$11769 ( \12112 , \12111 , \11480 );
xor \U$11770 ( \12113 , \11397 , \11490 );
xor \U$11771 ( \12114 , \12112 , \12113 );
xor \U$11772 ( \12115 , \11828 , \11830 );
xor \U$11773 ( \12116 , \12115 , \11833 );
xor \U$11774 ( \12117 , \11826 , \11843 );
xor \U$11775 ( \12118 , \12116 , \12117 );
xor \U$11776 ( \12119 , \12114 , \12118 );
xor \U$11777 ( \12120 , \12110 , \12119 );
xor \U$11778 ( \12121 , \12089 , \12091 );
xor \U$11779 ( \12122 , \12121 , \12106 );
and \U$11780 ( \12123 , \12120 , \12122 );
and \U$11781 ( \12124 , \12079 , \12120 );
or \U$11782 ( \12125 , \12108 , \12123 , \12124 );
xor \U$11783 ( \12126 , \11602 , \11610 );
xor \U$11784 ( \12127 , \12126 , \11619 );
xor \U$11785 ( \12128 , \11576 , \11583 );
xor \U$11786 ( \12129 , \12128 , \11591 );
and \U$11787 ( \12130 , \12127 , \12129 );
xor \U$11788 ( \12131 , \11630 , \11638 );
xor \U$11789 ( \12132 , \12131 , \11646 );
xor \U$11790 ( \12133 , \11576 , \11583 );
xor \U$11791 ( \12134 , \12133 , \11591 );
and \U$11792 ( \12135 , \12132 , \12134 );
and \U$11793 ( \12136 , \12127 , \12132 );
or \U$11794 ( \12137 , \12130 , \12135 , \12136 );
and \U$11795 ( \12138 , \416 , RI986fd90_71);
and \U$11796 ( \12139 , RI986fca0_69, \414 );
nor \U$11797 ( \12140 , \12138 , \12139 );
and \U$11798 ( \12141 , \12140 , \422 );
not \U$11799 ( \12142 , \12140 );
and \U$11800 ( \12143 , \12142 , \421 );
nor \U$11801 ( \12144 , \12141 , \12143 );
not \U$11802 ( \12145 , RI986fbb0_67);
nor \U$11803 ( \12146 , \12145 , \407 );
xor \U$11804 ( \12147 , \12144 , \12146 );
nand \U$11805 ( \12148 , RI986fac0_65, RI9871fc8_144);
and \U$11806 ( \12149 , \416 , RI986fbb0_67);
and \U$11807 ( \12150 , RI986fd90_71, \414 );
nor \U$11808 ( \12151 , \12149 , \12150 );
and \U$11809 ( \12152 , \12151 , \421 );
not \U$11810 ( \12153 , \12151 );
and \U$11811 ( \12154 , \12153 , \422 );
nor \U$11812 ( \12155 , \12152 , \12154 );
nand \U$11813 ( \12156 , \12148 , \12155 );
and \U$11814 ( \12157 , \12147 , \12156 );
and \U$11815 ( \12158 , \12144 , \12146 );
or \U$11816 ( \12159 , \12157 , \12158 );
xor \U$11817 ( \12160 , \12137 , \12159 );
xor \U$11818 ( \12161 , \11798 , \11806 );
xor \U$11819 ( \12162 , \12161 , \11814 );
xor \U$11820 ( \12163 , \11770 , \11778 );
xor \U$11821 ( \12164 , \12163 , \11786 );
xor \U$11822 ( \12165 , \12162 , \12164 );
xor \U$11823 ( \12166 , \11745 , \11752 );
xor \U$11824 ( \12167 , \12166 , \11760 );
and \U$11825 ( \12168 , \12165 , \12167 );
and \U$11826 ( \12169 , \12162 , \12164 );
or \U$11827 ( \12170 , \12168 , \12169 );
xor \U$11828 ( \12171 , \12160 , \12170 );
and \U$11829 ( \12172 , \4203 , RI986ecb0_35);
and \U$11830 ( \12173 , RI986f070_43, \4201 );
nor \U$11831 ( \12174 , \12172 , \12173 );
and \U$11832 ( \12175 , \12174 , \4207 );
not \U$11833 ( \12176 , \12174 );
and \U$11834 ( \12177 , \12176 , \3922 );
nor \U$11835 ( \12178 , \12175 , \12177 );
not \U$11836 ( \12179 , \2935 );
and \U$11837 ( \12180 , \3254 , RI986e800_25);
and \U$11838 ( \12181 , RI986ee90_39, \3252 );
nor \U$11839 ( \12182 , \12180 , \12181 );
not \U$11840 ( \12183 , \12182 );
or \U$11841 ( \12184 , \12179 , \12183 );
or \U$11842 ( \12185 , \12182 , \3406 );
nand \U$11843 ( \12186 , \12184 , \12185 );
xor \U$11844 ( \12187 , \12178 , \12186 );
not \U$11845 ( \12188 , \3918 );
and \U$11846 ( \12189 , \3683 , RI986eda0_37);
and \U$11847 ( \12190 , RI986ebc0_33, \3681 );
nor \U$11848 ( \12191 , \12189 , \12190 );
not \U$11849 ( \12192 , \12191 );
or \U$11850 ( \12193 , \12188 , \12192 );
or \U$11851 ( \12194 , \12191 , \3918 );
nand \U$11852 ( \12195 , \12193 , \12194 );
and \U$11853 ( \12196 , \12187 , \12195 );
and \U$11854 ( \12197 , \12178 , \12186 );
or \U$11855 ( \12198 , \12196 , \12197 );
and \U$11856 ( \12199 , \2464 , RI986e9e0_29);
and \U$11857 ( \12200 , RI986e8f0_27, \2462 );
nor \U$11858 ( \12201 , \12199 , \12200 );
and \U$11859 ( \12202 , \12201 , \2468 );
not \U$11860 ( \12203 , \12201 );
and \U$11861 ( \12204 , \12203 , \2263 );
nor \U$11862 ( \12205 , \12202 , \12204 );
not \U$11863 ( \12206 , \2034 );
and \U$11864 ( \12207 , \2042 , RI98717d0_127);
and \U$11865 ( \12208 , RI9871500_121, \2040 );
nor \U$11866 ( \12209 , \12207 , \12208 );
not \U$11867 ( \12210 , \12209 );
or \U$11868 ( \12211 , \12206 , \12210 );
or \U$11869 ( \12212 , \12209 , \1462 );
nand \U$11870 ( \12213 , \12211 , \12212 );
xor \U$11871 ( \12214 , \12205 , \12213 );
and \U$11872 ( \12215 , \2274 , RI98715f0_123);
and \U$11873 ( \12216 , RI986ead0_31, \2272 );
nor \U$11874 ( \12217 , \12215 , \12216 );
and \U$11875 ( \12218 , \12217 , \2030 );
not \U$11876 ( \12219 , \12217 );
and \U$11877 ( \12220 , \12219 , \2031 );
nor \U$11878 ( \12221 , \12218 , \12220 );
and \U$11879 ( \12222 , \12214 , \12221 );
and \U$11880 ( \12223 , \12205 , \12213 );
or \U$11881 ( \12224 , \12222 , \12223 );
xor \U$11882 ( \12225 , \12198 , \12224 );
and \U$11883 ( \12226 , \5881 , RI986e440_17);
and \U$11884 ( \12227 , RI986e710_23, \5879 );
nor \U$11885 ( \12228 , \12226 , \12227 );
and \U$11886 ( \12229 , \12228 , \5594 );
not \U$11887 ( \12230 , \12228 );
and \U$11888 ( \12231 , \12230 , \5885 );
nor \U$11889 ( \12232 , \12229 , \12231 );
not \U$11890 ( \12233 , \4519 );
and \U$11891 ( \12234 , \4710 , RI986ef80_41);
and \U$11892 ( \12235 , RI986f250_47, \4708 );
nor \U$11893 ( \12236 , \12234 , \12235 );
not \U$11894 ( \12237 , \12236 );
or \U$11895 ( \12238 , \12233 , \12237 );
or \U$11896 ( \12239 , \12236 , \4519 );
nand \U$11897 ( \12240 , \12238 , \12239 );
xor \U$11898 ( \12241 , \12232 , \12240 );
and \U$11899 ( \12242 , \5318 , RI986f160_45);
and \U$11900 ( \12243 , RI986e530_19, \5316 );
nor \U$11901 ( \12244 , \12242 , \12243 );
and \U$11902 ( \12245 , \12244 , \5052 );
not \U$11903 ( \12246 , \12244 );
and \U$11904 ( \12247 , \12246 , \5322 );
nor \U$11905 ( \12248 , \12245 , \12247 );
and \U$11906 ( \12249 , \12241 , \12248 );
and \U$11907 ( \12250 , \12232 , \12240 );
or \U$11908 ( \12251 , \12249 , \12250 );
and \U$11909 ( \12252 , \12225 , \12251 );
and \U$11910 ( \12253 , \12198 , \12224 );
or \U$11911 ( \12254 , \12252 , \12253 );
and \U$11912 ( \12255 , \6453 , RI986e620_21);
and \U$11913 ( \12256 , RI986f7f0_59, \6451 );
nor \U$11914 ( \12257 , \12255 , \12256 );
and \U$11915 ( \12258 , \12257 , \6190 );
not \U$11916 ( \12259 , \12257 );
and \U$11917 ( \12260 , \12259 , \6180 );
nor \U$11918 ( \12261 , \12258 , \12260 );
and \U$11919 ( \12262 , \7079 , RI986f700_57);
and \U$11920 ( \12263 , RI986f9d0_63, \7077 );
nor \U$11921 ( \12264 , \12262 , \12263 );
and \U$11922 ( \12265 , \12264 , \6710 );
not \U$11923 ( \12266 , \12264 );
and \U$11924 ( \12267 , \12266 , \6709 );
nor \U$11925 ( \12268 , \12265 , \12267 );
xor \U$11926 ( \12269 , \12261 , \12268 );
and \U$11927 ( \12270 , \7729 , RI986f8e0_61);
and \U$11928 ( \12271 , RI986f430_51, \7727 );
nor \U$11929 ( \12272 , \12270 , \12271 );
and \U$11930 ( \12273 , \12272 , \7480 );
not \U$11931 ( \12274 , \12272 );
and \U$11932 ( \12275 , \12274 , \7733 );
nor \U$11933 ( \12276 , \12273 , \12275 );
and \U$11934 ( \12277 , \12269 , \12276 );
and \U$11935 ( \12278 , \12261 , \12268 );
or \U$11936 ( \12279 , \12277 , \12278 );
and \U$11937 ( \12280 , \10424 , RI986dcc0_1);
and \U$11938 ( \12281 , RI986e170_11, \10422 );
nor \U$11939 ( \12282 , \12280 , \12281 );
and \U$11940 ( \12283 , \12282 , \9840 );
not \U$11941 ( \12284 , \12282 );
and \U$11942 ( \12285 , \12284 , \10428 );
nor \U$11943 ( \12286 , \12283 , \12285 );
and \U$11944 ( \12287 , RI9873210_183, RI9873300_185);
not \U$11945 ( \12288 , RI9873288_184);
and \U$11946 ( \12289 , \12288 , RI9873300_185);
nor \U$11947 ( \12290 , \12288 , RI9873300_185);
or \U$11948 ( \12291 , \12289 , \12290 );
nor \U$11949 ( \12292 , RI9873210_183, RI9873300_185);
nor \U$11950 ( \12293 , \12287 , \12291 , \12292 );
nand \U$11951 ( \12294 , RI986e350_15, \12293 );
and \U$11952 ( \12295 , \12294 , \11687 );
not \U$11953 ( \12296 , \12294 );
and \U$11954 ( \12297 , \12296 , \11686 );
nor \U$11955 ( \12298 , \12295 , \12297 );
xor \U$11956 ( \12299 , \12286 , \12298 );
and \U$11957 ( \12300 , \11696 , RI986e080_9);
and \U$11958 ( \12301 , RI986e260_13, \11694 );
nor \U$11959 ( \12302 , \12300 , \12301 );
and \U$11960 ( \12303 , \12302 , \10965 );
not \U$11961 ( \12304 , \12302 );
and \U$11962 ( \12305 , \12304 , \11702 );
nor \U$11963 ( \12306 , \12303 , \12305 );
and \U$11964 ( \12307 , \12299 , \12306 );
and \U$11965 ( \12308 , \12286 , \12298 );
or \U$11966 ( \12309 , \12307 , \12308 );
xor \U$11967 ( \12310 , \12279 , \12309 );
and \U$11968 ( \12311 , \8486 , RI986f340_49);
and \U$11969 ( \12312 , RI986f520_53, \8484 );
nor \U$11970 ( \12313 , \12311 , \12312 );
and \U$11971 ( \12314 , \12313 , \8050 );
not \U$11972 ( \12315 , \12313 );
and \U$11973 ( \12316 , \12315 , \8051 );
nor \U$11974 ( \12317 , \12314 , \12316 );
and \U$11975 ( \12318 , \9237 , RI986f610_55);
and \U$11976 ( \12319 , RI986df90_7, \9235 );
nor \U$11977 ( \12320 , \12318 , \12319 );
and \U$11978 ( \12321 , \12320 , \9241 );
not \U$11979 ( \12322 , \12320 );
and \U$11980 ( \12323 , \12322 , \8836 );
nor \U$11981 ( \12324 , \12321 , \12323 );
xor \U$11982 ( \12325 , \12317 , \12324 );
and \U$11983 ( \12326 , \9505 , RI986dea0_5);
and \U$11984 ( \12327 , RI986ddb0_3, \9503 );
nor \U$11985 ( \12328 , \12326 , \12327 );
and \U$11986 ( \12329 , \12328 , \9510 );
not \U$11987 ( \12330 , \12328 );
and \U$11988 ( \12331 , \12330 , \9513 );
nor \U$11989 ( \12332 , \12329 , \12331 );
and \U$11990 ( \12333 , \12325 , \12332 );
and \U$11991 ( \12334 , \12317 , \12324 );
or \U$11992 ( \12335 , \12333 , \12334 );
and \U$11993 ( \12336 , \12310 , \12335 );
and \U$11994 ( \12337 , \12279 , \12309 );
or \U$11995 ( \12338 , \12336 , \12337 );
xor \U$11996 ( \12339 , \12254 , \12338 );
not \U$11997 ( \12340 , \454 );
and \U$11998 ( \12341 , \465 , RI9870ab0_99);
and \U$11999 ( \12342 , RI9870d80_105, \463 );
nor \U$12000 ( \12343 , \12341 , \12342 );
not \U$12001 ( \12344 , \12343 );
or \U$12002 ( \12345 , \12340 , \12344 );
or \U$12003 ( \12346 , \12343 , \454 );
nand \U$12004 ( \12347 , \12345 , \12346 );
and \U$12005 ( \12348 , \776 , RI9870ba0_101);
and \U$12006 ( \12349 , RI9871050_111, \774 );
nor \U$12007 ( \12350 , \12348 , \12349 );
and \U$12008 ( \12351 , \12350 , \474 );
not \U$12009 ( \12352 , \12350 );
and \U$12010 ( \12353 , \12352 , \451 );
nor \U$12011 ( \12354 , \12351 , \12353 );
xor \U$12012 ( \12355 , \12347 , \12354 );
and \U$12013 ( \12356 , \438 , RI98709c0_97);
and \U$12014 ( \12357 , RI9870e70_107, \436 );
nor \U$12015 ( \12358 , \12356 , \12357 );
and \U$12016 ( \12359 , \12358 , \444 );
not \U$12017 ( \12360 , \12358 );
and \U$12018 ( \12361 , \12360 , \443 );
nor \U$12019 ( \12362 , \12359 , \12361 );
and \U$12020 ( \12363 , \12355 , \12362 );
and \U$12021 ( \12364 , \12347 , \12354 );
or \U$12022 ( \12365 , \12363 , \12364 );
not \U$12023 ( \12366 , \365 );
and \U$12024 ( \12367 , \376 , RI9870150_79);
and \U$12025 ( \12368 , RI9870f60_109, \374 );
nor \U$12026 ( \12369 , \12367 , \12368 );
not \U$12027 ( \12370 , \12369 );
or \U$12028 ( \12371 , \12366 , \12370 );
or \U$12029 ( \12372 , \12369 , \367 );
nand \U$12030 ( \12373 , \12371 , \12372 );
not \U$12031 ( \12374 , \487 );
and \U$12032 ( \12375 , \395 , RI986fe80_73);
and \U$12033 ( \12376 , RI9870060_77, \393 );
nor \U$12034 ( \12377 , \12375 , \12376 );
not \U$12035 ( \12378 , \12377 );
or \U$12036 ( \12379 , \12374 , \12378 );
or \U$12037 ( \12380 , \12377 , \386 );
nand \U$12038 ( \12381 , \12379 , \12380 );
xor \U$12039 ( \12382 , \12373 , \12381 );
not \U$12040 ( \12383 , \345 );
and \U$12041 ( \12384 , \354 , RI986fca0_69);
and \U$12042 ( \12385 , RI986ff70_75, \352 );
nor \U$12043 ( \12386 , \12384 , \12385 );
not \U$12044 ( \12387 , \12386 );
or \U$12045 ( \12388 , \12383 , \12387 );
or \U$12046 ( \12389 , \12386 , \345 );
nand \U$12047 ( \12390 , \12388 , \12389 );
and \U$12048 ( \12391 , \12382 , \12390 );
and \U$12049 ( \12392 , \12373 , \12381 );
or \U$12050 ( \12393 , \12391 , \12392 );
xor \U$12051 ( \12394 , \12365 , \12393 );
and \U$12052 ( \12395 , \1311 , RI9871410_119);
and \U$12053 ( \12396 , RI98716e0_125, \1309 );
nor \U$12054 ( \12397 , \12395 , \12396 );
and \U$12055 ( \12398 , \12397 , \1458 );
not \U$12056 ( \12399 , \12397 );
and \U$12057 ( \12400 , \12399 , \1318 );
nor \U$12058 ( \12401 , \12398 , \12400 );
not \U$12059 ( \12402 , \1128 );
and \U$12060 ( \12403 , \1293 , RI9870c90_103);
and \U$12061 ( \12404 , RI9871230_115, \1291 );
nor \U$12062 ( \12405 , \12403 , \12404 );
not \U$12063 ( \12406 , \12405 );
or \U$12064 ( \12407 , \12402 , \12406 );
or \U$12065 ( \12408 , \12405 , \1128 );
nand \U$12066 ( \12409 , \12407 , \12408 );
xor \U$12067 ( \12410 , \12401 , \12409 );
and \U$12068 ( \12411 , \1329 , RI9871140_113);
and \U$12069 ( \12412 , RI9871320_117, \1327 );
nor \U$12070 ( \12413 , \12411 , \12412 );
and \U$12071 ( \12414 , \12413 , \1336 );
not \U$12072 ( \12415 , \12413 );
and \U$12073 ( \12416 , \12415 , \1337 );
nor \U$12074 ( \12417 , \12414 , \12416 );
and \U$12075 ( \12418 , \12410 , \12417 );
and \U$12076 ( \12419 , \12401 , \12409 );
or \U$12077 ( \12420 , \12418 , \12419 );
and \U$12078 ( \12421 , \12394 , \12420 );
and \U$12079 ( \12422 , \12365 , \12393 );
or \U$12080 ( \12423 , \12421 , \12422 );
xor \U$12081 ( \12424 , \12339 , \12423 );
xor \U$12082 ( \12425 , \12171 , \12424 );
xor \U$12083 ( \12426 , \11863 , \11870 );
xor \U$12084 ( \12427 , \12426 , \11878 );
xor \U$12085 ( \12428 , \11893 , \11898 );
xor \U$12086 ( \12429 , \12428 , \11906 );
xor \U$12087 ( \12430 , \11684 , \11687 );
xor \U$12088 ( \12431 , \12430 , \11704 );
xor \U$12089 ( \12432 , \11659 , \11666 );
xor \U$12090 ( \12433 , \12432 , \11674 );
and \U$12091 ( \12434 , \12431 , \12433 );
xor \U$12092 ( \12435 , \11715 , \11722 );
xor \U$12093 ( \12436 , \12435 , \11730 );
xor \U$12094 ( \12437 , \11659 , \11666 );
xor \U$12095 ( \12438 , \12437 , \11674 );
and \U$12096 ( \12439 , \12436 , \12438 );
and \U$12097 ( \12440 , \12431 , \12436 );
or \U$12098 ( \12441 , \12434 , \12439 , \12440 );
xor \U$12099 ( \12442 , \12429 , \12441 );
xor \U$12100 ( \12443 , \12427 , \12442 );
and \U$12101 ( \12444 , \12425 , \12443 );
and \U$12102 ( \12445 , \12171 , \12424 );
or \U$12103 ( \12446 , \12444 , \12445 );
xor \U$12104 ( \12447 , \12178 , \12186 );
xor \U$12105 ( \12448 , \12447 , \12195 );
xor \U$12106 ( \12449 , \12261 , \12268 );
xor \U$12107 ( \12450 , \12449 , \12276 );
and \U$12108 ( \12451 , \12448 , \12450 );
xor \U$12109 ( \12452 , \12232 , \12240 );
xor \U$12110 ( \12453 , \12452 , \12248 );
xor \U$12111 ( \12454 , \12261 , \12268 );
xor \U$12112 ( \12455 , \12454 , \12276 );
and \U$12113 ( \12456 , \12453 , \12455 );
and \U$12114 ( \12457 , \12448 , \12453 );
or \U$12115 ( \12458 , \12451 , \12456 , \12457 );
not \U$12116 ( \12459 , \345 );
and \U$12117 ( \12460 , \354 , RI986fd90_71);
and \U$12118 ( \12461 , RI986fca0_69, \352 );
nor \U$12119 ( \12462 , \12460 , \12461 );
not \U$12120 ( \12463 , \12462 );
or \U$12121 ( \12464 , \12459 , \12463 );
or \U$12122 ( \12465 , \12462 , \345 );
nand \U$12123 ( \12466 , \12464 , \12465 );
not \U$12124 ( \12467 , RI98707e0_93);
nor \U$12125 ( \12468 , \12467 , \407 );
xor \U$12126 ( \12469 , \12466 , \12468 );
and \U$12127 ( \12470 , \416 , RI986fac0_65);
and \U$12128 ( \12471 , RI986fbb0_67, \414 );
nor \U$12129 ( \12472 , \12470 , \12471 );
and \U$12130 ( \12473 , \12472 , \422 );
not \U$12131 ( \12474 , \12472 );
and \U$12132 ( \12475 , \12474 , \421 );
nor \U$12133 ( \12476 , \12473 , \12475 );
and \U$12134 ( \12477 , \12469 , \12476 );
and \U$12135 ( \12478 , \12466 , \12468 );
or \U$12136 ( \12479 , \12477 , \12478 );
or \U$12137 ( \12480 , \12155 , \12148 );
nand \U$12138 ( \12481 , \12480 , \12156 );
xor \U$12139 ( \12482 , \12479 , \12481 );
xor \U$12140 ( \12483 , \12373 , \12381 );
xor \U$12141 ( \12484 , \12483 , \12390 );
and \U$12142 ( \12485 , \12482 , \12484 );
and \U$12143 ( \12486 , \12479 , \12481 );
or \U$12144 ( \12487 , \12485 , \12486 );
xor \U$12145 ( \12488 , \12458 , \12487 );
xor \U$12146 ( \12489 , \12347 , \12354 );
xor \U$12147 ( \12490 , \12489 , \12362 );
xor \U$12148 ( \12491 , \12401 , \12409 );
xor \U$12149 ( \12492 , \12491 , \12417 );
xor \U$12150 ( \12493 , \12490 , \12492 );
xor \U$12151 ( \12494 , \12205 , \12213 );
xor \U$12152 ( \12495 , \12494 , \12221 );
and \U$12153 ( \12496 , \12493 , \12495 );
and \U$12154 ( \12497 , \12490 , \12492 );
or \U$12155 ( \12498 , \12496 , \12497 );
and \U$12156 ( \12499 , \12488 , \12498 );
and \U$12157 ( \12500 , \12458 , \12487 );
or \U$12158 ( \12501 , \12499 , \12500 );
not \U$12159 ( \12502 , \454 );
and \U$12160 ( \12503 , \465 , RI9870f60_109);
and \U$12161 ( \12504 , RI9870ab0_99, \463 );
nor \U$12162 ( \12505 , \12503 , \12504 );
not \U$12163 ( \12506 , \12505 );
or \U$12164 ( \12507 , \12502 , \12506 );
or \U$12165 ( \12508 , \12505 , \456 );
nand \U$12166 ( \12509 , \12507 , \12508 );
not \U$12167 ( \12510 , \367 );
and \U$12168 ( \12511 , \376 , RI9870060_77);
and \U$12169 ( \12512 , RI9870150_79, \374 );
nor \U$12170 ( \12513 , \12511 , \12512 );
not \U$12171 ( \12514 , \12513 );
or \U$12172 ( \12515 , \12510 , \12514 );
or \U$12173 ( \12516 , \12513 , \367 );
nand \U$12174 ( \12517 , \12515 , \12516 );
xor \U$12175 ( \12518 , \12509 , \12517 );
not \U$12176 ( \12519 , \487 );
and \U$12177 ( \12520 , \395 , RI986ff70_75);
and \U$12178 ( \12521 , RI986fe80_73, \393 );
nor \U$12179 ( \12522 , \12520 , \12521 );
not \U$12180 ( \12523 , \12522 );
or \U$12181 ( \12524 , \12519 , \12523 );
or \U$12182 ( \12525 , \12522 , \487 );
nand \U$12183 ( \12526 , \12524 , \12525 );
and \U$12184 ( \12527 , \12518 , \12526 );
and \U$12185 ( \12528 , \12509 , \12517 );
or \U$12186 ( \12529 , \12527 , \12528 );
and \U$12187 ( \12530 , \776 , RI9870e70_107);
and \U$12188 ( \12531 , RI9870ba0_101, \774 );
nor \U$12189 ( \12532 , \12530 , \12531 );
and \U$12190 ( \12533 , \12532 , \474 );
not \U$12191 ( \12534 , \12532 );
and \U$12192 ( \12535 , \12534 , \451 );
nor \U$12193 ( \12536 , \12533 , \12535 );
and \U$12194 ( \12537 , \438 , RI9870d80_105);
and \U$12195 ( \12538 , RI98709c0_97, \436 );
nor \U$12196 ( \12539 , \12537 , \12538 );
and \U$12197 ( \12540 , \12539 , \444 );
not \U$12198 ( \12541 , \12539 );
and \U$12199 ( \12542 , \12541 , \443 );
nor \U$12200 ( \12543 , \12540 , \12542 );
xor \U$12201 ( \12544 , \12536 , \12543 );
not \U$12202 ( \12545 , \1128 );
and \U$12203 ( \12546 , \1293 , RI9871050_111);
and \U$12204 ( \12547 , RI9870c90_103, \1291 );
nor \U$12205 ( \12548 , \12546 , \12547 );
not \U$12206 ( \12549 , \12548 );
or \U$12207 ( \12550 , \12545 , \12549 );
or \U$12208 ( \12551 , \12548 , \1301 );
nand \U$12209 ( \12552 , \12550 , \12551 );
and \U$12210 ( \12553 , \12544 , \12552 );
and \U$12211 ( \12554 , \12536 , \12543 );
or \U$12212 ( \12555 , \12553 , \12554 );
xor \U$12213 ( \12556 , \12529 , \12555 );
and \U$12214 ( \12557 , \1329 , RI9871230_115);
and \U$12215 ( \12558 , RI9871140_113, \1327 );
nor \U$12216 ( \12559 , \12557 , \12558 );
and \U$12217 ( \12560 , \12559 , \1336 );
not \U$12218 ( \12561 , \12559 );
and \U$12219 ( \12562 , \12561 , \1337 );
nor \U$12220 ( \12563 , \12560 , \12562 );
and \U$12221 ( \12564 , \1311 , RI9871320_117);
and \U$12222 ( \12565 , RI9871410_119, \1309 );
nor \U$12223 ( \12566 , \12564 , \12565 );
and \U$12224 ( \12567 , \12566 , \1319 );
not \U$12225 ( \12568 , \12566 );
and \U$12226 ( \12569 , \12568 , \1318 );
nor \U$12227 ( \12570 , \12567 , \12569 );
xor \U$12228 ( \12571 , \12563 , \12570 );
not \U$12229 ( \12572 , \1462 );
and \U$12230 ( \12573 , \2042 , RI98716e0_125);
and \U$12231 ( \12574 , RI98717d0_127, \2040 );
nor \U$12232 ( \12575 , \12573 , \12574 );
not \U$12233 ( \12576 , \12575 );
or \U$12234 ( \12577 , \12572 , \12576 );
or \U$12235 ( \12578 , \12575 , \1462 );
nand \U$12236 ( \12579 , \12577 , \12578 );
and \U$12237 ( \12580 , \12571 , \12579 );
and \U$12238 ( \12581 , \12563 , \12570 );
or \U$12239 ( \12582 , \12580 , \12581 );
and \U$12240 ( \12583 , \12556 , \12582 );
and \U$12241 ( \12584 , \12529 , \12555 );
or \U$12242 ( \12585 , \12583 , \12584 );
and \U$12243 ( \12586 , \9505 , RI986df90_7);
and \U$12244 ( \12587 , RI986dea0_5, \9503 );
nor \U$12245 ( \12588 , \12586 , \12587 );
and \U$12246 ( \12589 , \12588 , \9513 );
not \U$12247 ( \12590 , \12588 );
and \U$12248 ( \12591 , \12590 , \9510 );
nor \U$12249 ( \12592 , \12589 , \12591 );
and \U$12250 ( \12593 , \10424 , RI986ddb0_3);
and \U$12251 ( \12594 , RI986dcc0_1, \10422 );
nor \U$12252 ( \12595 , \12593 , \12594 );
and \U$12253 ( \12596 , \12595 , \10428 );
not \U$12254 ( \12597 , \12595 );
and \U$12255 ( \12598 , \12597 , \9840 );
nor \U$12256 ( \12599 , \12596 , \12598 );
xor \U$12257 ( \12600 , \12592 , \12599 );
and \U$12258 ( \12601 , \9237 , RI986f520_53);
and \U$12259 ( \12602 , RI986f610_55, \9235 );
nor \U$12260 ( \12603 , \12601 , \12602 );
and \U$12261 ( \12604 , \12603 , \8836 );
not \U$12262 ( \12605 , \12603 );
and \U$12263 ( \12606 , \12605 , \9241 );
nor \U$12264 ( \12607 , \12604 , \12606 );
and \U$12265 ( \12608 , \12600 , \12607 );
and \U$12266 ( \12609 , \12592 , \12599 );
nor \U$12267 ( \12610 , \12608 , \12609 );
and \U$12268 ( \12611 , \11696 , RI986e170_11);
and \U$12269 ( \12612 , RI986e080_9, \11694 );
nor \U$12270 ( \12613 , \12611 , \12612 );
and \U$12271 ( \12614 , \12613 , \11702 );
not \U$12272 ( \12615 , \12613 );
and \U$12273 ( \12616 , \12615 , \10965 );
nor \U$12274 ( \12617 , \12614 , \12616 );
nand \U$12275 ( \12618 , RI98733f0_187, RI9873378_186);
and \U$12276 ( \12619 , \12618 , RI9873288_184);
or \U$12277 ( \12620 , \12617 , \12619 );
not \U$12278 ( \12621 , \12619 );
not \U$12279 ( \12622 , \12617 );
or \U$12280 ( \12623 , \12621 , \12622 );
and \U$12281 ( \12624 , \12293 , RI986e260_13);
and \U$12282 ( \12625 , RI986e350_15, \12291 );
nor \U$12283 ( \12626 , \12624 , \12625 );
and \U$12284 ( \12627 , \12626 , \11687 );
not \U$12285 ( \12628 , \12626 );
and \U$12286 ( \12629 , \12628 , \11686 );
nor \U$12287 ( \12630 , \12627 , \12629 );
nand \U$12288 ( \12631 , \12623 , \12630 );
nand \U$12289 ( \12632 , \12620 , \12631 );
xor \U$12290 ( \12633 , \12610 , \12632 );
and \U$12291 ( \12634 , \8486 , RI986f430_51);
and \U$12292 ( \12635 , RI986f340_49, \8484 );
nor \U$12293 ( \12636 , \12634 , \12635 );
and \U$12294 ( \12637 , \12636 , \8050 );
not \U$12295 ( \12638 , \12636 );
and \U$12296 ( \12639 , \12638 , \8051 );
nor \U$12297 ( \12640 , \12637 , \12639 );
and \U$12298 ( \12641 , \7079 , RI986f7f0_59);
and \U$12299 ( \12642 , RI986f700_57, \7077 );
nor \U$12300 ( \12643 , \12641 , \12642 );
and \U$12301 ( \12644 , \12643 , \6710 );
not \U$12302 ( \12645 , \12643 );
and \U$12303 ( \12646 , \12645 , \6709 );
nor \U$12304 ( \12647 , \12644 , \12646 );
xor \U$12305 ( \12648 , \12640 , \12647 );
and \U$12306 ( \12649 , \7729 , RI986f9d0_63);
and \U$12307 ( \12650 , RI986f8e0_61, \7727 );
nor \U$12308 ( \12651 , \12649 , \12650 );
and \U$12309 ( \12652 , \12651 , \7480 );
not \U$12310 ( \12653 , \12651 );
and \U$12311 ( \12654 , \12653 , \7733 );
nor \U$12312 ( \12655 , \12652 , \12654 );
and \U$12313 ( \12656 , \12648 , \12655 );
and \U$12314 ( \12657 , \12640 , \12647 );
or \U$12315 ( \12658 , \12656 , \12657 );
and \U$12316 ( \12659 , \12633 , \12658 );
and \U$12317 ( \12660 , \12610 , \12632 );
or \U$12318 ( \12661 , \12659 , \12660 );
xor \U$12319 ( \12662 , \12585 , \12661 );
not \U$12320 ( \12663 , \4521 );
and \U$12321 ( \12664 , \4710 , RI986f070_43);
and \U$12322 ( \12665 , RI986ef80_41, \4708 );
nor \U$12323 ( \12666 , \12664 , \12665 );
not \U$12324 ( \12667 , \12666 );
or \U$12325 ( \12668 , \12663 , \12667 );
or \U$12326 ( \12669 , \12666 , \4519 );
nand \U$12327 ( \12670 , \12668 , \12669 );
not \U$12328 ( \12671 , \3918 );
and \U$12329 ( \12672 , \3683 , RI986ee90_39);
and \U$12330 ( \12673 , RI986eda0_37, \3681 );
nor \U$12331 ( \12674 , \12672 , \12673 );
not \U$12332 ( \12675 , \12674 );
or \U$12333 ( \12676 , \12671 , \12675 );
or \U$12334 ( \12677 , \12674 , \3918 );
nand \U$12335 ( \12678 , \12676 , \12677 );
xor \U$12336 ( \12679 , \12670 , \12678 );
and \U$12337 ( \12680 , \4203 , RI986ebc0_33);
and \U$12338 ( \12681 , RI986ecb0_35, \4201 );
nor \U$12339 ( \12682 , \12680 , \12681 );
and \U$12340 ( \12683 , \12682 , \4207 );
not \U$12341 ( \12684 , \12682 );
and \U$12342 ( \12685 , \12684 , \3922 );
nor \U$12343 ( \12686 , \12683 , \12685 );
and \U$12344 ( \12687 , \12679 , \12686 );
and \U$12345 ( \12688 , \12670 , \12678 );
or \U$12346 ( \12689 , \12687 , \12688 );
not \U$12347 ( \12690 , \2935 );
and \U$12348 ( \12691 , \3254 , RI986e8f0_27);
and \U$12349 ( \12692 , RI986e800_25, \3252 );
nor \U$12350 ( \12693 , \12691 , \12692 );
not \U$12351 ( \12694 , \12693 );
or \U$12352 ( \12695 , \12690 , \12694 );
or \U$12353 ( \12696 , \12693 , \2935 );
nand \U$12354 ( \12697 , \12695 , \12696 );
and \U$12355 ( \12698 , \2274 , RI9871500_121);
and \U$12356 ( \12699 , RI98715f0_123, \2272 );
nor \U$12357 ( \12700 , \12698 , \12699 );
and \U$12358 ( \12701 , \12700 , \2030 );
not \U$12359 ( \12702 , \12700 );
and \U$12360 ( \12703 , \12702 , \2031 );
nor \U$12361 ( \12704 , \12701 , \12703 );
xor \U$12362 ( \12705 , \12697 , \12704 );
and \U$12363 ( \12706 , \2464 , RI986ead0_31);
and \U$12364 ( \12707 , RI986e9e0_29, \2462 );
nor \U$12365 ( \12708 , \12706 , \12707 );
and \U$12366 ( \12709 , \12708 , \2468 );
not \U$12367 ( \12710 , \12708 );
and \U$12368 ( \12711 , \12710 , \2263 );
nor \U$12369 ( \12712 , \12709 , \12711 );
and \U$12370 ( \12713 , \12705 , \12712 );
and \U$12371 ( \12714 , \12697 , \12704 );
or \U$12372 ( \12715 , \12713 , \12714 );
xor \U$12373 ( \12716 , \12689 , \12715 );
and \U$12374 ( \12717 , \6453 , RI986e710_23);
and \U$12375 ( \12718 , RI986e620_21, \6451 );
nor \U$12376 ( \12719 , \12717 , \12718 );
and \U$12377 ( \12720 , \12719 , \6190 );
not \U$12378 ( \12721 , \12719 );
and \U$12379 ( \12722 , \12721 , \6705 );
nor \U$12380 ( \12723 , \12720 , \12722 );
and \U$12381 ( \12724 , \5318 , RI986f250_47);
and \U$12382 ( \12725 , RI986f160_45, \5316 );
nor \U$12383 ( \12726 , \12724 , \12725 );
and \U$12384 ( \12727 , \12726 , \5052 );
not \U$12385 ( \12728 , \12726 );
and \U$12386 ( \12729 , \12728 , \5322 );
nor \U$12387 ( \12730 , \12727 , \12729 );
xor \U$12388 ( \12731 , \12723 , \12730 );
and \U$12389 ( \12732 , \5881 , RI986e530_19);
and \U$12390 ( \12733 , RI986e440_17, \5879 );
nor \U$12391 ( \12734 , \12732 , \12733 );
and \U$12392 ( \12735 , \12734 , \5594 );
not \U$12393 ( \12736 , \12734 );
and \U$12394 ( \12737 , \12736 , \5885 );
nor \U$12395 ( \12738 , \12735 , \12737 );
and \U$12396 ( \12739 , \12731 , \12738 );
and \U$12397 ( \12740 , \12723 , \12730 );
or \U$12398 ( \12741 , \12739 , \12740 );
and \U$12399 ( \12742 , \12716 , \12741 );
and \U$12400 ( \12743 , \12689 , \12715 );
or \U$12401 ( \12744 , \12742 , \12743 );
and \U$12402 ( \12745 , \12662 , \12744 );
and \U$12403 ( \12746 , \12585 , \12661 );
or \U$12404 ( \12747 , \12745 , \12746 );
xor \U$12405 ( \12748 , \12501 , \12747 );
xor \U$12406 ( \12749 , \11659 , \11666 );
xor \U$12407 ( \12750 , \12749 , \11674 );
xor \U$12408 ( \12751 , \12431 , \12436 );
xor \U$12409 ( \12752 , \12750 , \12751 );
xor \U$12410 ( \12753 , \12162 , \12164 );
xor \U$12411 ( \12754 , \12753 , \12167 );
and \U$12412 ( \12755 , \12752 , \12754 );
xor \U$12413 ( \12756 , \11576 , \11583 );
xor \U$12414 ( \12757 , \12756 , \11591 );
xor \U$12415 ( \12758 , \12127 , \12132 );
xor \U$12416 ( \12759 , \12757 , \12758 );
xor \U$12417 ( \12760 , \12162 , \12164 );
xor \U$12418 ( \12761 , \12760 , \12167 );
and \U$12419 ( \12762 , \12759 , \12761 );
and \U$12420 ( \12763 , \12752 , \12759 );
or \U$12421 ( \12764 , \12755 , \12762 , \12763 );
and \U$12422 ( \12765 , \12748 , \12764 );
and \U$12423 ( \12766 , \12501 , \12747 );
or \U$12424 ( \12767 , \12765 , \12766 );
xor \U$12425 ( \12768 , \12446 , \12767 );
xor \U$12426 ( \12769 , \12144 , \12146 );
xor \U$12427 ( \12770 , \12769 , \12156 );
xor \U$12428 ( \12771 , \12365 , \12393 );
xor \U$12429 ( \12772 , \12771 , \12420 );
and \U$12430 ( \12773 , \12770 , \12772 );
xor \U$12431 ( \12774 , \12198 , \12224 );
xor \U$12432 ( \12775 , \12774 , \12251 );
xor \U$12433 ( \12776 , \12365 , \12393 );
xor \U$12434 ( \12777 , \12776 , \12420 );
and \U$12435 ( \12778 , \12775 , \12777 );
and \U$12436 ( \12779 , \12770 , \12775 );
or \U$12437 ( \12780 , \12773 , \12778 , \12779 );
xor \U$12438 ( \12781 , \12081 , \12083 );
xor \U$12439 ( \12782 , \12781 , \12086 );
and \U$12440 ( \12783 , \12780 , \12782 );
xor \U$12441 ( \12784 , \11557 , \11559 );
xor \U$12442 ( \12785 , \12784 , \11562 );
xor \U$12443 ( \12786 , \12094 , \12101 );
xor \U$12444 ( \12787 , \12785 , \12786 );
xor \U$12445 ( \12788 , \12081 , \12083 );
xor \U$12446 ( \12789 , \12788 , \12086 );
and \U$12447 ( \12790 , \12787 , \12789 );
and \U$12448 ( \12791 , \12780 , \12787 );
or \U$12449 ( \12792 , \12783 , \12790 , \12791 );
and \U$12450 ( \12793 , \12768 , \12792 );
and \U$12451 ( \12794 , \12446 , \12767 );
or \U$12452 ( \12795 , \12793 , \12794 );
xor \U$12453 ( \12796 , \12125 , \12795 );
xor \U$12454 ( \12797 , \11495 , \11497 );
xor \U$12455 ( \12798 , \12797 , \11506 );
xor \U$12456 ( \12799 , \11568 , \11823 );
xor \U$12457 ( \12800 , \12799 , \11848 );
xor \U$12458 ( \12801 , \11926 , \11934 );
xor \U$12459 ( \12802 , \12801 , \11939 );
xor \U$12460 ( \12803 , \11918 , \11951 );
xor \U$12461 ( \12804 , \12802 , \12803 );
xor \U$12462 ( \12805 , \12800 , \12804 );
xor \U$12463 ( \12806 , \12798 , \12805 );
and \U$12464 ( \12807 , \12796 , \12806 );
and \U$12465 ( \12808 , \12125 , \12795 );
or \U$12466 ( \12809 , \12807 , \12808 );
xor \U$12467 ( \12810 , \11509 , \11851 );
xor \U$12468 ( \12811 , \12810 , \11956 );
xor \U$12469 ( \12812 , \12809 , \12811 );
xor \U$12470 ( \12813 , \11495 , \11497 );
xor \U$12471 ( \12814 , \12813 , \11506 );
and \U$12472 ( \12815 , \12800 , \12814 );
xor \U$12473 ( \12816 , \11495 , \11497 );
xor \U$12474 ( \12817 , \12816 , \11506 );
and \U$12475 ( \12818 , \12804 , \12817 );
and \U$12476 ( \12819 , \12800 , \12804 );
or \U$12477 ( \12820 , \12815 , \12818 , \12819 );
xor \U$12478 ( \12821 , \12089 , \12091 );
and \U$12479 ( \12822 , \12821 , \12106 );
and \U$12480 ( \12823 , \12089 , \12091 );
or \U$12481 ( \12824 , \12822 , \12823 );
xor \U$12482 ( \12825 , \12254 , \12338 );
and \U$12483 ( \12826 , \12825 , \12423 );
and \U$12484 ( \12827 , \12254 , \12338 );
or \U$12485 ( \12828 , \12826 , \12827 );
xor \U$12486 ( \12829 , \11863 , \11870 );
xor \U$12487 ( \12830 , \12829 , \11878 );
and \U$12488 ( \12831 , \12429 , \12830 );
xor \U$12489 ( \12832 , \11863 , \11870 );
xor \U$12490 ( \12833 , \12832 , \11878 );
and \U$12491 ( \12834 , \12441 , \12833 );
and \U$12492 ( \12835 , \12429 , \12441 );
or \U$12493 ( \12836 , \12831 , \12834 , \12835 );
xor \U$12494 ( \12837 , \12828 , \12836 );
xor \U$12495 ( \12838 , \12137 , \12159 );
and \U$12496 ( \12839 , \12838 , \12170 );
and \U$12497 ( \12840 , \12137 , \12159 );
or \U$12498 ( \12841 , \12839 , \12840 );
and \U$12499 ( \12842 , \12837 , \12841 );
and \U$12500 ( \12843 , \12828 , \12836 );
or \U$12501 ( \12844 , \12842 , \12843 );
xor \U$12502 ( \12845 , \12824 , \12844 );
xor \U$12503 ( \12846 , \11542 , \11554 );
xor \U$12504 ( \12847 , \12846 , \11565 );
and \U$12505 ( \12848 , \12114 , \12847 );
xor \U$12506 ( \12849 , \11542 , \11554 );
xor \U$12507 ( \12850 , \12849 , \11565 );
and \U$12508 ( \12851 , \12118 , \12850 );
and \U$12509 ( \12852 , \12114 , \12118 );
or \U$12510 ( \12853 , \12848 , \12851 , \12852 );
and \U$12511 ( \12854 , \12845 , \12853 );
and \U$12512 ( \12855 , \12824 , \12844 );
or \U$12513 ( \12856 , \12854 , \12855 );
xor \U$12514 ( \12857 , \12820 , \12856 );
xor \U$12515 ( \12858 , \11968 , \11972 );
xor \U$12516 ( \12859 , \12858 , \11981 );
xor \U$12517 ( \12860 , \11964 , \11999 );
xor \U$12518 ( \12861 , \12859 , \12860 );
xor \U$12519 ( \12862 , \12857 , \12861 );
and \U$12520 ( \12863 , \12812 , \12862 );
and \U$12521 ( \12864 , \12809 , \12811 );
or \U$12522 ( \12865 , \12863 , \12864 );
xor \U$12523 ( \12866 , \12820 , \12856 );
and \U$12524 ( \12867 , \12866 , \12861 );
and \U$12525 ( \12868 , \12820 , \12856 );
or \U$12526 ( \12869 , \12867 , \12868 );
xor \U$12527 ( \12870 , \12024 , \12025 );
xor \U$12528 ( \12871 , \12870 , \12034 );
xor \U$12529 ( \12872 , \12869 , \12871 );
xor \U$12530 ( \12873 , \11959 , \12004 );
xor \U$12531 ( \12874 , \12873 , \12014 );
xor \U$12532 ( \12875 , \12872 , \12874 );
and \U$12533 ( \12876 , \12865 , \12875 );
not \U$12534 ( \12877 , \12876 );
xor \U$12535 ( \12878 , \12869 , \12871 );
and \U$12536 ( \12879 , \12878 , \12874 );
and \U$12537 ( \12880 , \12869 , \12871 );
or \U$12538 ( \12881 , \12879 , \12880 );
xor \U$12539 ( \12882 , \12017 , \12019 );
xor \U$12540 ( \12883 , \12882 , \12051 );
xor \U$12541 ( \12884 , \12881 , \12883 );
not \U$12542 ( \12885 , \12884 );
or \U$12543 ( \12886 , \12877 , \12885 );
xor \U$12544 ( \12887 , \12446 , \12767 );
xor \U$12545 ( \12888 , \12887 , \12792 );
xor \U$12546 ( \12889 , \12089 , \12091 );
xor \U$12547 ( \12890 , \12889 , \12106 );
xor \U$12548 ( \12891 , \12079 , \12120 );
xor \U$12549 ( \12892 , \12890 , \12891 );
and \U$12550 ( \12893 , \12888 , \12892 );
xor \U$12551 ( \12894 , \12824 , \12844 );
xor \U$12552 ( \12895 , \12894 , \12853 );
xor \U$12553 ( \12896 , \12893 , \12895 );
xor \U$12554 ( \12897 , \12585 , \12661 );
xor \U$12555 ( \12898 , \12897 , \12744 );
xor \U$12556 ( \12899 , \12458 , \12487 );
xor \U$12557 ( \12900 , \12899 , \12498 );
and \U$12558 ( \12901 , \12898 , \12900 );
xor \U$12559 ( \12902 , \12162 , \12164 );
xor \U$12560 ( \12903 , \12902 , \12167 );
xor \U$12561 ( \12904 , \12752 , \12759 );
xor \U$12562 ( \12905 , \12903 , \12904 );
xor \U$12563 ( \12906 , \12458 , \12487 );
xor \U$12564 ( \12907 , \12906 , \12498 );
and \U$12565 ( \12908 , \12905 , \12907 );
and \U$12566 ( \12909 , \12898 , \12905 );
or \U$12567 ( \12910 , \12901 , \12908 , \12909 );
xor \U$12568 ( \12911 , \12317 , \12324 );
xor \U$12569 ( \12912 , \12911 , \12332 );
xor \U$12570 ( \12913 , \12286 , \12298 );
xor \U$12571 ( \12914 , \12913 , \12306 );
xor \U$12572 ( \12915 , \12912 , \12914 );
xor \U$12573 ( \12916 , \12261 , \12268 );
xor \U$12574 ( \12917 , \12916 , \12276 );
xor \U$12575 ( \12918 , \12448 , \12453 );
xor \U$12576 ( \12919 , \12917 , \12918 );
and \U$12577 ( \12920 , \12915 , \12919 );
and \U$12578 ( \12921 , \12912 , \12914 );
or \U$12579 ( \12922 , \12920 , \12921 );
not \U$12580 ( \12923 , \1128 );
and \U$12581 ( \12924 , \1293 , RI9870ba0_101);
and \U$12582 ( \12925 , RI9871050_111, \1291 );
nor \U$12583 ( \12926 , \12924 , \12925 );
not \U$12584 ( \12927 , \12926 );
or \U$12585 ( \12928 , \12923 , \12927 );
or \U$12586 ( \12929 , \12926 , \1128 );
nand \U$12587 ( \12930 , \12928 , \12929 );
and \U$12588 ( \12931 , \776 , RI98709c0_97);
and \U$12589 ( \12932 , RI9870e70_107, \774 );
nor \U$12590 ( \12933 , \12931 , \12932 );
and \U$12591 ( \12934 , \12933 , \474 );
not \U$12592 ( \12935 , \12933 );
and \U$12593 ( \12936 , \12935 , \451 );
nor \U$12594 ( \12937 , \12934 , \12936 );
xor \U$12595 ( \12938 , \12930 , \12937 );
and \U$12596 ( \12939 , \438 , RI9870ab0_99);
and \U$12597 ( \12940 , RI9870d80_105, \436 );
nor \U$12598 ( \12941 , \12939 , \12940 );
and \U$12599 ( \12942 , \12941 , \444 );
not \U$12600 ( \12943 , \12941 );
and \U$12601 ( \12944 , \12943 , \443 );
nor \U$12602 ( \12945 , \12942 , \12944 );
and \U$12603 ( \12946 , \12938 , \12945 );
and \U$12604 ( \12947 , \12930 , \12937 );
or \U$12605 ( \12948 , \12946 , \12947 );
not \U$12606 ( \12949 , \454 );
and \U$12607 ( \12950 , \465 , RI9870150_79);
and \U$12608 ( \12951 , RI9870f60_109, \463 );
nor \U$12609 ( \12952 , \12950 , \12951 );
not \U$12610 ( \12953 , \12952 );
or \U$12611 ( \12954 , \12949 , \12953 );
or \U$12612 ( \12955 , \12952 , \456 );
nand \U$12613 ( \12956 , \12954 , \12955 );
not \U$12614 ( \12957 , \367 );
and \U$12615 ( \12958 , \376 , RI986fe80_73);
and \U$12616 ( \12959 , RI9870060_77, \374 );
nor \U$12617 ( \12960 , \12958 , \12959 );
not \U$12618 ( \12961 , \12960 );
or \U$12619 ( \12962 , \12957 , \12961 );
or \U$12620 ( \12963 , \12960 , \365 );
nand \U$12621 ( \12964 , \12962 , \12963 );
xor \U$12622 ( \12965 , \12956 , \12964 );
not \U$12623 ( \12966 , \386 );
and \U$12624 ( \12967 , \395 , RI986fca0_69);
and \U$12625 ( \12968 , RI986ff70_75, \393 );
nor \U$12626 ( \12969 , \12967 , \12968 );
not \U$12627 ( \12970 , \12969 );
or \U$12628 ( \12971 , \12966 , \12970 );
or \U$12629 ( \12972 , \12969 , \487 );
nand \U$12630 ( \12973 , \12971 , \12972 );
and \U$12631 ( \12974 , \12965 , \12973 );
and \U$12632 ( \12975 , \12956 , \12964 );
or \U$12633 ( \12976 , \12974 , \12975 );
xor \U$12634 ( \12977 , \12948 , \12976 );
and \U$12635 ( \12978 , \1329 , RI9870c90_103);
and \U$12636 ( \12979 , RI9871230_115, \1327 );
nor \U$12637 ( \12980 , \12978 , \12979 );
and \U$12638 ( \12981 , \12980 , \1336 );
not \U$12639 ( \12982 , \12980 );
and \U$12640 ( \12983 , \12982 , \1337 );
nor \U$12641 ( \12984 , \12981 , \12983 );
and \U$12642 ( \12985 , \1311 , RI9871140_113);
and \U$12643 ( \12986 , RI9871320_117, \1309 );
nor \U$12644 ( \12987 , \12985 , \12986 );
and \U$12645 ( \12988 , \12987 , \1458 );
not \U$12646 ( \12989 , \12987 );
and \U$12647 ( \12990 , \12989 , \1318 );
nor \U$12648 ( \12991 , \12988 , \12990 );
xor \U$12649 ( \12992 , \12984 , \12991 );
not \U$12650 ( \12993 , \2034 );
and \U$12651 ( \12994 , \2042 , RI9871410_119);
and \U$12652 ( \12995 , RI98716e0_125, \2040 );
nor \U$12653 ( \12996 , \12994 , \12995 );
not \U$12654 ( \12997 , \12996 );
or \U$12655 ( \12998 , \12993 , \12997 );
or \U$12656 ( \12999 , \12996 , \2034 );
nand \U$12657 ( \13000 , \12998 , \12999 );
and \U$12658 ( \13001 , \12992 , \13000 );
and \U$12659 ( \13002 , \12984 , \12991 );
or \U$12660 ( \13003 , \13001 , \13002 );
and \U$12661 ( \13004 , \12977 , \13003 );
and \U$12662 ( \13005 , \12948 , \12976 );
or \U$12663 ( \13006 , \13004 , \13005 );
and \U$12664 ( \13007 , \8486 , RI986f8e0_61);
and \U$12665 ( \13008 , RI986f430_51, \8484 );
nor \U$12666 ( \13009 , \13007 , \13008 );
and \U$12667 ( \13010 , \13009 , \8050 );
not \U$12668 ( \13011 , \13009 );
and \U$12669 ( \13012 , \13011 , \8051 );
nor \U$12670 ( \13013 , \13010 , \13012 );
and \U$12671 ( \13014 , \7079 , RI986e620_21);
and \U$12672 ( \13015 , RI986f7f0_59, \7077 );
nor \U$12673 ( \13016 , \13014 , \13015 );
and \U$12674 ( \13017 , \13016 , \6710 );
not \U$12675 ( \13018 , \13016 );
and \U$12676 ( \13019 , \13018 , \6709 );
nor \U$12677 ( \13020 , \13017 , \13019 );
xor \U$12678 ( \13021 , \13013 , \13020 );
and \U$12679 ( \13022 , \7729 , RI986f700_57);
and \U$12680 ( \13023 , RI986f9d0_63, \7727 );
nor \U$12681 ( \13024 , \13022 , \13023 );
and \U$12682 ( \13025 , \13024 , \7480 );
not \U$12683 ( \13026 , \13024 );
and \U$12684 ( \13027 , \13026 , \7733 );
nor \U$12685 ( \13028 , \13025 , \13027 );
and \U$12686 ( \13029 , \13021 , \13028 );
and \U$12687 ( \13030 , \13013 , \13020 );
or \U$12688 ( \13031 , \13029 , \13030 );
and \U$12689 ( \13032 , \11696 , RI986dcc0_1);
and \U$12690 ( \13033 , RI986e170_11, \11694 );
nor \U$12691 ( \13034 , \13032 , \13033 );
and \U$12692 ( \13035 , \13034 , \10965 );
not \U$12693 ( \13036 , \13034 );
and \U$12694 ( \13037 , \13036 , \11702 );
nor \U$12695 ( \13038 , \13035 , \13037 );
and \U$12696 ( \13039 , RI9873288_184, RI9873378_186);
not \U$12697 ( \13040 , RI98733f0_187);
and \U$12698 ( \13041 , \13040 , RI9873378_186);
nor \U$12699 ( \13042 , \13040 , RI9873378_186);
or \U$12700 ( \13043 , \13041 , \13042 );
nor \U$12701 ( \13044 , RI9873288_184, RI9873378_186);
nor \U$12702 ( \13045 , \13039 , \13043 , \13044 );
nand \U$12703 ( \13046 , RI986e350_15, \13045 );
not \U$12704 ( \13047 , \12619 );
and \U$12705 ( \13048 , \13046 , \13047 );
not \U$12706 ( \13049 , \13046 );
and \U$12707 ( \13050 , \13049 , \12619 );
nor \U$12708 ( \13051 , \13048 , \13050 );
xor \U$12709 ( \13052 , \13038 , \13051 );
and \U$12710 ( \13053 , \12293 , RI986e080_9);
and \U$12711 ( \13054 , RI986e260_13, \12291 );
nor \U$12712 ( \13055 , \13053 , \13054 );
and \U$12713 ( \13056 , \13055 , \11687 );
not \U$12714 ( \13057 , \13055 );
and \U$12715 ( \13058 , \13057 , \11686 );
nor \U$12716 ( \13059 , \13056 , \13058 );
and \U$12717 ( \13060 , \13052 , \13059 );
and \U$12718 ( \13061 , \13038 , \13051 );
or \U$12719 ( \13062 , \13060 , \13061 );
xor \U$12720 ( \13063 , \13031 , \13062 );
and \U$12721 ( \13064 , \9505 , RI986f610_55);
and \U$12722 ( \13065 , RI986df90_7, \9503 );
nor \U$12723 ( \13066 , \13064 , \13065 );
and \U$12724 ( \13067 , \13066 , \9510 );
not \U$12725 ( \13068 , \13066 );
and \U$12726 ( \13069 , \13068 , \9513 );
nor \U$12727 ( \13070 , \13067 , \13069 );
and \U$12728 ( \13071 , \9237 , RI986f340_49);
and \U$12729 ( \13072 , RI986f520_53, \9235 );
nor \U$12730 ( \13073 , \13071 , \13072 );
and \U$12731 ( \13074 , \13073 , \9241 );
not \U$12732 ( \13075 , \13073 );
and \U$12733 ( \13076 , \13075 , \8836 );
nor \U$12734 ( \13077 , \13074 , \13076 );
xor \U$12735 ( \13078 , \13070 , \13077 );
and \U$12736 ( \13079 , \10424 , RI986dea0_5);
and \U$12737 ( \13080 , RI986ddb0_3, \10422 );
nor \U$12738 ( \13081 , \13079 , \13080 );
and \U$12739 ( \13082 , \13081 , \9840 );
not \U$12740 ( \13083 , \13081 );
and \U$12741 ( \13084 , \13083 , \10428 );
nor \U$12742 ( \13085 , \13082 , \13084 );
and \U$12743 ( \13086 , \13078 , \13085 );
and \U$12744 ( \13087 , \13070 , \13077 );
or \U$12745 ( \13088 , \13086 , \13087 );
and \U$12746 ( \13089 , \13063 , \13088 );
and \U$12747 ( \13090 , \13031 , \13062 );
or \U$12748 ( \13091 , \13089 , \13090 );
xor \U$12749 ( \13092 , \13006 , \13091 );
and \U$12750 ( \13093 , \5881 , RI986f160_45);
and \U$12751 ( \13094 , RI986e530_19, \5879 );
nor \U$12752 ( \13095 , \13093 , \13094 );
and \U$12753 ( \13096 , \13095 , \5594 );
not \U$12754 ( \13097 , \13095 );
and \U$12755 ( \13098 , \13097 , \5885 );
nor \U$12756 ( \13099 , \13096 , \13098 );
and \U$12757 ( \13100 , \5318 , RI986ef80_41);
and \U$12758 ( \13101 , RI986f250_47, \5316 );
nor \U$12759 ( \13102 , \13100 , \13101 );
and \U$12760 ( \13103 , \13102 , \5052 );
not \U$12761 ( \13104 , \13102 );
and \U$12762 ( \13105 , \13104 , \5322 );
nor \U$12763 ( \13106 , \13103 , \13105 );
xor \U$12764 ( \13107 , \13099 , \13106 );
and \U$12765 ( \13108 , \6453 , RI986e440_17);
and \U$12766 ( \13109 , RI986e710_23, \6451 );
nor \U$12767 ( \13110 , \13108 , \13109 );
and \U$12768 ( \13111 , \13110 , \6190 );
not \U$12769 ( \13112 , \13110 );
and \U$12770 ( \13113 , \13112 , \6180 );
nor \U$12771 ( \13114 , \13111 , \13113 );
and \U$12772 ( \13115 , \13107 , \13114 );
and \U$12773 ( \13116 , \13099 , \13106 );
or \U$12774 ( \13117 , \13115 , \13116 );
not \U$12775 ( \13118 , \3406 );
and \U$12776 ( \13119 , \3254 , RI986e9e0_29);
and \U$12777 ( \13120 , RI986e8f0_27, \3252 );
nor \U$12778 ( \13121 , \13119 , \13120 );
not \U$12779 ( \13122 , \13121 );
or \U$12780 ( \13123 , \13118 , \13122 );
or \U$12781 ( \13124 , \13121 , \3406 );
nand \U$12782 ( \13125 , \13123 , \13124 );
and \U$12783 ( \13126 , \2274 , RI98717d0_127);
and \U$12784 ( \13127 , RI9871500_121, \2272 );
nor \U$12785 ( \13128 , \13126 , \13127 );
and \U$12786 ( \13129 , \13128 , \2030 );
not \U$12787 ( \13130 , \13128 );
and \U$12788 ( \13131 , \13130 , \2031 );
nor \U$12789 ( \13132 , \13129 , \13131 );
xor \U$12790 ( \13133 , \13125 , \13132 );
and \U$12791 ( \13134 , \2464 , RI98715f0_123);
and \U$12792 ( \13135 , RI986ead0_31, \2462 );
nor \U$12793 ( \13136 , \13134 , \13135 );
and \U$12794 ( \13137 , \13136 , \2468 );
not \U$12795 ( \13138 , \13136 );
and \U$12796 ( \13139 , \13138 , \2263 );
nor \U$12797 ( \13140 , \13137 , \13139 );
and \U$12798 ( \13141 , \13133 , \13140 );
and \U$12799 ( \13142 , \13125 , \13132 );
or \U$12800 ( \13143 , \13141 , \13142 );
xor \U$12801 ( \13144 , \13117 , \13143 );
and \U$12802 ( \13145 , \4203 , RI986eda0_37);
and \U$12803 ( \13146 , RI986ebc0_33, \4201 );
nor \U$12804 ( \13147 , \13145 , \13146 );
and \U$12805 ( \13148 , \13147 , \4207 );
not \U$12806 ( \13149 , \13147 );
and \U$12807 ( \13150 , \13149 , \3923 );
nor \U$12808 ( \13151 , \13148 , \13150 );
not \U$12809 ( \13152 , \3412 );
and \U$12810 ( \13153 , \3683 , RI986e800_25);
and \U$12811 ( \13154 , RI986ee90_39, \3681 );
nor \U$12812 ( \13155 , \13153 , \13154 );
not \U$12813 ( \13156 , \13155 );
or \U$12814 ( \13157 , \13152 , \13156 );
or \U$12815 ( \13158 , \13155 , \3412 );
nand \U$12816 ( \13159 , \13157 , \13158 );
xor \U$12817 ( \13160 , \13151 , \13159 );
not \U$12818 ( \13161 , \4521 );
and \U$12819 ( \13162 , \4710 , RI986ecb0_35);
and \U$12820 ( \13163 , RI986f070_43, \4708 );
nor \U$12821 ( \13164 , \13162 , \13163 );
not \U$12822 ( \13165 , \13164 );
or \U$12823 ( \13166 , \13161 , \13165 );
or \U$12824 ( \13167 , \13164 , \4521 );
nand \U$12825 ( \13168 , \13166 , \13167 );
and \U$12826 ( \13169 , \13160 , \13168 );
and \U$12827 ( \13170 , \13151 , \13159 );
or \U$12828 ( \13171 , \13169 , \13170 );
and \U$12829 ( \13172 , \13144 , \13171 );
and \U$12830 ( \13173 , \13117 , \13143 );
or \U$12831 ( \13174 , \13172 , \13173 );
and \U$12832 ( \13175 , \13092 , \13174 );
and \U$12833 ( \13176 , \13006 , \13091 );
or \U$12834 ( \13177 , \13175 , \13176 );
xor \U$12835 ( \13178 , \12922 , \13177 );
xor \U$12836 ( \13179 , \12536 , \12543 );
xor \U$12837 ( \13180 , \13179 , \12552 );
xor \U$12838 ( \13181 , \12697 , \12704 );
xor \U$12839 ( \13182 , \13181 , \12712 );
and \U$12840 ( \13183 , \13180 , \13182 );
xor \U$12841 ( \13184 , \12563 , \12570 );
xor \U$12842 ( \13185 , \13184 , \12579 );
xor \U$12843 ( \13186 , \12697 , \12704 );
xor \U$12844 ( \13187 , \13186 , \12712 );
and \U$12845 ( \13188 , \13185 , \13187 );
and \U$12846 ( \13189 , \13180 , \13185 );
or \U$12847 ( \13190 , \13183 , \13188 , \13189 );
and \U$12848 ( \13191 , \416 , RI98707e0_93);
and \U$12849 ( \13192 , RI986fac0_65, \414 );
nor \U$12850 ( \13193 , \13191 , \13192 );
and \U$12851 ( \13194 , \13193 , \421 );
not \U$12852 ( \13195 , \13193 );
and \U$12853 ( \13196 , \13195 , \422 );
nor \U$12854 ( \13197 , \13194 , \13196 );
nand \U$12855 ( \13198 , RI98708d0_95, RI9871fc8_144);
or \U$12856 ( \13199 , \13197 , \13198 );
not \U$12857 ( \13200 , \13198 );
not \U$12858 ( \13201 , \13197 );
or \U$12859 ( \13202 , \13200 , \13201 );
not \U$12860 ( \13203 , \345 );
and \U$12861 ( \13204 , \354 , RI986fbb0_67);
and \U$12862 ( \13205 , RI986fd90_71, \352 );
nor \U$12863 ( \13206 , \13204 , \13205 );
not \U$12864 ( \13207 , \13206 );
or \U$12865 ( \13208 , \13203 , \13207 );
or \U$12866 ( \13209 , \13206 , \361 );
nand \U$12867 ( \13210 , \13208 , \13209 );
nand \U$12868 ( \13211 , \13202 , \13210 );
nand \U$12869 ( \13212 , \13199 , \13211 );
xor \U$12870 ( \13213 , \12509 , \12517 );
xor \U$12871 ( \13214 , \13213 , \12526 );
and \U$12872 ( \13215 , \13212 , \13214 );
xor \U$12873 ( \13216 , \12466 , \12468 );
xor \U$12874 ( \13217 , \13216 , \12476 );
xor \U$12875 ( \13218 , \12509 , \12517 );
xor \U$12876 ( \13219 , \13218 , \12526 );
and \U$12877 ( \13220 , \13217 , \13219 );
and \U$12878 ( \13221 , \13212 , \13217 );
or \U$12879 ( \13222 , \13215 , \13220 , \13221 );
xor \U$12880 ( \13223 , \13190 , \13222 );
xor \U$12881 ( \13224 , \12670 , \12678 );
xor \U$12882 ( \13225 , \13224 , \12686 );
xor \U$12883 ( \13226 , \12723 , \12730 );
xor \U$12884 ( \13227 , \13226 , \12738 );
xor \U$12885 ( \13228 , \13225 , \13227 );
xor \U$12886 ( \13229 , \12640 , \12647 );
xor \U$12887 ( \13230 , \13229 , \12655 );
and \U$12888 ( \13231 , \13228 , \13230 );
and \U$12889 ( \13232 , \13225 , \13227 );
or \U$12890 ( \13233 , \13231 , \13232 );
and \U$12891 ( \13234 , \13223 , \13233 );
and \U$12892 ( \13235 , \13190 , \13222 );
or \U$12893 ( \13236 , \13234 , \13235 );
and \U$12894 ( \13237 , \13178 , \13236 );
and \U$12895 ( \13238 , \12922 , \13177 );
or \U$12896 ( \13239 , \13237 , \13238 );
xor \U$12897 ( \13240 , \12910 , \13239 );
xor \U$12898 ( \13241 , \12529 , \12555 );
xor \U$12899 ( \13242 , \13241 , \12582 );
xor \U$12900 ( \13243 , \12490 , \12492 );
xor \U$12901 ( \13244 , \13243 , \12495 );
and \U$12902 ( \13245 , \13242 , \13244 );
xor \U$12903 ( \13246 , \12479 , \12481 );
xor \U$12904 ( \13247 , \13246 , \12484 );
xor \U$12905 ( \13248 , \12490 , \12492 );
xor \U$12906 ( \13249 , \13248 , \12495 );
and \U$12907 ( \13250 , \13247 , \13249 );
and \U$12908 ( \13251 , \13242 , \13247 );
or \U$12909 ( \13252 , \13245 , \13250 , \13251 );
xor \U$12910 ( \13253 , \12279 , \12309 );
xor \U$12911 ( \13254 , \13253 , \12335 );
xor \U$12912 ( \13255 , \13252 , \13254 );
xor \U$12913 ( \13256 , \12365 , \12393 );
xor \U$12914 ( \13257 , \13256 , \12420 );
xor \U$12915 ( \13258 , \12770 , \12775 );
xor \U$12916 ( \13259 , \13257 , \13258 );
and \U$12917 ( \13260 , \13255 , \13259 );
and \U$12918 ( \13261 , \13252 , \13254 );
or \U$12919 ( \13262 , \13260 , \13261 );
and \U$12920 ( \13263 , \13240 , \13262 );
and \U$12921 ( \13264 , \12910 , \13239 );
or \U$12922 ( \13265 , \13263 , \13264 );
xor \U$12923 ( \13266 , \12828 , \12836 );
xor \U$12924 ( \13267 , \13266 , \12841 );
xor \U$12925 ( \13268 , \13265 , \13267 );
xor \U$12926 ( \13269 , \12501 , \12747 );
xor \U$12927 ( \13270 , \13269 , \12764 );
xor \U$12928 ( \13271 , \12171 , \12424 );
xor \U$12929 ( \13272 , \13271 , \12443 );
and \U$12930 ( \13273 , \13270 , \13272 );
xor \U$12931 ( \13274 , \12081 , \12083 );
xor \U$12932 ( \13275 , \13274 , \12086 );
xor \U$12933 ( \13276 , \12780 , \12787 );
xor \U$12934 ( \13277 , \13275 , \13276 );
xor \U$12935 ( \13278 , \12171 , \12424 );
xor \U$12936 ( \13279 , \13278 , \12443 );
and \U$12937 ( \13280 , \13277 , \13279 );
and \U$12938 ( \13281 , \13270 , \13277 );
or \U$12939 ( \13282 , \13273 , \13280 , \13281 );
and \U$12940 ( \13283 , \13268 , \13282 );
and \U$12941 ( \13284 , \13265 , \13267 );
or \U$12942 ( \13285 , \13283 , \13284 );
and \U$12943 ( \13286 , \12896 , \13285 );
and \U$12944 ( \13287 , \12893 , \12895 );
or \U$12945 ( \13288 , \13286 , \13287 );
xor \U$12946 ( \13289 , \12809 , \12811 );
xor \U$12947 ( \13290 , \13289 , \12862 );
xor \U$12948 ( \13291 , \13288 , \13290 );
not \U$12949 ( \13292 , \13291 );
xor \U$12950 ( \13293 , \12922 , \13177 );
xor \U$12951 ( \13294 , \13293 , \13236 );
xor \U$12952 ( \13295 , \13252 , \13254 );
xor \U$12953 ( \13296 , \13295 , \13259 );
and \U$12954 ( \13297 , \13294 , \13296 );
xor \U$12955 ( \13298 , \12458 , \12487 );
xor \U$12956 ( \13299 , \13298 , \12498 );
xor \U$12957 ( \13300 , \12898 , \12905 );
xor \U$12958 ( \13301 , \13299 , \13300 );
xor \U$12959 ( \13302 , \13252 , \13254 );
xor \U$12960 ( \13303 , \13302 , \13259 );
and \U$12961 ( \13304 , \13301 , \13303 );
and \U$12962 ( \13305 , \13294 , \13301 );
or \U$12963 ( \13306 , \13297 , \13304 , \13305 );
xor \U$12964 ( \13307 , \12610 , \12632 );
xor \U$12965 ( \13308 , \13307 , \12658 );
xor \U$12966 ( \13309 , \12912 , \12914 );
xor \U$12967 ( \13310 , \13309 , \12919 );
and \U$12968 ( \13311 , \13308 , \13310 );
xor \U$12969 ( \13312 , \12490 , \12492 );
xor \U$12970 ( \13313 , \13312 , \12495 );
xor \U$12971 ( \13314 , \13242 , \13247 );
xor \U$12972 ( \13315 , \13313 , \13314 );
xor \U$12973 ( \13316 , \12912 , \12914 );
xor \U$12974 ( \13317 , \13316 , \12919 );
and \U$12975 ( \13318 , \13315 , \13317 );
and \U$12976 ( \13319 , \13308 , \13315 );
or \U$12977 ( \13320 , \13311 , \13318 , \13319 );
and \U$12978 ( \13321 , \7729 , RI986f7f0_59);
and \U$12979 ( \13322 , RI986f700_57, \7727 );
nor \U$12980 ( \13323 , \13321 , \13322 );
and \U$12981 ( \13324 , \13323 , \7733 );
not \U$12982 ( \13325 , \13323 );
and \U$12983 ( \13326 , \13325 , \7480 );
nor \U$12984 ( \13327 , \13324 , \13326 );
and \U$12985 ( \13328 , \8486 , RI986f9d0_63);
and \U$12986 ( \13329 , RI986f8e0_61, \8484 );
nor \U$12987 ( \13330 , \13328 , \13329 );
and \U$12988 ( \13331 , \13330 , \8051 );
not \U$12989 ( \13332 , \13330 );
and \U$12990 ( \13333 , \13332 , \8050 );
nor \U$12991 ( \13334 , \13331 , \13333 );
or \U$12992 ( \13335 , \13327 , \13334 );
not \U$12993 ( \13336 , \13334 );
not \U$12994 ( \13337 , \13327 );
or \U$12995 ( \13338 , \13336 , \13337 );
and \U$12996 ( \13339 , \9237 , RI986f430_51);
and \U$12997 ( \13340 , RI986f340_49, \9235 );
nor \U$12998 ( \13341 , \13339 , \13340 );
and \U$12999 ( \13342 , \13341 , \9241 );
not \U$13000 ( \13343 , \13341 );
and \U$13001 ( \13344 , \13343 , \8836 );
nor \U$13002 ( \13345 , \13342 , \13344 );
nand \U$13003 ( \13346 , \13338 , \13345 );
nand \U$13004 ( \13347 , \13335 , \13346 );
and \U$13005 ( \13348 , \12293 , RI986e170_11);
and \U$13006 ( \13349 , RI986e080_9, \12291 );
nor \U$13007 ( \13350 , \13348 , \13349 );
and \U$13008 ( \13351 , \13350 , \11686 );
not \U$13009 ( \13352 , \13350 );
and \U$13010 ( \13353 , \13352 , \11687 );
nor \U$13011 ( \13354 , \13351 , \13353 );
not \U$13012 ( \13355 , RI98734e0_189);
not \U$13013 ( \13356 , RI9873468_188);
or \U$13014 ( \13357 , \13355 , \13356 );
nand \U$13015 ( \13358 , \13357 , RI98733f0_187);
not \U$13016 ( \13359 , \13358 );
or \U$13017 ( \13360 , \13354 , \13359 );
not \U$13018 ( \13361 , \13359 );
not \U$13019 ( \13362 , \13354 );
or \U$13020 ( \13363 , \13361 , \13362 );
and \U$13021 ( \13364 , \13045 , RI986e260_13);
and \U$13022 ( \13365 , RI986e350_15, \13043 );
nor \U$13023 ( \13366 , \13364 , \13365 );
and \U$13024 ( \13367 , \13366 , \13047 );
not \U$13025 ( \13368 , \13366 );
and \U$13026 ( \13369 , \13368 , \12619 );
nor \U$13027 ( \13370 , \13367 , \13369 );
nand \U$13028 ( \13371 , \13363 , \13370 );
nand \U$13029 ( \13372 , \13360 , \13371 );
xor \U$13030 ( \13373 , \13347 , \13372 );
and \U$13031 ( \13374 , \9505 , RI986f520_53);
and \U$13032 ( \13375 , RI986f610_55, \9503 );
nor \U$13033 ( \13376 , \13374 , \13375 );
and \U$13034 ( \13377 , \13376 , \9513 );
not \U$13035 ( \13378 , \13376 );
and \U$13036 ( \13379 , \13378 , \9510 );
nor \U$13037 ( \13380 , \13377 , \13379 );
and \U$13038 ( \13381 , \10424 , RI986df90_7);
and \U$13039 ( \13382 , RI986dea0_5, \10422 );
nor \U$13040 ( \13383 , \13381 , \13382 );
and \U$13041 ( \13384 , \13383 , \10428 );
not \U$13042 ( \13385 , \13383 );
and \U$13043 ( \13386 , \13385 , \9840 );
nor \U$13044 ( \13387 , \13384 , \13386 );
or \U$13045 ( \13388 , \13380 , \13387 );
not \U$13046 ( \13389 , \13387 );
not \U$13047 ( \13390 , \13380 );
or \U$13048 ( \13391 , \13389 , \13390 );
and \U$13049 ( \13392 , \11696 , RI986ddb0_3);
and \U$13050 ( \13393 , RI986dcc0_1, \11694 );
nor \U$13051 ( \13394 , \13392 , \13393 );
and \U$13052 ( \13395 , \13394 , \10965 );
not \U$13053 ( \13396 , \13394 );
and \U$13054 ( \13397 , \13396 , \11702 );
nor \U$13055 ( \13398 , \13395 , \13397 );
nand \U$13056 ( \13399 , \13391 , \13398 );
nand \U$13057 ( \13400 , \13388 , \13399 );
and \U$13058 ( \13401 , \13373 , \13400 );
and \U$13059 ( \13402 , \13347 , \13372 );
nor \U$13060 ( \13403 , \13401 , \13402 );
and \U$13061 ( \13404 , \6453 , RI986e530_19);
and \U$13062 ( \13405 , RI986e440_17, \6451 );
nor \U$13063 ( \13406 , \13404 , \13405 );
and \U$13064 ( \13407 , \13406 , \6180 );
not \U$13065 ( \13408 , \13406 );
and \U$13066 ( \13409 , \13408 , \6190 );
nor \U$13067 ( \13410 , \13407 , \13409 );
and \U$13068 ( \13411 , \7079 , RI986e710_23);
and \U$13069 ( \13412 , RI986e620_21, \7077 );
nor \U$13070 ( \13413 , \13411 , \13412 );
and \U$13071 ( \13414 , \13413 , \6709 );
not \U$13072 ( \13415 , \13413 );
and \U$13073 ( \13416 , \13415 , \6710 );
nor \U$13074 ( \13417 , \13414 , \13416 );
xor \U$13075 ( \13418 , \13410 , \13417 );
and \U$13076 ( \13419 , \5881 , RI986f250_47);
and \U$13077 ( \13420 , RI986f160_45, \5879 );
nor \U$13078 ( \13421 , \13419 , \13420 );
and \U$13079 ( \13422 , \13421 , \5885 );
not \U$13080 ( \13423 , \13421 );
and \U$13081 ( \13424 , \13423 , \5594 );
nor \U$13082 ( \13425 , \13422 , \13424 );
and \U$13083 ( \13426 , \13418 , \13425 );
and \U$13084 ( \13427 , \13410 , \13417 );
nor \U$13085 ( \13428 , \13426 , \13427 );
and \U$13086 ( \13429 , \4203 , RI986ee90_39);
and \U$13087 ( \13430 , RI986eda0_37, \4201 );
nor \U$13088 ( \13431 , \13429 , \13430 );
and \U$13089 ( \13432 , \13431 , \3922 );
not \U$13090 ( \13433 , \13431 );
and \U$13091 ( \13434 , \13433 , \4207 );
nor \U$13092 ( \13435 , \13432 , \13434 );
and \U$13093 ( \13436 , \4710 , RI986ebc0_33);
and \U$13094 ( \13437 , RI986ecb0_35, \4708 );
nor \U$13095 ( \13438 , \13436 , \13437 );
not \U$13096 ( \13439 , \13438 );
not \U$13097 ( \13440 , \4521 );
and \U$13098 ( \13441 , \13439 , \13440 );
and \U$13099 ( \13442 , \13438 , \4519 );
nor \U$13100 ( \13443 , \13441 , \13442 );
or \U$13101 ( \13444 , \13435 , \13443 );
not \U$13102 ( \13445 , \13443 );
not \U$13103 ( \13446 , \13435 );
or \U$13104 ( \13447 , \13445 , \13446 );
and \U$13105 ( \13448 , \5318 , RI986f070_43);
and \U$13106 ( \13449 , RI986ef80_41, \5316 );
nor \U$13107 ( \13450 , \13448 , \13449 );
and \U$13108 ( \13451 , \13450 , \5052 );
not \U$13109 ( \13452 , \13450 );
and \U$13110 ( \13453 , \13452 , \5322 );
nor \U$13111 ( \13454 , \13451 , \13453 );
nand \U$13112 ( \13455 , \13447 , \13454 );
nand \U$13113 ( \13456 , \13444 , \13455 );
xor \U$13114 ( \13457 , \13428 , \13456 );
and \U$13115 ( \13458 , \2464 , RI9871500_121);
and \U$13116 ( \13459 , RI98715f0_123, \2462 );
nor \U$13117 ( \13460 , \13458 , \13459 );
and \U$13118 ( \13461 , \13460 , \2263 );
not \U$13119 ( \13462 , \13460 );
and \U$13120 ( \13463 , \13462 , \2468 );
nor \U$13121 ( \13464 , \13461 , \13463 );
and \U$13122 ( \13465 , \3254 , RI986ead0_31);
and \U$13123 ( \13466 , RI986e9e0_29, \3252 );
nor \U$13124 ( \13467 , \13465 , \13466 );
not \U$13125 ( \13468 , \13467 );
not \U$13126 ( \13469 , \2935 );
and \U$13127 ( \13470 , \13468 , \13469 );
and \U$13128 ( \13471 , \13467 , \3406 );
nor \U$13129 ( \13472 , \13470 , \13471 );
or \U$13130 ( \13473 , \13464 , \13472 );
not \U$13131 ( \13474 , \13472 );
not \U$13132 ( \13475 , \13464 );
or \U$13133 ( \13476 , \13474 , \13475 );
not \U$13134 ( \13477 , \3918 );
and \U$13135 ( \13478 , \3683 , RI986e8f0_27);
and \U$13136 ( \13479 , RI986e800_25, \3681 );
nor \U$13137 ( \13480 , \13478 , \13479 );
not \U$13138 ( \13481 , \13480 );
or \U$13139 ( \13482 , \13477 , \13481 );
or \U$13140 ( \13483 , \13480 , \3918 );
nand \U$13141 ( \13484 , \13482 , \13483 );
nand \U$13142 ( \13485 , \13476 , \13484 );
nand \U$13143 ( \13486 , \13473 , \13485 );
and \U$13144 ( \13487 , \13457 , \13486 );
and \U$13145 ( \13488 , \13428 , \13456 );
nor \U$13146 ( \13489 , \13487 , \13488 );
xor \U$13147 ( \13490 , \13403 , \13489 );
and \U$13148 ( \13491 , \776 , RI9870d80_105);
and \U$13149 ( \13492 , RI98709c0_97, \774 );
nor \U$13150 ( \13493 , \13491 , \13492 );
and \U$13151 ( \13494 , \13493 , \451 );
not \U$13152 ( \13495 , \13493 );
and \U$13153 ( \13496 , \13495 , \474 );
nor \U$13154 ( \13497 , \13494 , \13496 );
and \U$13155 ( \13498 , \1293 , RI9870e70_107);
and \U$13156 ( \13499 , RI9870ba0_101, \1291 );
nor \U$13157 ( \13500 , \13498 , \13499 );
not \U$13158 ( \13501 , \13500 );
not \U$13159 ( \13502 , \1128 );
and \U$13160 ( \13503 , \13501 , \13502 );
and \U$13161 ( \13504 , \13500 , \1128 );
nor \U$13162 ( \13505 , \13503 , \13504 );
or \U$13163 ( \13506 , \13497 , \13505 );
not \U$13164 ( \13507 , \13505 );
not \U$13165 ( \13508 , \13497 );
or \U$13166 ( \13509 , \13507 , \13508 );
and \U$13167 ( \13510 , \1329 , RI9871050_111);
and \U$13168 ( \13511 , RI9870c90_103, \1327 );
nor \U$13169 ( \13512 , \13510 , \13511 );
and \U$13170 ( \13513 , \13512 , \1336 );
not \U$13171 ( \13514 , \13512 );
and \U$13172 ( \13515 , \13514 , \1337 );
nor \U$13173 ( \13516 , \13513 , \13515 );
nand \U$13174 ( \13517 , \13509 , \13516 );
nand \U$13175 ( \13518 , \13506 , \13517 );
and \U$13176 ( \13519 , \465 , RI9870060_77);
and \U$13177 ( \13520 , RI9870150_79, \463 );
nor \U$13178 ( \13521 , \13519 , \13520 );
not \U$13179 ( \13522 , \13521 );
not \U$13180 ( \13523 , \454 );
and \U$13181 ( \13524 , \13522 , \13523 );
and \U$13182 ( \13525 , \13521 , \456 );
nor \U$13183 ( \13526 , \13524 , \13525 );
and \U$13184 ( \13527 , \376 , RI986ff70_75);
and \U$13185 ( \13528 , RI986fe80_73, \374 );
nor \U$13186 ( \13529 , \13527 , \13528 );
not \U$13187 ( \13530 , \13529 );
not \U$13188 ( \13531 , \367 );
and \U$13189 ( \13532 , \13530 , \13531 );
and \U$13190 ( \13533 , \13529 , \367 );
nor \U$13191 ( \13534 , \13532 , \13533 );
or \U$13192 ( \13535 , \13526 , \13534 );
not \U$13193 ( \13536 , \13534 );
not \U$13194 ( \13537 , \13526 );
or \U$13195 ( \13538 , \13536 , \13537 );
and \U$13196 ( \13539 , \438 , RI9870f60_109);
and \U$13197 ( \13540 , RI9870ab0_99, \436 );
nor \U$13198 ( \13541 , \13539 , \13540 );
and \U$13199 ( \13542 , \13541 , \444 );
not \U$13200 ( \13543 , \13541 );
and \U$13201 ( \13544 , \13543 , \443 );
nor \U$13202 ( \13545 , \13542 , \13544 );
nand \U$13203 ( \13546 , \13538 , \13545 );
nand \U$13204 ( \13547 , \13535 , \13546 );
xor \U$13205 ( \13548 , \13518 , \13547 );
and \U$13206 ( \13549 , \2274 , RI98716e0_125);
and \U$13207 ( \13550 , RI98717d0_127, \2272 );
nor \U$13208 ( \13551 , \13549 , \13550 );
and \U$13209 ( \13552 , \13551 , \2030 );
not \U$13210 ( \13553 , \13551 );
and \U$13211 ( \13554 , \13553 , \2031 );
nor \U$13212 ( \13555 , \13552 , \13554 );
and \U$13213 ( \13556 , \1311 , RI9871230_115);
and \U$13214 ( \13557 , RI9871140_113, \1309 );
nor \U$13215 ( \13558 , \13556 , \13557 );
and \U$13216 ( \13559 , \13558 , \1458 );
not \U$13217 ( \13560 , \13558 );
and \U$13218 ( \13561 , \13560 , \1318 );
nor \U$13219 ( \13562 , \13559 , \13561 );
xor \U$13220 ( \13563 , \13555 , \13562 );
not \U$13221 ( \13564 , \1462 );
and \U$13222 ( \13565 , \2042 , RI9871320_117);
and \U$13223 ( \13566 , RI9871410_119, \2040 );
nor \U$13224 ( \13567 , \13565 , \13566 );
not \U$13225 ( \13568 , \13567 );
or \U$13226 ( \13569 , \13564 , \13568 );
or \U$13227 ( \13570 , \13567 , \2034 );
nand \U$13228 ( \13571 , \13569 , \13570 );
and \U$13229 ( \13572 , \13563 , \13571 );
and \U$13230 ( \13573 , \13555 , \13562 );
or \U$13231 ( \13574 , \13572 , \13573 );
and \U$13232 ( \13575 , \13548 , \13574 );
and \U$13233 ( \13576 , \13518 , \13547 );
nor \U$13234 ( \13577 , \13575 , \13576 );
and \U$13235 ( \13578 , \13490 , \13577 );
and \U$13236 ( \13579 , \13403 , \13489 );
nor \U$13237 ( \13580 , \13578 , \13579 );
and \U$13238 ( \13581 , \12630 , \13047 );
not \U$13239 ( \13582 , \12630 );
and \U$13240 ( \13583 , \13582 , \12619 );
nor \U$13241 ( \13584 , \13581 , \13583 );
not \U$13242 ( \13585 , \13584 );
not \U$13243 ( \13586 , \12617 );
and \U$13244 ( \13587 , \13585 , \13586 );
and \U$13245 ( \13588 , \13584 , \12617 );
nor \U$13246 ( \13589 , \13587 , \13588 );
xor \U$13247 ( \13590 , \12592 , \12599 );
xor \U$13248 ( \13591 , \13590 , \12607 );
or \U$13249 ( \13592 , \13589 , \13591 );
not \U$13250 ( \13593 , \13591 );
not \U$13251 ( \13594 , \13589 );
or \U$13252 ( \13595 , \13593 , \13594 );
xor \U$13253 ( \13596 , \13038 , \13051 );
xor \U$13254 ( \13597 , \13596 , \13059 );
xor \U$13255 ( \13598 , \13013 , \13020 );
xor \U$13256 ( \13599 , \13598 , \13028 );
and \U$13257 ( \13600 , \13597 , \13599 );
xor \U$13258 ( \13601 , \13070 , \13077 );
xor \U$13259 ( \13602 , \13601 , \13085 );
xor \U$13260 ( \13603 , \13013 , \13020 );
xor \U$13261 ( \13604 , \13603 , \13028 );
and \U$13262 ( \13605 , \13602 , \13604 );
and \U$13263 ( \13606 , \13597 , \13602 );
or \U$13264 ( \13607 , \13600 , \13605 , \13606 );
nand \U$13265 ( \13608 , \13595 , \13607 );
nand \U$13266 ( \13609 , \13592 , \13608 );
xor \U$13267 ( \13610 , \13580 , \13609 );
xor \U$13268 ( \13611 , \12956 , \12964 );
xor \U$13269 ( \13612 , \13611 , \12973 );
xor \U$13270 ( \13613 , \12984 , \12991 );
xor \U$13271 ( \13614 , \13613 , \13000 );
and \U$13272 ( \13615 , \13612 , \13614 );
xor \U$13273 ( \13616 , \12930 , \12937 );
xor \U$13274 ( \13617 , \13616 , \12945 );
xor \U$13275 ( \13618 , \12984 , \12991 );
xor \U$13276 ( \13619 , \13618 , \13000 );
and \U$13277 ( \13620 , \13617 , \13619 );
and \U$13278 ( \13621 , \13612 , \13617 );
or \U$13279 ( \13622 , \13615 , \13620 , \13621 );
not \U$13280 ( \13623 , \386 );
and \U$13281 ( \13624 , \395 , RI986fd90_71);
and \U$13282 ( \13625 , RI986fca0_69, \393 );
nor \U$13283 ( \13626 , \13624 , \13625 );
not \U$13284 ( \13627 , \13626 );
or \U$13285 ( \13628 , \13623 , \13627 );
or \U$13286 ( \13629 , \13626 , \487 );
nand \U$13287 ( \13630 , \13628 , \13629 );
not \U$13288 ( \13631 , \345 );
and \U$13289 ( \13632 , \354 , RI986fac0_65);
and \U$13290 ( \13633 , RI986fbb0_67, \352 );
nor \U$13291 ( \13634 , \13632 , \13633 );
not \U$13292 ( \13635 , \13634 );
or \U$13293 ( \13636 , \13631 , \13635 );
or \U$13294 ( \13637 , \13634 , \361 );
nand \U$13295 ( \13638 , \13636 , \13637 );
xor \U$13296 ( \13639 , \13630 , \13638 );
and \U$13297 ( \13640 , \416 , RI98708d0_95);
and \U$13298 ( \13641 , RI98707e0_93, \414 );
nor \U$13299 ( \13642 , \13640 , \13641 );
and \U$13300 ( \13643 , \13642 , \422 );
not \U$13301 ( \13644 , \13642 );
and \U$13302 ( \13645 , \13644 , \421 );
nor \U$13303 ( \13646 , \13643 , \13645 );
and \U$13304 ( \13647 , \13639 , \13646 );
and \U$13305 ( \13648 , \13630 , \13638 );
nor \U$13306 ( \13649 , \13647 , \13648 );
not \U$13307 ( \13650 , \13197 );
not \U$13308 ( \13651 , \13210 );
or \U$13309 ( \13652 , \13650 , \13651 );
or \U$13310 ( \13653 , \13197 , \13210 );
nand \U$13311 ( \13654 , \13652 , \13653 );
not \U$13312 ( \13655 , \13654 );
not \U$13313 ( \13656 , \13198 );
and \U$13314 ( \13657 , \13655 , \13656 );
and \U$13315 ( \13658 , \13654 , \13198 );
nor \U$13316 ( \13659 , \13657 , \13658 );
nand \U$13317 ( \13660 , \13649 , \13659 );
xor \U$13318 ( \13661 , \13622 , \13660 );
xor \U$13319 ( \13662 , \13125 , \13132 );
xor \U$13320 ( \13663 , \13662 , \13140 );
xor \U$13321 ( \13664 , \13099 , \13106 );
xor \U$13322 ( \13665 , \13664 , \13114 );
and \U$13323 ( \13666 , \13663 , \13665 );
xor \U$13324 ( \13667 , \13151 , \13159 );
xor \U$13325 ( \13668 , \13667 , \13168 );
xor \U$13326 ( \13669 , \13099 , \13106 );
xor \U$13327 ( \13670 , \13669 , \13114 );
and \U$13328 ( \13671 , \13668 , \13670 );
and \U$13329 ( \13672 , \13663 , \13668 );
or \U$13330 ( \13673 , \13666 , \13671 , \13672 );
and \U$13331 ( \13674 , \13661 , \13673 );
and \U$13332 ( \13675 , \13622 , \13660 );
or \U$13333 ( \13676 , \13674 , \13675 );
and \U$13334 ( \13677 , \13610 , \13676 );
and \U$13335 ( \13678 , \13580 , \13609 );
or \U$13336 ( \13679 , \13677 , \13678 );
xor \U$13337 ( \13680 , \13320 , \13679 );
xor \U$13338 ( \13681 , \13031 , \13062 );
xor \U$13339 ( \13682 , \13681 , \13088 );
xor \U$13340 ( \13683 , \12948 , \12976 );
xor \U$13341 ( \13684 , \13683 , \13003 );
xor \U$13342 ( \13685 , \13682 , \13684 );
xor \U$13343 ( \13686 , \13117 , \13143 );
xor \U$13344 ( \13687 , \13686 , \13171 );
and \U$13345 ( \13688 , \13685 , \13687 );
and \U$13346 ( \13689 , \13682 , \13684 );
or \U$13347 ( \13690 , \13688 , \13689 );
xor \U$13348 ( \13691 , \12689 , \12715 );
xor \U$13349 ( \13692 , \13691 , \12741 );
xor \U$13350 ( \13693 , \13690 , \13692 );
xor \U$13351 ( \13694 , \12509 , \12517 );
xor \U$13352 ( \13695 , \13694 , \12526 );
xor \U$13353 ( \13696 , \13212 , \13217 );
xor \U$13354 ( \13697 , \13695 , \13696 );
xor \U$13355 ( \13698 , \13225 , \13227 );
xor \U$13356 ( \13699 , \13698 , \13230 );
and \U$13357 ( \13700 , \13697 , \13699 );
xor \U$13358 ( \13701 , \12697 , \12704 );
xor \U$13359 ( \13702 , \13701 , \12712 );
xor \U$13360 ( \13703 , \13180 , \13185 );
xor \U$13361 ( \13704 , \13702 , \13703 );
xor \U$13362 ( \13705 , \13225 , \13227 );
xor \U$13363 ( \13706 , \13705 , \13230 );
and \U$13364 ( \13707 , \13704 , \13706 );
and \U$13365 ( \13708 , \13697 , \13704 );
or \U$13366 ( \13709 , \13700 , \13707 , \13708 );
and \U$13367 ( \13710 , \13693 , \13709 );
and \U$13368 ( \13711 , \13690 , \13692 );
or \U$13369 ( \13712 , \13710 , \13711 );
and \U$13370 ( \13713 , \13680 , \13712 );
and \U$13371 ( \13714 , \13320 , \13679 );
or \U$13372 ( \13715 , \13713 , \13714 );
xor \U$13373 ( \13716 , \13306 , \13715 );
xor \U$13374 ( \13717 , \12171 , \12424 );
xor \U$13375 ( \13718 , \13717 , \12443 );
xor \U$13376 ( \13719 , \13270 , \13277 );
xor \U$13377 ( \13720 , \13718 , \13719 );
and \U$13378 ( \13721 , \13716 , \13720 );
and \U$13379 ( \13722 , \13306 , \13715 );
or \U$13380 ( \13723 , \13721 , \13722 );
xor \U$13381 ( \13724 , \12888 , \12892 );
xor \U$13382 ( \13725 , \13723 , \13724 );
xor \U$13383 ( \13726 , \13265 , \13267 );
xor \U$13384 ( \13727 , \13726 , \13282 );
and \U$13385 ( \13728 , \13725 , \13727 );
and \U$13386 ( \13729 , \13723 , \13724 );
or \U$13387 ( \13730 , \13728 , \13729 );
xor \U$13388 ( \13731 , \12125 , \12795 );
xor \U$13389 ( \13732 , \13731 , \12806 );
xor \U$13390 ( \13733 , \13730 , \13732 );
xor \U$13391 ( \13734 , \12893 , \12895 );
xor \U$13392 ( \13735 , \13734 , \13285 );
and \U$13393 ( \13736 , \13733 , \13735 );
and \U$13394 ( \13737 , \13730 , \13732 );
or \U$13395 ( \13738 , \13736 , \13737 );
not \U$13396 ( \13739 , \13738 );
or \U$13397 ( \13740 , \13292 , \13739 );
not \U$13398 ( \13741 , \13591 );
not \U$13399 ( \13742 , \13607 );
or \U$13400 ( \13743 , \13741 , \13742 );
or \U$13401 ( \13744 , \13607 , \13591 );
nand \U$13402 ( \13745 , \13743 , \13744 );
not \U$13403 ( \13746 , \13745 );
not \U$13404 ( \13747 , \13589 );
and \U$13405 ( \13748 , \13746 , \13747 );
and \U$13406 ( \13749 , \13745 , \13589 );
nor \U$13407 ( \13750 , \13748 , \13749 );
xor \U$13408 ( \13751 , \13403 , \13489 );
xor \U$13409 ( \13752 , \13751 , \13577 );
or \U$13410 ( \13753 , \13750 , \13752 );
not \U$13411 ( \13754 , \13752 );
not \U$13412 ( \13755 , \13750 );
or \U$13413 ( \13756 , \13754 , \13755 );
xor \U$13414 ( \13757 , \13622 , \13660 );
xor \U$13415 ( \13758 , \13757 , \13673 );
nand \U$13416 ( \13759 , \13756 , \13758 );
nand \U$13417 ( \13760 , \13753 , \13759 );
not \U$13418 ( \13761 , \1128 );
and \U$13419 ( \13762 , \1293 , RI98709c0_97);
and \U$13420 ( \13763 , RI9870e70_107, \1291 );
nor \U$13421 ( \13764 , \13762 , \13763 );
not \U$13422 ( \13765 , \13764 );
or \U$13423 ( \13766 , \13761 , \13765 );
or \U$13424 ( \13767 , \13764 , \1301 );
nand \U$13425 ( \13768 , \13766 , \13767 );
and \U$13426 ( \13769 , \776 , RI9870ab0_99);
and \U$13427 ( \13770 , RI9870d80_105, \774 );
nor \U$13428 ( \13771 , \13769 , \13770 );
and \U$13429 ( \13772 , \13771 , \474 );
not \U$13430 ( \13773 , \13771 );
and \U$13431 ( \13774 , \13773 , \451 );
nor \U$13432 ( \13775 , \13772 , \13774 );
xor \U$13433 ( \13776 , \13768 , \13775 );
and \U$13434 ( \13777 , \1329 , RI9870ba0_101);
and \U$13435 ( \13778 , RI9871050_111, \1327 );
nor \U$13436 ( \13779 , \13777 , \13778 );
and \U$13437 ( \13780 , \13779 , \1336 );
not \U$13438 ( \13781 , \13779 );
and \U$13439 ( \13782 , \13781 , \1337 );
nor \U$13440 ( \13783 , \13780 , \13782 );
and \U$13441 ( \13784 , \13776 , \13783 );
and \U$13442 ( \13785 , \13768 , \13775 );
or \U$13443 ( \13786 , \13784 , \13785 );
not \U$13444 ( \13787 , \456 );
and \U$13445 ( \13788 , \465 , RI986fe80_73);
and \U$13446 ( \13789 , RI9870060_77, \463 );
nor \U$13447 ( \13790 , \13788 , \13789 );
not \U$13448 ( \13791 , \13790 );
or \U$13449 ( \13792 , \13787 , \13791 );
or \U$13450 ( \13793 , \13790 , \454 );
nand \U$13451 ( \13794 , \13792 , \13793 );
and \U$13452 ( \13795 , \438 , RI9870150_79);
and \U$13453 ( \13796 , RI9870f60_109, \436 );
nor \U$13454 ( \13797 , \13795 , \13796 );
and \U$13455 ( \13798 , \13797 , \444 );
not \U$13456 ( \13799 , \13797 );
and \U$13457 ( \13800 , \13799 , \443 );
nor \U$13458 ( \13801 , \13798 , \13800 );
xor \U$13459 ( \13802 , \13794 , \13801 );
not \U$13460 ( \13803 , \367 );
and \U$13461 ( \13804 , \376 , RI986fca0_69);
and \U$13462 ( \13805 , RI986ff70_75, \374 );
nor \U$13463 ( \13806 , \13804 , \13805 );
not \U$13464 ( \13807 , \13806 );
or \U$13465 ( \13808 , \13803 , \13807 );
or \U$13466 ( \13809 , \13806 , \367 );
nand \U$13467 ( \13810 , \13808 , \13809 );
and \U$13468 ( \13811 , \13802 , \13810 );
and \U$13469 ( \13812 , \13794 , \13801 );
or \U$13470 ( \13813 , \13811 , \13812 );
xor \U$13471 ( \13814 , \13786 , \13813 );
and \U$13472 ( \13815 , \2274 , RI9871410_119);
and \U$13473 ( \13816 , RI98716e0_125, \2272 );
nor \U$13474 ( \13817 , \13815 , \13816 );
and \U$13475 ( \13818 , \13817 , \2030 );
not \U$13476 ( \13819 , \13817 );
and \U$13477 ( \13820 , \13819 , \2031 );
nor \U$13478 ( \13821 , \13818 , \13820 );
and \U$13479 ( \13822 , \1311 , RI9870c90_103);
and \U$13480 ( \13823 , RI9871230_115, \1309 );
nor \U$13481 ( \13824 , \13822 , \13823 );
and \U$13482 ( \13825 , \13824 , \1458 );
not \U$13483 ( \13826 , \13824 );
and \U$13484 ( \13827 , \13826 , \1318 );
nor \U$13485 ( \13828 , \13825 , \13827 );
xor \U$13486 ( \13829 , \13821 , \13828 );
not \U$13487 ( \13830 , \2034 );
and \U$13488 ( \13831 , \2042 , RI9871140_113);
and \U$13489 ( \13832 , RI9871320_117, \2040 );
nor \U$13490 ( \13833 , \13831 , \13832 );
not \U$13491 ( \13834 , \13833 );
or \U$13492 ( \13835 , \13830 , \13834 );
or \U$13493 ( \13836 , \13833 , \1462 );
nand \U$13494 ( \13837 , \13835 , \13836 );
and \U$13495 ( \13838 , \13829 , \13837 );
and \U$13496 ( \13839 , \13821 , \13828 );
or \U$13497 ( \13840 , \13838 , \13839 );
and \U$13498 ( \13841 , \13814 , \13840 );
and \U$13499 ( \13842 , \13786 , \13813 );
or \U$13500 ( \13843 , \13841 , \13842 );
and \U$13501 ( \13844 , \8486 , RI986f700_57);
and \U$13502 ( \13845 , RI986f9d0_63, \8484 );
nor \U$13503 ( \13846 , \13844 , \13845 );
and \U$13504 ( \13847 , \13846 , \8050 );
not \U$13505 ( \13848 , \13846 );
and \U$13506 ( \13849 , \13848 , \8051 );
nor \U$13507 ( \13850 , \13847 , \13849 );
and \U$13508 ( \13851 , \7729 , RI986e620_21);
and \U$13509 ( \13852 , RI986f7f0_59, \7727 );
nor \U$13510 ( \13853 , \13851 , \13852 );
and \U$13511 ( \13854 , \13853 , \7480 );
not \U$13512 ( \13855 , \13853 );
and \U$13513 ( \13856 , \13855 , \7733 );
nor \U$13514 ( \13857 , \13854 , \13856 );
xor \U$13515 ( \13858 , \13850 , \13857 );
and \U$13516 ( \13859 , \9237 , RI986f8e0_61);
and \U$13517 ( \13860 , RI986f430_51, \9235 );
nor \U$13518 ( \13861 , \13859 , \13860 );
and \U$13519 ( \13862 , \13861 , \9241 );
not \U$13520 ( \13863 , \13861 );
and \U$13521 ( \13864 , \13863 , \8836 );
nor \U$13522 ( \13865 , \13862 , \13864 );
and \U$13523 ( \13866 , \13858 , \13865 );
and \U$13524 ( \13867 , \13850 , \13857 );
or \U$13525 ( \13868 , \13866 , \13867 );
and \U$13526 ( \13869 , \12293 , RI986dcc0_1);
and \U$13527 ( \13870 , RI986e170_11, \12291 );
nor \U$13528 ( \13871 , \13869 , \13870 );
and \U$13529 ( \13872 , \13871 , \11687 );
not \U$13530 ( \13873 , \13871 );
and \U$13531 ( \13874 , \13873 , \11686 );
nor \U$13532 ( \13875 , \13872 , \13874 );
and \U$13533 ( \13876 , RI98733f0_187, RI9873468_188);
not \U$13534 ( \13877 , RI98734e0_189);
and \U$13535 ( \13878 , \13877 , RI9873468_188);
nor \U$13536 ( \13879 , \13877 , RI9873468_188);
or \U$13537 ( \13880 , \13878 , \13879 );
nor \U$13538 ( \13881 , RI98733f0_187, RI9873468_188);
nor \U$13539 ( \13882 , \13876 , \13880 , \13881 );
nand \U$13540 ( \13883 , RI986e350_15, \13882 );
and \U$13541 ( \13884 , \13883 , \13358 );
not \U$13542 ( \13885 , \13883 );
and \U$13543 ( \13886 , \13885 , \13359 );
nor \U$13544 ( \13887 , \13884 , \13886 );
xor \U$13545 ( \13888 , \13875 , \13887 );
and \U$13546 ( \13889 , \13045 , RI986e080_9);
and \U$13547 ( \13890 , RI986e260_13, \13043 );
nor \U$13548 ( \13891 , \13889 , \13890 );
and \U$13549 ( \13892 , \13891 , \13047 );
not \U$13550 ( \13893 , \13891 );
and \U$13551 ( \13894 , \13893 , \12619 );
nor \U$13552 ( \13895 , \13892 , \13894 );
and \U$13553 ( \13896 , \13888 , \13895 );
and \U$13554 ( \13897 , \13875 , \13887 );
or \U$13555 ( \13898 , \13896 , \13897 );
xor \U$13556 ( \13899 , \13868 , \13898 );
and \U$13557 ( \13900 , \11696 , RI986dea0_5);
and \U$13558 ( \13901 , RI986ddb0_3, \11694 );
nor \U$13559 ( \13902 , \13900 , \13901 );
and \U$13560 ( \13903 , \13902 , \10965 );
not \U$13561 ( \13904 , \13902 );
and \U$13562 ( \13905 , \13904 , \11702 );
nor \U$13563 ( \13906 , \13903 , \13905 );
and \U$13564 ( \13907 , \9505 , RI986f340_49);
and \U$13565 ( \13908 , RI986f520_53, \9503 );
nor \U$13566 ( \13909 , \13907 , \13908 );
and \U$13567 ( \13910 , \13909 , \9510 );
not \U$13568 ( \13911 , \13909 );
and \U$13569 ( \13912 , \13911 , \9513 );
nor \U$13570 ( \13913 , \13910 , \13912 );
xor \U$13571 ( \13914 , \13906 , \13913 );
and \U$13572 ( \13915 , \10424 , RI986f610_55);
and \U$13573 ( \13916 , RI986df90_7, \10422 );
nor \U$13574 ( \13917 , \13915 , \13916 );
and \U$13575 ( \13918 , \13917 , \9840 );
not \U$13576 ( \13919 , \13917 );
and \U$13577 ( \13920 , \13919 , \10428 );
nor \U$13578 ( \13921 , \13918 , \13920 );
and \U$13579 ( \13922 , \13914 , \13921 );
and \U$13580 ( \13923 , \13906 , \13913 );
or \U$13581 ( \13924 , \13922 , \13923 );
and \U$13582 ( \13925 , \13899 , \13924 );
and \U$13583 ( \13926 , \13868 , \13898 );
or \U$13584 ( \13927 , \13925 , \13926 );
xor \U$13585 ( \13928 , \13843 , \13927 );
and \U$13586 ( \13929 , \7079 , RI986e440_17);
and \U$13587 ( \13930 , RI986e710_23, \7077 );
nor \U$13588 ( \13931 , \13929 , \13930 );
and \U$13589 ( \13932 , \13931 , \6710 );
not \U$13590 ( \13933 , \13931 );
and \U$13591 ( \13934 , \13933 , \6709 );
nor \U$13592 ( \13935 , \13932 , \13934 );
and \U$13593 ( \13936 , \5881 , RI986ef80_41);
and \U$13594 ( \13937 , RI986f250_47, \5879 );
nor \U$13595 ( \13938 , \13936 , \13937 );
and \U$13596 ( \13939 , \13938 , \5594 );
not \U$13597 ( \13940 , \13938 );
and \U$13598 ( \13941 , \13940 , \5885 );
nor \U$13599 ( \13942 , \13939 , \13941 );
xor \U$13600 ( \13943 , \13935 , \13942 );
and \U$13601 ( \13944 , \6453 , RI986f160_45);
and \U$13602 ( \13945 , RI986e530_19, \6451 );
nor \U$13603 ( \13946 , \13944 , \13945 );
and \U$13604 ( \13947 , \13946 , \6190 );
not \U$13605 ( \13948 , \13946 );
and \U$13606 ( \13949 , \13948 , \6180 );
nor \U$13607 ( \13950 , \13947 , \13949 );
and \U$13608 ( \13951 , \13943 , \13950 );
and \U$13609 ( \13952 , \13935 , \13942 );
or \U$13610 ( \13953 , \13951 , \13952 );
not \U$13611 ( \13954 , \3406 );
and \U$13612 ( \13955 , \3254 , RI98715f0_123);
and \U$13613 ( \13956 , RI986ead0_31, \3252 );
nor \U$13614 ( \13957 , \13955 , \13956 );
not \U$13615 ( \13958 , \13957 );
or \U$13616 ( \13959 , \13954 , \13958 );
or \U$13617 ( \13960 , \13957 , \2935 );
nand \U$13618 ( \13961 , \13959 , \13960 );
and \U$13619 ( \13962 , \2464 , RI98717d0_127);
and \U$13620 ( \13963 , RI9871500_121, \2462 );
nor \U$13621 ( \13964 , \13962 , \13963 );
and \U$13622 ( \13965 , \13964 , \2468 );
not \U$13623 ( \13966 , \13964 );
and \U$13624 ( \13967 , \13966 , \2263 );
nor \U$13625 ( \13968 , \13965 , \13967 );
xor \U$13626 ( \13969 , \13961 , \13968 );
not \U$13627 ( \13970 , \3918 );
and \U$13628 ( \13971 , \3683 , RI986e9e0_29);
and \U$13629 ( \13972 , RI986e8f0_27, \3681 );
nor \U$13630 ( \13973 , \13971 , \13972 );
not \U$13631 ( \13974 , \13973 );
or \U$13632 ( \13975 , \13970 , \13974 );
or \U$13633 ( \13976 , \13973 , \3918 );
nand \U$13634 ( \13977 , \13975 , \13976 );
and \U$13635 ( \13978 , \13969 , \13977 );
and \U$13636 ( \13979 , \13961 , \13968 );
or \U$13637 ( \13980 , \13978 , \13979 );
xor \U$13638 ( \13981 , \13953 , \13980 );
and \U$13639 ( \13982 , \5318 , RI986ecb0_35);
and \U$13640 ( \13983 , RI986f070_43, \5316 );
nor \U$13641 ( \13984 , \13982 , \13983 );
and \U$13642 ( \13985 , \13984 , \5052 );
not \U$13643 ( \13986 , \13984 );
and \U$13644 ( \13987 , \13986 , \5322 );
nor \U$13645 ( \13988 , \13985 , \13987 );
and \U$13646 ( \13989 , \4203 , RI986e800_25);
and \U$13647 ( \13990 , RI986ee90_39, \4201 );
nor \U$13648 ( \13991 , \13989 , \13990 );
and \U$13649 ( \13992 , \13991 , \4207 );
not \U$13650 ( \13993 , \13991 );
and \U$13651 ( \13994 , \13993 , \3923 );
nor \U$13652 ( \13995 , \13992 , \13994 );
xor \U$13653 ( \13996 , \13988 , \13995 );
not \U$13654 ( \13997 , \4521 );
and \U$13655 ( \13998 , \4710 , RI986eda0_37);
and \U$13656 ( \13999 , RI986ebc0_33, \4708 );
nor \U$13657 ( \14000 , \13998 , \13999 );
not \U$13658 ( \14001 , \14000 );
or \U$13659 ( \14002 , \13997 , \14001 );
or \U$13660 ( \14003 , \14000 , \4521 );
nand \U$13661 ( \14004 , \14002 , \14003 );
and \U$13662 ( \14005 , \13996 , \14004 );
and \U$13663 ( \14006 , \13988 , \13995 );
or \U$13664 ( \14007 , \14005 , \14006 );
and \U$13665 ( \14008 , \13981 , \14007 );
and \U$13666 ( \14009 , \13953 , \13980 );
or \U$13667 ( \14010 , \14008 , \14009 );
and \U$13668 ( \14011 , \13928 , \14010 );
and \U$13669 ( \14012 , \13843 , \13927 );
nor \U$13670 ( \14013 , \14011 , \14012 );
not \U$13671 ( \14014 , \13526 );
not \U$13672 ( \14015 , \13545 );
or \U$13673 ( \14016 , \14014 , \14015 );
or \U$13674 ( \14017 , \13526 , \13545 );
nand \U$13675 ( \14018 , \14016 , \14017 );
not \U$13676 ( \14019 , \14018 );
not \U$13677 ( \14020 , \13534 );
and \U$13678 ( \14021 , \14019 , \14020 );
and \U$13679 ( \14022 , \14018 , \13534 );
nor \U$13680 ( \14023 , \14021 , \14022 );
not \U$13681 ( \14024 , \13505 );
not \U$13682 ( \14025 , \13516 );
or \U$13683 ( \14026 , \14024 , \14025 );
or \U$13684 ( \14027 , \13505 , \13516 );
nand \U$13685 ( \14028 , \14026 , \14027 );
not \U$13686 ( \14029 , \14028 );
not \U$13687 ( \14030 , \13497 );
and \U$13688 ( \14031 , \14029 , \14030 );
and \U$13689 ( \14032 , \14028 , \13497 );
nor \U$13690 ( \14033 , \14031 , \14032 );
or \U$13691 ( \14034 , \14023 , \14033 );
not \U$13692 ( \14035 , \14033 );
not \U$13693 ( \14036 , \14023 );
or \U$13694 ( \14037 , \14035 , \14036 );
xor \U$13695 ( \14038 , \13630 , \13638 );
xor \U$13696 ( \14039 , \14038 , \13646 );
nand \U$13697 ( \14040 , \14037 , \14039 );
nand \U$13698 ( \14041 , \14034 , \14040 );
nand \U$13699 ( \14042 , RI98706f0_91, RI9871fc8_144);
nand \U$13700 ( \14043 , RI9870600_89, RI9871fc8_144);
or \U$13701 ( \14044 , \14042 , \14043 );
not \U$13702 ( \14045 , \14043 );
not \U$13703 ( \14046 , \14042 );
or \U$13704 ( \14047 , \14045 , \14046 );
not \U$13705 ( \14048 , \361 );
and \U$13706 ( \14049 , \354 , RI98707e0_93);
and \U$13707 ( \14050 , RI986fac0_65, \352 );
nor \U$13708 ( \14051 , \14049 , \14050 );
not \U$13709 ( \14052 , \14051 );
or \U$13710 ( \14053 , \14048 , \14052 );
or \U$13711 ( \14054 , \14051 , \361 );
nand \U$13712 ( \14055 , \14053 , \14054 );
not \U$13713 ( \14056 , \386 );
and \U$13714 ( \14057 , \395 , RI986fbb0_67);
and \U$13715 ( \14058 , RI986fd90_71, \393 );
nor \U$13716 ( \14059 , \14057 , \14058 );
not \U$13717 ( \14060 , \14059 );
or \U$13718 ( \14061 , \14056 , \14060 );
or \U$13719 ( \14062 , \14059 , \487 );
nand \U$13720 ( \14063 , \14061 , \14062 );
xor \U$13721 ( \14064 , \14055 , \14063 );
and \U$13722 ( \14065 , \416 , RI9870600_89);
and \U$13723 ( \14066 , RI98708d0_95, \414 );
nor \U$13724 ( \14067 , \14065 , \14066 );
and \U$13725 ( \14068 , \14067 , \422 );
not \U$13726 ( \14069 , \14067 );
and \U$13727 ( \14070 , \14069 , \421 );
nor \U$13728 ( \14071 , \14068 , \14070 );
and \U$13729 ( \14072 , \14064 , \14071 );
and \U$13730 ( \14073 , \14055 , \14063 );
or \U$13731 ( \14074 , \14072 , \14073 );
nand \U$13732 ( \14075 , \14047 , \14074 );
nand \U$13733 ( \14076 , \14044 , \14075 );
xor \U$13734 ( \14077 , \14041 , \14076 );
not \U$13735 ( \14078 , \13472 );
not \U$13736 ( \14079 , \13484 );
or \U$13737 ( \14080 , \14078 , \14079 );
or \U$13738 ( \14081 , \13472 , \13484 );
nand \U$13739 ( \14082 , \14080 , \14081 );
not \U$13740 ( \14083 , \14082 );
not \U$13741 ( \14084 , \13464 );
and \U$13742 ( \14085 , \14083 , \14084 );
and \U$13743 ( \14086 , \14082 , \13464 );
nor \U$13744 ( \14087 , \14085 , \14086 );
not \U$13745 ( \14088 , \13443 );
not \U$13746 ( \14089 , \13454 );
or \U$13747 ( \14090 , \14088 , \14089 );
or \U$13748 ( \14091 , \13443 , \13454 );
nand \U$13749 ( \14092 , \14090 , \14091 );
not \U$13750 ( \14093 , \14092 );
not \U$13751 ( \14094 , \13435 );
and \U$13752 ( \14095 , \14093 , \14094 );
and \U$13753 ( \14096 , \14092 , \13435 );
nor \U$13754 ( \14097 , \14095 , \14096 );
or \U$13755 ( \14098 , \14087 , \14097 );
not \U$13756 ( \14099 , \14097 );
not \U$13757 ( \14100 , \14087 );
or \U$13758 ( \14101 , \14099 , \14100 );
xor \U$13759 ( \14102 , \13555 , \13562 );
xor \U$13760 ( \14103 , \14102 , \13571 );
nand \U$13761 ( \14104 , \14101 , \14103 );
nand \U$13762 ( \14105 , \14098 , \14104 );
and \U$13763 ( \14106 , \14077 , \14105 );
and \U$13764 ( \14107 , \14041 , \14076 );
nor \U$13765 ( \14108 , \14106 , \14107 );
xor \U$13766 ( \14109 , \14013 , \14108 );
xor \U$13767 ( \14110 , \13013 , \13020 );
xor \U$13768 ( \14111 , \14110 , \13028 );
xor \U$13769 ( \14112 , \13597 , \13602 );
xor \U$13770 ( \14113 , \14111 , \14112 );
xor \U$13771 ( \14114 , \13099 , \13106 );
xor \U$13772 ( \14115 , \14114 , \13114 );
xor \U$13773 ( \14116 , \13663 , \13668 );
xor \U$13774 ( \14117 , \14115 , \14116 );
and \U$13775 ( \14118 , \14113 , \14117 );
not \U$13776 ( \14119 , \14113 );
not \U$13777 ( \14120 , \14117 );
and \U$13778 ( \14121 , \14119 , \14120 );
xor \U$13779 ( \14122 , \13410 , \13417 );
xor \U$13780 ( \14123 , \14122 , \13425 );
not \U$13781 ( \14124 , \13334 );
not \U$13782 ( \14125 , \13345 );
or \U$13783 ( \14126 , \14124 , \14125 );
or \U$13784 ( \14127 , \13334 , \13345 );
nand \U$13785 ( \14128 , \14126 , \14127 );
not \U$13786 ( \14129 , \14128 );
not \U$13787 ( \14130 , \13327 );
and \U$13788 ( \14131 , \14129 , \14130 );
and \U$13789 ( \14132 , \14128 , \13327 );
nor \U$13790 ( \14133 , \14131 , \14132 );
xor \U$13791 ( \14134 , \14123 , \14133 );
not \U$13792 ( \14135 , \13387 );
not \U$13793 ( \14136 , \13398 );
or \U$13794 ( \14137 , \14135 , \14136 );
or \U$13795 ( \14138 , \13387 , \13398 );
nand \U$13796 ( \14139 , \14137 , \14138 );
not \U$13797 ( \14140 , \14139 );
not \U$13798 ( \14141 , \13380 );
and \U$13799 ( \14142 , \14140 , \14141 );
and \U$13800 ( \14143 , \14139 , \13380 );
nor \U$13801 ( \14144 , \14142 , \14143 );
and \U$13802 ( \14145 , \14134 , \14144 );
and \U$13803 ( \14146 , \14123 , \14133 );
or \U$13804 ( \14147 , \14145 , \14146 );
nor \U$13805 ( \14148 , \14121 , \14147 );
nor \U$13806 ( \14149 , \14118 , \14148 );
and \U$13807 ( \14150 , \14109 , \14149 );
and \U$13808 ( \14151 , \14013 , \14108 );
nor \U$13809 ( \14152 , \14150 , \14151 );
xor \U$13810 ( \14153 , \13760 , \14152 );
xor \U$13811 ( \14154 , \13518 , \13547 );
xor \U$13812 ( \14155 , \14154 , \13574 );
or \U$13813 ( \14156 , \13659 , \13649 );
nand \U$13814 ( \14157 , \14156 , \13660 );
xor \U$13815 ( \14158 , \14155 , \14157 );
xor \U$13816 ( \14159 , \12984 , \12991 );
xor \U$13817 ( \14160 , \14159 , \13000 );
xor \U$13818 ( \14161 , \13612 , \13617 );
xor \U$13819 ( \14162 , \14160 , \14161 );
and \U$13820 ( \14163 , \14158 , \14162 );
and \U$13821 ( \14164 , \14155 , \14157 );
or \U$13822 ( \14165 , \14163 , \14164 );
xor \U$13823 ( \14166 , \13682 , \13684 );
xor \U$13824 ( \14167 , \14166 , \13687 );
and \U$13825 ( \14168 , \14165 , \14167 );
xor \U$13826 ( \14169 , \13225 , \13227 );
xor \U$13827 ( \14170 , \14169 , \13230 );
xor \U$13828 ( \14171 , \13697 , \13704 );
xor \U$13829 ( \14172 , \14170 , \14171 );
xor \U$13830 ( \14173 , \13682 , \13684 );
xor \U$13831 ( \14174 , \14173 , \13687 );
and \U$13832 ( \14175 , \14172 , \14174 );
and \U$13833 ( \14176 , \14165 , \14172 );
or \U$13834 ( \14177 , \14168 , \14175 , \14176 );
and \U$13835 ( \14178 , \14153 , \14177 );
and \U$13836 ( \14179 , \13760 , \14152 );
or \U$13837 ( \14180 , \14178 , \14179 );
xor \U$13838 ( \14181 , \13190 , \13222 );
xor \U$13839 ( \14182 , \14181 , \13233 );
xor \U$13840 ( \14183 , \13006 , \13091 );
xor \U$13841 ( \14184 , \14183 , \13174 );
xor \U$13842 ( \14185 , \14182 , \14184 );
xor \U$13843 ( \14186 , \12912 , \12914 );
xor \U$13844 ( \14187 , \14186 , \12919 );
xor \U$13845 ( \14188 , \13308 , \13315 );
xor \U$13846 ( \14189 , \14187 , \14188 );
and \U$13847 ( \14190 , \14185 , \14189 );
and \U$13848 ( \14191 , \14182 , \14184 );
or \U$13849 ( \14192 , \14190 , \14191 );
xor \U$13850 ( \14193 , \14180 , \14192 );
xor \U$13851 ( \14194 , \13252 , \13254 );
xor \U$13852 ( \14195 , \14194 , \13259 );
xor \U$13853 ( \14196 , \13294 , \13301 );
xor \U$13854 ( \14197 , \14195 , \14196 );
and \U$13855 ( \14198 , \14193 , \14197 );
and \U$13856 ( \14199 , \14180 , \14192 );
or \U$13857 ( \14200 , \14198 , \14199 );
xor \U$13858 ( \14201 , \12910 , \13239 );
xor \U$13859 ( \14202 , \14201 , \13262 );
xor \U$13860 ( \14203 , \14200 , \14202 );
xor \U$13861 ( \14204 , \13306 , \13715 );
xor \U$13862 ( \14205 , \14204 , \13720 );
and \U$13863 ( \14206 , \14203 , \14205 );
and \U$13864 ( \14207 , \14200 , \14202 );
or \U$13865 ( \14208 , \14206 , \14207 );
xor \U$13866 ( \14209 , \13723 , \13724 );
xor \U$13867 ( \14210 , \14209 , \13727 );
xor \U$13868 ( \14211 , \14208 , \14210 );
not \U$13869 ( \14212 , \14211 );
xor \U$13870 ( \14213 , \13320 , \13679 );
xor \U$13871 ( \14214 , \14213 , \13712 );
xor \U$13872 ( \14215 , \13580 , \13609 );
xor \U$13873 ( \14216 , \14215 , \13676 );
xor \U$13874 ( \14217 , \14182 , \14184 );
xor \U$13875 ( \14218 , \14217 , \14189 );
and \U$13876 ( \14219 , \14216 , \14218 );
xor \U$13877 ( \14220 , \13760 , \14152 );
xor \U$13878 ( \14221 , \14220 , \14177 );
xor \U$13879 ( \14222 , \14182 , \14184 );
xor \U$13880 ( \14223 , \14222 , \14189 );
and \U$13881 ( \14224 , \14221 , \14223 );
and \U$13882 ( \14225 , \14216 , \14221 );
or \U$13883 ( \14226 , \14219 , \14224 , \14225 );
xor \U$13884 ( \14227 , \14214 , \14226 );
xor \U$13885 ( \14228 , \13868 , \13898 );
xor \U$13886 ( \14229 , \14228 , \13924 );
xor \U$13887 ( \14230 , \13786 , \13813 );
xor \U$13888 ( \14231 , \14230 , \13840 );
and \U$13889 ( \14232 , \14229 , \14231 );
xor \U$13890 ( \14233 , \13953 , \13980 );
xor \U$13891 ( \14234 , \14233 , \14007 );
xor \U$13892 ( \14235 , \13786 , \13813 );
xor \U$13893 ( \14236 , \14235 , \13840 );
and \U$13894 ( \14237 , \14234 , \14236 );
and \U$13895 ( \14238 , \14229 , \14234 );
or \U$13896 ( \14239 , \14232 , \14237 , \14238 );
xor \U$13897 ( \14240 , \13428 , \13456 );
xor \U$13898 ( \14241 , \14240 , \13486 );
xor \U$13899 ( \14242 , \14239 , \14241 );
not \U$13900 ( \14243 , \14042 );
not \U$13901 ( \14244 , \14074 );
or \U$13902 ( \14245 , \14243 , \14244 );
or \U$13903 ( \14246 , \14074 , \14042 );
nand \U$13904 ( \14247 , \14245 , \14246 );
not \U$13905 ( \14248 , \14247 );
not \U$13906 ( \14249 , \14043 );
and \U$13907 ( \14250 , \14248 , \14249 );
and \U$13908 ( \14251 , \14247 , \14043 );
nor \U$13909 ( \14252 , \14250 , \14251 );
not \U$13910 ( \14253 , \14039 );
not \U$13911 ( \14254 , \14023 );
or \U$13912 ( \14255 , \14253 , \14254 );
or \U$13913 ( \14256 , \14023 , \14039 );
nand \U$13914 ( \14257 , \14255 , \14256 );
not \U$13915 ( \14258 , \14257 );
not \U$13916 ( \14259 , \14033 );
and \U$13917 ( \14260 , \14258 , \14259 );
and \U$13918 ( \14261 , \14257 , \14033 );
nor \U$13919 ( \14262 , \14260 , \14261 );
xor \U$13920 ( \14263 , \14252 , \14262 );
not \U$13921 ( \14264 , \14097 );
not \U$13922 ( \14265 , \14103 );
or \U$13923 ( \14266 , \14264 , \14265 );
or \U$13924 ( \14267 , \14097 , \14103 );
nand \U$13925 ( \14268 , \14266 , \14267 );
not \U$13926 ( \14269 , \14268 );
not \U$13927 ( \14270 , \14087 );
and \U$13928 ( \14271 , \14269 , \14270 );
and \U$13929 ( \14272 , \14268 , \14087 );
nor \U$13930 ( \14273 , \14271 , \14272 );
and \U$13931 ( \14274 , \14263 , \14273 );
and \U$13932 ( \14275 , \14252 , \14262 );
nor \U$13933 ( \14276 , \14274 , \14275 );
and \U$13934 ( \14277 , \14242 , \14276 );
and \U$13935 ( \14278 , \14239 , \14241 );
or \U$13936 ( \14279 , \14277 , \14278 );
xor \U$13937 ( \14280 , \13988 , \13995 );
xor \U$13938 ( \14281 , \14280 , \14004 );
xor \U$13939 ( \14282 , \13961 , \13968 );
xor \U$13940 ( \14283 , \14282 , \13977 );
and \U$13941 ( \14284 , \14281 , \14283 );
xor \U$13942 ( \14285 , \13935 , \13942 );
xor \U$13943 ( \14286 , \14285 , \13950 );
xor \U$13944 ( \14287 , \13961 , \13968 );
xor \U$13945 ( \14288 , \14287 , \13977 );
and \U$13946 ( \14289 , \14286 , \14288 );
and \U$13947 ( \14290 , \14281 , \14286 );
or \U$13948 ( \14291 , \14284 , \14289 , \14290 );
not \U$13949 ( \14292 , \365 );
and \U$13950 ( \14293 , \376 , RI986fd90_71);
and \U$13951 ( \14294 , RI986fca0_69, \374 );
nor \U$13952 ( \14295 , \14293 , \14294 );
not \U$13953 ( \14296 , \14295 );
or \U$13954 ( \14297 , \14292 , \14296 );
or \U$13955 ( \14298 , \14295 , \365 );
nand \U$13956 ( \14299 , \14297 , \14298 );
not \U$13957 ( \14300 , \487 );
and \U$13958 ( \14301 , \395 , RI986fac0_65);
and \U$13959 ( \14302 , RI986fbb0_67, \393 );
nor \U$13960 ( \14303 , \14301 , \14302 );
not \U$13961 ( \14304 , \14303 );
or \U$13962 ( \14305 , \14300 , \14304 );
or \U$13963 ( \14306 , \14303 , \487 );
nand \U$13964 ( \14307 , \14305 , \14306 );
xor \U$13965 ( \14308 , \14299 , \14307 );
not \U$13966 ( \14309 , \361 );
and \U$13967 ( \14310 , \354 , RI98708d0_95);
and \U$13968 ( \14311 , RI98707e0_93, \352 );
nor \U$13969 ( \14312 , \14310 , \14311 );
not \U$13970 ( \14313 , \14312 );
or \U$13971 ( \14314 , \14309 , \14313 );
or \U$13972 ( \14315 , \14312 , \345 );
nand \U$13973 ( \14316 , \14314 , \14315 );
and \U$13974 ( \14317 , \14308 , \14316 );
and \U$13975 ( \14318 , \14299 , \14307 );
or \U$13976 ( \14319 , \14317 , \14318 );
xor \U$13977 ( \14320 , \14319 , \14042 );
xor \U$13978 ( \14321 , \14055 , \14063 );
xor \U$13979 ( \14322 , \14321 , \14071 );
and \U$13980 ( \14323 , \14320 , \14322 );
and \U$13981 ( \14324 , \14319 , \14042 );
or \U$13982 ( \14325 , \14323 , \14324 );
xor \U$13983 ( \14326 , \14291 , \14325 );
xor \U$13984 ( \14327 , \13821 , \13828 );
xor \U$13985 ( \14328 , \14327 , \13837 );
xor \U$13986 ( \14329 , \13794 , \13801 );
xor \U$13987 ( \14330 , \14329 , \13810 );
xor \U$13988 ( \14331 , \14328 , \14330 );
xor \U$13989 ( \14332 , \13768 , \13775 );
xor \U$13990 ( \14333 , \14332 , \13783 );
and \U$13991 ( \14334 , \14331 , \14333 );
and \U$13992 ( \14335 , \14328 , \14330 );
or \U$13993 ( \14336 , \14334 , \14335 );
and \U$13994 ( \14337 , \14326 , \14336 );
and \U$13995 ( \14338 , \14291 , \14325 );
or \U$13996 ( \14339 , \14337 , \14338 );
and \U$13997 ( \14340 , \7729 , RI986e710_23);
and \U$13998 ( \14341 , RI986e620_21, \7727 );
nor \U$13999 ( \14342 , \14340 , \14341 );
and \U$14000 ( \14343 , \14342 , \7480 );
not \U$14001 ( \14344 , \14342 );
and \U$14002 ( \14345 , \14344 , \7733 );
nor \U$14003 ( \14346 , \14343 , \14345 );
and \U$14004 ( \14347 , \6453 , RI986f250_47);
and \U$14005 ( \14348 , RI986f160_45, \6451 );
nor \U$14006 ( \14349 , \14347 , \14348 );
and \U$14007 ( \14350 , \14349 , \6190 );
not \U$14008 ( \14351 , \14349 );
and \U$14009 ( \14352 , \14351 , \6705 );
nor \U$14010 ( \14353 , \14350 , \14352 );
xor \U$14011 ( \14354 , \14346 , \14353 );
and \U$14012 ( \14355 , \7079 , RI986e530_19);
and \U$14013 ( \14356 , RI986e440_17, \7077 );
nor \U$14014 ( \14357 , \14355 , \14356 );
and \U$14015 ( \14358 , \14357 , \6710 );
not \U$14016 ( \14359 , \14357 );
and \U$14017 ( \14360 , \14359 , \6709 );
nor \U$14018 ( \14361 , \14358 , \14360 );
and \U$14019 ( \14362 , \14354 , \14361 );
and \U$14020 ( \14363 , \14346 , \14353 );
or \U$14021 ( \14364 , \14362 , \14363 );
not \U$14022 ( \14365 , \3406 );
and \U$14023 ( \14366 , \3254 , RI9871500_121);
and \U$14024 ( \14367 , RI98715f0_123, \3252 );
nor \U$14025 ( \14368 , \14366 , \14367 );
not \U$14026 ( \14369 , \14368 );
or \U$14027 ( \14370 , \14365 , \14369 );
or \U$14028 ( \14371 , \14368 , \3406 );
nand \U$14029 ( \14372 , \14370 , \14371 );
not \U$14030 ( \14373 , \3918 );
and \U$14031 ( \14374 , \3683 , RI986ead0_31);
and \U$14032 ( \14375 , RI986e9e0_29, \3681 );
nor \U$14033 ( \14376 , \14374 , \14375 );
not \U$14034 ( \14377 , \14376 );
or \U$14035 ( \14378 , \14373 , \14377 );
or \U$14036 ( \14379 , \14376 , \3412 );
nand \U$14037 ( \14380 , \14378 , \14379 );
xor \U$14038 ( \14381 , \14372 , \14380 );
and \U$14039 ( \14382 , \4203 , RI986e8f0_27);
and \U$14040 ( \14383 , RI986e800_25, \4201 );
nor \U$14041 ( \14384 , \14382 , \14383 );
and \U$14042 ( \14385 , \14384 , \4207 );
not \U$14043 ( \14386 , \14384 );
and \U$14044 ( \14387 , \14386 , \3922 );
nor \U$14045 ( \14388 , \14385 , \14387 );
and \U$14046 ( \14389 , \14381 , \14388 );
and \U$14047 ( \14390 , \14372 , \14380 );
or \U$14048 ( \14391 , \14389 , \14390 );
xor \U$14049 ( \14392 , \14364 , \14391 );
and \U$14050 ( \14393 , \5881 , RI986f070_43);
and \U$14051 ( \14394 , RI986ef80_41, \5879 );
nor \U$14052 ( \14395 , \14393 , \14394 );
and \U$14053 ( \14396 , \14395 , \5594 );
not \U$14054 ( \14397 , \14395 );
and \U$14055 ( \14398 , \14397 , \5885 );
nor \U$14056 ( \14399 , \14396 , \14398 );
not \U$14057 ( \14400 , \4519 );
and \U$14058 ( \14401 , \4710 , RI986ee90_39);
and \U$14059 ( \14402 , RI986eda0_37, \4708 );
nor \U$14060 ( \14403 , \14401 , \14402 );
not \U$14061 ( \14404 , \14403 );
or \U$14062 ( \14405 , \14400 , \14404 );
or \U$14063 ( \14406 , \14403 , \4521 );
nand \U$14064 ( \14407 , \14405 , \14406 );
xor \U$14065 ( \14408 , \14399 , \14407 );
and \U$14066 ( \14409 , \5318 , RI986ebc0_33);
and \U$14067 ( \14410 , RI986ecb0_35, \5316 );
nor \U$14068 ( \14411 , \14409 , \14410 );
and \U$14069 ( \14412 , \14411 , \5052 );
not \U$14070 ( \14413 , \14411 );
and \U$14071 ( \14414 , \14413 , \5322 );
nor \U$14072 ( \14415 , \14412 , \14414 );
and \U$14073 ( \14416 , \14408 , \14415 );
and \U$14074 ( \14417 , \14399 , \14407 );
or \U$14075 ( \14418 , \14416 , \14417 );
and \U$14076 ( \14419 , \14392 , \14418 );
and \U$14077 ( \14420 , \14364 , \14391 );
or \U$14078 ( \14421 , \14419 , \14420 );
and \U$14079 ( \14422 , \1329 , RI9870e70_107);
and \U$14080 ( \14423 , RI9870ba0_101, \1327 );
nor \U$14081 ( \14424 , \14422 , \14423 );
and \U$14082 ( \14425 , \14424 , \1336 );
not \U$14083 ( \14426 , \14424 );
and \U$14084 ( \14427 , \14426 , \1337 );
nor \U$14085 ( \14428 , \14425 , \14427 );
not \U$14086 ( \14429 , \1128 );
and \U$14087 ( \14430 , \1293 , RI9870d80_105);
and \U$14088 ( \14431 , RI98709c0_97, \1291 );
nor \U$14089 ( \14432 , \14430 , \14431 );
not \U$14090 ( \14433 , \14432 );
or \U$14091 ( \14434 , \14429 , \14433 );
or \U$14092 ( \14435 , \14432 , \1128 );
nand \U$14093 ( \14436 , \14434 , \14435 );
xor \U$14094 ( \14437 , \14428 , \14436 );
and \U$14095 ( \14438 , \1311 , RI9871050_111);
and \U$14096 ( \14439 , RI9870c90_103, \1309 );
nor \U$14097 ( \14440 , \14438 , \14439 );
and \U$14098 ( \14441 , \14440 , \1458 );
not \U$14099 ( \14442 , \14440 );
and \U$14100 ( \14443 , \14442 , \1315 );
nor \U$14101 ( \14444 , \14441 , \14443 );
and \U$14102 ( \14445 , \14437 , \14444 );
and \U$14103 ( \14446 , \14428 , \14436 );
or \U$14104 ( \14447 , \14445 , \14446 );
and \U$14105 ( \14448 , \438 , RI9870060_77);
and \U$14106 ( \14449 , RI9870150_79, \436 );
nor \U$14107 ( \14450 , \14448 , \14449 );
and \U$14108 ( \14451 , \14450 , \444 );
not \U$14109 ( \14452 , \14450 );
and \U$14110 ( \14453 , \14452 , \443 );
nor \U$14111 ( \14454 , \14451 , \14453 );
and \U$14112 ( \14455 , \776 , RI9870f60_109);
and \U$14113 ( \14456 , RI9870ab0_99, \774 );
nor \U$14114 ( \14457 , \14455 , \14456 );
and \U$14115 ( \14458 , \14457 , \474 );
not \U$14116 ( \14459 , \14457 );
and \U$14117 ( \14460 , \14459 , \451 );
nor \U$14118 ( \14461 , \14458 , \14460 );
xor \U$14119 ( \14462 , \14454 , \14461 );
not \U$14120 ( \14463 , \454 );
and \U$14121 ( \14464 , \465 , RI986ff70_75);
and \U$14122 ( \14465 , RI986fe80_73, \463 );
nor \U$14123 ( \14466 , \14464 , \14465 );
not \U$14124 ( \14467 , \14466 );
or \U$14125 ( \14468 , \14463 , \14467 );
or \U$14126 ( \14469 , \14466 , \456 );
nand \U$14127 ( \14470 , \14468 , \14469 );
and \U$14128 ( \14471 , \14462 , \14470 );
and \U$14129 ( \14472 , \14454 , \14461 );
or \U$14130 ( \14473 , \14471 , \14472 );
xor \U$14131 ( \14474 , \14447 , \14473 );
and \U$14132 ( \14475 , \2464 , RI98716e0_125);
and \U$14133 ( \14476 , RI98717d0_127, \2462 );
nor \U$14134 ( \14477 , \14475 , \14476 );
and \U$14135 ( \14478 , \14477 , \2468 );
not \U$14136 ( \14479 , \14477 );
and \U$14137 ( \14480 , \14479 , \2263 );
nor \U$14138 ( \14481 , \14478 , \14480 );
not \U$14139 ( \14482 , \2034 );
and \U$14140 ( \14483 , \2042 , RI9871230_115);
and \U$14141 ( \14484 , RI9871140_113, \2040 );
nor \U$14142 ( \14485 , \14483 , \14484 );
not \U$14143 ( \14486 , \14485 );
or \U$14144 ( \14487 , \14482 , \14486 );
or \U$14145 ( \14488 , \14485 , \2034 );
nand \U$14146 ( \14489 , \14487 , \14488 );
xor \U$14147 ( \14490 , \14481 , \14489 );
and \U$14148 ( \14491 , \2274 , RI9871320_117);
and \U$14149 ( \14492 , RI9871410_119, \2272 );
nor \U$14150 ( \14493 , \14491 , \14492 );
and \U$14151 ( \14494 , \14493 , \2030 );
not \U$14152 ( \14495 , \14493 );
and \U$14153 ( \14496 , \14495 , \2031 );
nor \U$14154 ( \14497 , \14494 , \14496 );
and \U$14155 ( \14498 , \14490 , \14497 );
and \U$14156 ( \14499 , \14481 , \14489 );
or \U$14157 ( \14500 , \14498 , \14499 );
and \U$14158 ( \14501 , \14474 , \14500 );
and \U$14159 ( \14502 , \14447 , \14473 );
or \U$14160 ( \14503 , \14501 , \14502 );
xor \U$14161 ( \14504 , \14421 , \14503 );
and \U$14162 ( \14505 , \9505 , RI986f430_51);
and \U$14163 ( \14506 , RI986f340_49, \9503 );
nor \U$14164 ( \14507 , \14505 , \14506 );
and \U$14165 ( \14508 , \14507 , \9510 );
not \U$14166 ( \14509 , \14507 );
and \U$14167 ( \14510 , \14509 , \9513 );
nor \U$14168 ( \14511 , \14508 , \14510 );
and \U$14169 ( \14512 , \8486 , RI986f7f0_59);
and \U$14170 ( \14513 , RI986f700_57, \8484 );
nor \U$14171 ( \14514 , \14512 , \14513 );
and \U$14172 ( \14515 , \14514 , \8050 );
not \U$14173 ( \14516 , \14514 );
and \U$14174 ( \14517 , \14516 , \8051 );
nor \U$14175 ( \14518 , \14515 , \14517 );
xor \U$14176 ( \14519 , \14511 , \14518 );
and \U$14177 ( \14520 , \9237 , RI986f9d0_63);
and \U$14178 ( \14521 , RI986f8e0_61, \9235 );
nor \U$14179 ( \14522 , \14520 , \14521 );
and \U$14180 ( \14523 , \14522 , \9241 );
not \U$14181 ( \14524 , \14522 );
and \U$14182 ( \14525 , \14524 , \8836 );
nor \U$14183 ( \14526 , \14523 , \14525 );
and \U$14184 ( \14527 , \14519 , \14526 );
and \U$14185 ( \14528 , \14511 , \14518 );
or \U$14186 ( \14529 , \14527 , \14528 );
and \U$14187 ( \14530 , \13882 , RI986e260_13);
and \U$14188 ( \14531 , RI986e350_15, \13880 );
nor \U$14189 ( \14532 , \14530 , \14531 );
and \U$14190 ( \14533 , \14532 , \13358 );
not \U$14191 ( \14534 , \14532 );
and \U$14192 ( \14535 , \14534 , \13359 );
nor \U$14193 ( \14536 , \14533 , \14535 );
nand \U$14194 ( \14537 , RI9873558_190, RI98735d0_191);
and \U$14195 ( \14538 , \14537 , RI98734e0_189);
not \U$14196 ( \14539 , \14538 );
xor \U$14197 ( \14540 , \14536 , \14539 );
and \U$14198 ( \14541 , \13045 , RI986e170_11);
and \U$14199 ( \14542 , RI986e080_9, \13043 );
nor \U$14200 ( \14543 , \14541 , \14542 );
and \U$14201 ( \14544 , \14543 , \13047 );
not \U$14202 ( \14545 , \14543 );
and \U$14203 ( \14546 , \14545 , \12619 );
nor \U$14204 ( \14547 , \14544 , \14546 );
and \U$14205 ( \14548 , \14540 , \14547 );
and \U$14206 ( \14549 , \14536 , \14539 );
or \U$14207 ( \14550 , \14548 , \14549 );
xor \U$14208 ( \14551 , \14529 , \14550 );
and \U$14209 ( \14552 , \10424 , RI986f520_53);
and \U$14210 ( \14553 , RI986f610_55, \10422 );
nor \U$14211 ( \14554 , \14552 , \14553 );
and \U$14212 ( \14555 , \14554 , \9840 );
not \U$14213 ( \14556 , \14554 );
and \U$14214 ( \14557 , \14556 , \10428 );
nor \U$14215 ( \14558 , \14555 , \14557 );
and \U$14216 ( \14559 , \11696 , RI986df90_7);
and \U$14217 ( \14560 , RI986dea0_5, \11694 );
nor \U$14218 ( \14561 , \14559 , \14560 );
and \U$14219 ( \14562 , \14561 , \10965 );
not \U$14220 ( \14563 , \14561 );
and \U$14221 ( \14564 , \14563 , \11702 );
nor \U$14222 ( \14565 , \14562 , \14564 );
xor \U$14223 ( \14566 , \14558 , \14565 );
and \U$14224 ( \14567 , \12293 , RI986ddb0_3);
and \U$14225 ( \14568 , RI986dcc0_1, \12291 );
nor \U$14226 ( \14569 , \14567 , \14568 );
and \U$14227 ( \14570 , \14569 , \11687 );
not \U$14228 ( \14571 , \14569 );
and \U$14229 ( \14572 , \14571 , \11686 );
nor \U$14230 ( \14573 , \14570 , \14572 );
and \U$14231 ( \14574 , \14566 , \14573 );
and \U$14232 ( \14575 , \14558 , \14565 );
or \U$14233 ( \14576 , \14574 , \14575 );
and \U$14234 ( \14577 , \14551 , \14576 );
and \U$14235 ( \14578 , \14529 , \14550 );
or \U$14236 ( \14579 , \14577 , \14578 );
and \U$14237 ( \14580 , \14504 , \14579 );
and \U$14238 ( \14581 , \14421 , \14503 );
or \U$14239 ( \14582 , \14580 , \14581 );
xor \U$14240 ( \14583 , \14339 , \14582 );
xor \U$14241 ( \14584 , \14123 , \14133 );
xor \U$14242 ( \14585 , \14584 , \14144 );
and \U$14243 ( \14586 , \13370 , \13358 );
not \U$14244 ( \14587 , \13370 );
and \U$14245 ( \14588 , \14587 , \13359 );
nor \U$14246 ( \14589 , \14586 , \14588 );
not \U$14247 ( \14590 , \14589 );
not \U$14248 ( \14591 , \13354 );
and \U$14249 ( \14592 , \14590 , \14591 );
and \U$14250 ( \14593 , \14589 , \13354 );
nor \U$14251 ( \14594 , \14592 , \14593 );
or \U$14252 ( \14595 , \14585 , \14594 );
not \U$14253 ( \14596 , \14594 );
not \U$14254 ( \14597 , \14585 );
or \U$14255 ( \14598 , \14596 , \14597 );
xor \U$14256 ( \14599 , \13850 , \13857 );
xor \U$14257 ( \14600 , \14599 , \13865 );
xor \U$14258 ( \14601 , \13875 , \13887 );
xor \U$14259 ( \14602 , \14601 , \13895 );
and \U$14260 ( \14603 , \14600 , \14602 );
xor \U$14261 ( \14604 , \13906 , \13913 );
xor \U$14262 ( \14605 , \14604 , \13921 );
xor \U$14263 ( \14606 , \13875 , \13887 );
xor \U$14264 ( \14607 , \14606 , \13895 );
and \U$14265 ( \14608 , \14605 , \14607 );
and \U$14266 ( \14609 , \14600 , \14605 );
or \U$14267 ( \14610 , \14603 , \14608 , \14609 );
nand \U$14268 ( \14611 , \14598 , \14610 );
nand \U$14269 ( \14612 , \14595 , \14611 );
and \U$14270 ( \14613 , \14583 , \14612 );
and \U$14271 ( \14614 , \14339 , \14582 );
or \U$14272 ( \14615 , \14613 , \14614 );
xor \U$14273 ( \14616 , \14279 , \14615 );
xor \U$14274 ( \14617 , \13347 , \13372 );
xor \U$14275 ( \14618 , \14617 , \13400 );
xor \U$14276 ( \14619 , \14155 , \14157 );
xor \U$14277 ( \14620 , \14619 , \14162 );
and \U$14278 ( \14621 , \14618 , \14620 );
not \U$14279 ( \14622 , \14147 );
not \U$14280 ( \14623 , \14113 );
or \U$14281 ( \14624 , \14622 , \14623 );
or \U$14282 ( \14625 , \14113 , \14147 );
nand \U$14283 ( \14626 , \14624 , \14625 );
xor \U$14284 ( \14627 , \14117 , \14626 );
xor \U$14285 ( \14628 , \14155 , \14157 );
xor \U$14286 ( \14629 , \14628 , \14162 );
and \U$14287 ( \14630 , \14627 , \14629 );
and \U$14288 ( \14631 , \14618 , \14627 );
or \U$14289 ( \14632 , \14621 , \14630 , \14631 );
and \U$14290 ( \14633 , \14616 , \14632 );
and \U$14291 ( \14634 , \14279 , \14615 );
or \U$14292 ( \14635 , \14633 , \14634 );
xor \U$14293 ( \14636 , \13690 , \13692 );
xor \U$14294 ( \14637 , \14636 , \13709 );
xor \U$14295 ( \14638 , \14635 , \14637 );
not \U$14296 ( \14639 , \13752 );
not \U$14297 ( \14640 , \13758 );
or \U$14298 ( \14641 , \14639 , \14640 );
or \U$14299 ( \14642 , \13758 , \13752 );
nand \U$14300 ( \14643 , \14641 , \14642 );
not \U$14301 ( \14644 , \14643 );
not \U$14302 ( \14645 , \13750 );
and \U$14303 ( \14646 , \14644 , \14645 );
and \U$14304 ( \14647 , \14643 , \13750 );
nor \U$14305 ( \14648 , \14646 , \14647 );
xor \U$14306 ( \14649 , \14013 , \14108 );
xor \U$14307 ( \14650 , \14649 , \14149 );
or \U$14308 ( \14651 , \14648 , \14650 );
not \U$14309 ( \14652 , \14650 );
not \U$14310 ( \14653 , \14648 );
or \U$14311 ( \14654 , \14652 , \14653 );
xor \U$14312 ( \14655 , \13682 , \13684 );
xor \U$14313 ( \14656 , \14655 , \13687 );
xor \U$14314 ( \14657 , \14165 , \14172 );
xor \U$14315 ( \14658 , \14656 , \14657 );
nand \U$14316 ( \14659 , \14654 , \14658 );
nand \U$14317 ( \14660 , \14651 , \14659 );
and \U$14318 ( \14661 , \14638 , \14660 );
and \U$14319 ( \14662 , \14635 , \14637 );
or \U$14320 ( \14663 , \14661 , \14662 );
and \U$14321 ( \14664 , \14227 , \14663 );
and \U$14322 ( \14665 , \14214 , \14226 );
nor \U$14323 ( \14666 , \14664 , \14665 );
not \U$14324 ( \14667 , \14666 );
xor \U$14325 ( \14668 , \14200 , \14202 );
xor \U$14326 ( \14669 , \14668 , \14205 );
nand \U$14327 ( \14670 , \14667 , \14669 );
or \U$14328 ( \14671 , \14212 , \14670 );
not \U$14329 ( \14672 , \14211 );
not \U$14330 ( \14673 , \14670 );
and \U$14331 ( \14674 , \14672 , \14673 );
and \U$14332 ( \14675 , \14211 , \14670 );
nor \U$14333 ( \14676 , \14674 , \14675 );
xor \U$14334 ( \14677 , \14182 , \14184 );
xor \U$14335 ( \14678 , \14677 , \14189 );
xor \U$14336 ( \14679 , \14216 , \14221 );
xor \U$14337 ( \14680 , \14678 , \14679 );
not \U$14338 ( \14681 , \14680 );
xor \U$14339 ( \14682 , \14635 , \14637 );
xor \U$14340 ( \14683 , \14682 , \14660 );
not \U$14341 ( \14684 , \14683 );
or \U$14342 ( \14685 , \14681 , \14684 );
or \U$14343 ( \14686 , \14683 , \14680 );
xnor \U$14344 ( \14687 , \14650 , \14648 );
not \U$14345 ( \14688 , \14687 );
not \U$14346 ( \14689 , \14658 );
and \U$14347 ( \14690 , \14688 , \14689 );
and \U$14348 ( \14691 , \14687 , \14658 );
nor \U$14349 ( \14692 , \14690 , \14691 );
not \U$14350 ( \14693 , \14692 );
xor \U$14351 ( \14694 , \13843 , \13927 );
xor \U$14352 ( \14695 , \14694 , \14010 );
xor \U$14353 ( \14696 , \14041 , \14076 );
xor \U$14354 ( \14697 , \14696 , \14105 );
xor \U$14355 ( \14698 , \14695 , \14697 );
xor \U$14356 ( \14699 , \14155 , \14157 );
xor \U$14357 ( \14700 , \14699 , \14162 );
xor \U$14358 ( \14701 , \14618 , \14627 );
xor \U$14359 ( \14702 , \14700 , \14701 );
and \U$14360 ( \14703 , \14698 , \14702 );
and \U$14361 ( \14704 , \14695 , \14697 );
nor \U$14362 ( \14705 , \14703 , \14704 );
not \U$14363 ( \14706 , \14705 );
and \U$14364 ( \14707 , \14693 , \14706 );
and \U$14365 ( \14708 , \14692 , \14705 );
xor \U$14366 ( \14709 , \14319 , \14042 );
xor \U$14367 ( \14710 , \14709 , \14322 );
xor \U$14368 ( \14711 , \14328 , \14330 );
xor \U$14369 ( \14712 , \14711 , \14333 );
and \U$14370 ( \14713 , \14710 , \14712 );
xor \U$14371 ( \14714 , \13961 , \13968 );
xor \U$14372 ( \14715 , \14714 , \13977 );
xor \U$14373 ( \14716 , \14281 , \14286 );
xor \U$14374 ( \14717 , \14715 , \14716 );
xor \U$14375 ( \14718 , \14328 , \14330 );
xor \U$14376 ( \14719 , \14718 , \14333 );
and \U$14377 ( \14720 , \14717 , \14719 );
and \U$14378 ( \14721 , \14710 , \14717 );
or \U$14379 ( \14722 , \14713 , \14720 , \14721 );
xor \U$14380 ( \14723 , \14447 , \14473 );
xor \U$14381 ( \14724 , \14723 , \14500 );
xor \U$14382 ( \14725 , \14529 , \14550 );
xor \U$14383 ( \14726 , \14725 , \14576 );
and \U$14384 ( \14727 , \14724 , \14726 );
xor \U$14385 ( \14728 , \14364 , \14391 );
xor \U$14386 ( \14729 , \14728 , \14418 );
xor \U$14387 ( \14730 , \14529 , \14550 );
xor \U$14388 ( \14731 , \14730 , \14576 );
and \U$14389 ( \14732 , \14729 , \14731 );
and \U$14390 ( \14733 , \14724 , \14729 );
or \U$14391 ( \14734 , \14727 , \14732 , \14733 );
xor \U$14392 ( \14735 , \14722 , \14734 );
xor \U$14393 ( \14736 , \13786 , \13813 );
xor \U$14394 ( \14737 , \14736 , \13840 );
xor \U$14395 ( \14738 , \14229 , \14234 );
xor \U$14396 ( \14739 , \14737 , \14738 );
and \U$14397 ( \14740 , \14735 , \14739 );
and \U$14398 ( \14741 , \14722 , \14734 );
or \U$14399 ( \14742 , \14740 , \14741 );
not \U$14400 ( \14743 , RI9870240_81);
nor \U$14401 ( \14744 , \14743 , \407 );
xor \U$14402 ( \14745 , \14299 , \14307 );
xor \U$14403 ( \14746 , \14745 , \14316 );
and \U$14404 ( \14747 , \14744 , \14746 );
xor \U$14405 ( \14748 , \14454 , \14461 );
xor \U$14406 ( \14749 , \14748 , \14470 );
xor \U$14407 ( \14750 , \14299 , \14307 );
xor \U$14408 ( \14751 , \14750 , \14316 );
and \U$14409 ( \14752 , \14749 , \14751 );
and \U$14410 ( \14753 , \14744 , \14749 );
or \U$14411 ( \14754 , \14747 , \14752 , \14753 );
nand \U$14412 ( \14755 , RI9870330_83, RI9871fc8_144);
and \U$14413 ( \14756 , \416 , RI9870240_81);
and \U$14414 ( \14757 , RI98706f0_91, \414 );
nor \U$14415 ( \14758 , \14756 , \14757 );
and \U$14416 ( \14759 , \14758 , \421 );
not \U$14417 ( \14760 , \14758 );
and \U$14418 ( \14761 , \14760 , \422 );
nor \U$14419 ( \14762 , \14759 , \14761 );
nand \U$14420 ( \14763 , \14755 , \14762 );
and \U$14421 ( \14764 , \416 , RI98706f0_91);
and \U$14422 ( \14765 , RI9870600_89, \414 );
nor \U$14423 ( \14766 , \14764 , \14765 );
and \U$14424 ( \14767 , \14766 , \422 );
not \U$14425 ( \14768 , \14766 );
and \U$14426 ( \14769 , \14768 , \421 );
nor \U$14427 ( \14770 , \14767 , \14769 );
xor \U$14428 ( \14771 , \14763 , \14770 );
not \U$14429 ( \14772 , \487 );
and \U$14430 ( \14773 , \395 , RI98707e0_93);
and \U$14431 ( \14774 , RI986fac0_65, \393 );
nor \U$14432 ( \14775 , \14773 , \14774 );
not \U$14433 ( \14776 , \14775 );
or \U$14434 ( \14777 , \14772 , \14776 );
or \U$14435 ( \14778 , \14775 , \487 );
nand \U$14436 ( \14779 , \14777 , \14778 );
not \U$14437 ( \14780 , \367 );
and \U$14438 ( \14781 , \376 , RI986fbb0_67);
and \U$14439 ( \14782 , RI986fd90_71, \374 );
nor \U$14440 ( \14783 , \14781 , \14782 );
not \U$14441 ( \14784 , \14783 );
or \U$14442 ( \14785 , \14780 , \14784 );
or \U$14443 ( \14786 , \14783 , \367 );
nand \U$14444 ( \14787 , \14785 , \14786 );
xor \U$14445 ( \14788 , \14779 , \14787 );
not \U$14446 ( \14789 , \345 );
and \U$14447 ( \14790 , \354 , RI9870600_89);
and \U$14448 ( \14791 , RI98708d0_95, \352 );
nor \U$14449 ( \14792 , \14790 , \14791 );
not \U$14450 ( \14793 , \14792 );
or \U$14451 ( \14794 , \14789 , \14793 );
or \U$14452 ( \14795 , \14792 , \345 );
nand \U$14453 ( \14796 , \14794 , \14795 );
and \U$14454 ( \14797 , \14788 , \14796 );
and \U$14455 ( \14798 , \14779 , \14787 );
or \U$14456 ( \14799 , \14797 , \14798 );
and \U$14457 ( \14800 , \14771 , \14799 );
and \U$14458 ( \14801 , \14763 , \14770 );
or \U$14459 ( \14802 , \14800 , \14801 );
xor \U$14460 ( \14803 , \14754 , \14802 );
xor \U$14461 ( \14804 , \14481 , \14489 );
xor \U$14462 ( \14805 , \14804 , \14497 );
xor \U$14463 ( \14806 , \14428 , \14436 );
xor \U$14464 ( \14807 , \14806 , \14444 );
xor \U$14465 ( \14808 , \14805 , \14807 );
xor \U$14466 ( \14809 , \14372 , \14380 );
xor \U$14467 ( \14810 , \14809 , \14388 );
and \U$14468 ( \14811 , \14808 , \14810 );
and \U$14469 ( \14812 , \14805 , \14807 );
or \U$14470 ( \14813 , \14811 , \14812 );
and \U$14471 ( \14814 , \14803 , \14813 );
and \U$14472 ( \14815 , \14754 , \14802 );
or \U$14473 ( \14816 , \14814 , \14815 );
and \U$14474 ( \14817 , \1329 , RI98709c0_97);
and \U$14475 ( \14818 , RI9870e70_107, \1327 );
nor \U$14476 ( \14819 , \14817 , \14818 );
and \U$14477 ( \14820 , \14819 , \1336 );
not \U$14478 ( \14821 , \14819 );
and \U$14479 ( \14822 , \14821 , \1337 );
nor \U$14480 ( \14823 , \14820 , \14822 );
not \U$14481 ( \14824 , \1301 );
and \U$14482 ( \14825 , \1293 , RI9870ab0_99);
and \U$14483 ( \14826 , RI9870d80_105, \1291 );
nor \U$14484 ( \14827 , \14825 , \14826 );
not \U$14485 ( \14828 , \14827 );
or \U$14486 ( \14829 , \14824 , \14828 );
or \U$14487 ( \14830 , \14827 , \1301 );
nand \U$14488 ( \14831 , \14829 , \14830 );
xor \U$14489 ( \14832 , \14823 , \14831 );
and \U$14490 ( \14833 , \1311 , RI9870ba0_101);
and \U$14491 ( \14834 , RI9871050_111, \1309 );
nor \U$14492 ( \14835 , \14833 , \14834 );
and \U$14493 ( \14836 , \14835 , \1458 );
not \U$14494 ( \14837 , \14835 );
and \U$14495 ( \14838 , \14837 , \1318 );
nor \U$14496 ( \14839 , \14836 , \14838 );
and \U$14497 ( \14840 , \14832 , \14839 );
and \U$14498 ( \14841 , \14823 , \14831 );
or \U$14499 ( \14842 , \14840 , \14841 );
and \U$14500 ( \14843 , \776 , RI9870150_79);
and \U$14501 ( \14844 , RI9870f60_109, \774 );
nor \U$14502 ( \14845 , \14843 , \14844 );
and \U$14503 ( \14846 , \14845 , \474 );
not \U$14504 ( \14847 , \14845 );
and \U$14505 ( \14848 , \14847 , \451 );
nor \U$14506 ( \14849 , \14846 , \14848 );
and \U$14507 ( \14850 , \438 , RI986fe80_73);
and \U$14508 ( \14851 , RI9870060_77, \436 );
nor \U$14509 ( \14852 , \14850 , \14851 );
and \U$14510 ( \14853 , \14852 , \444 );
not \U$14511 ( \14854 , \14852 );
and \U$14512 ( \14855 , \14854 , \443 );
nor \U$14513 ( \14856 , \14853 , \14855 );
xor \U$14514 ( \14857 , \14849 , \14856 );
not \U$14515 ( \14858 , \456 );
and \U$14516 ( \14859 , \465 , RI986fca0_69);
and \U$14517 ( \14860 , RI986ff70_75, \463 );
nor \U$14518 ( \14861 , \14859 , \14860 );
not \U$14519 ( \14862 , \14861 );
or \U$14520 ( \14863 , \14858 , \14862 );
or \U$14521 ( \14864 , \14861 , \456 );
nand \U$14522 ( \14865 , \14863 , \14864 );
and \U$14523 ( \14866 , \14857 , \14865 );
and \U$14524 ( \14867 , \14849 , \14856 );
or \U$14525 ( \14868 , \14866 , \14867 );
xor \U$14526 ( \14869 , \14842 , \14868 );
and \U$14527 ( \14870 , \2274 , RI9871140_113);
and \U$14528 ( \14871 , RI9871320_117, \2272 );
nor \U$14529 ( \14872 , \14870 , \14871 );
and \U$14530 ( \14873 , \14872 , \2030 );
not \U$14531 ( \14874 , \14872 );
and \U$14532 ( \14875 , \14874 , \2031 );
nor \U$14533 ( \14876 , \14873 , \14875 );
not \U$14534 ( \14877 , \1462 );
and \U$14535 ( \14878 , \2042 , RI9870c90_103);
and \U$14536 ( \14879 , RI9871230_115, \2040 );
nor \U$14537 ( \14880 , \14878 , \14879 );
not \U$14538 ( \14881 , \14880 );
or \U$14539 ( \14882 , \14877 , \14881 );
or \U$14540 ( \14883 , \14880 , \1462 );
nand \U$14541 ( \14884 , \14882 , \14883 );
xor \U$14542 ( \14885 , \14876 , \14884 );
and \U$14543 ( \14886 , \2464 , RI9871410_119);
and \U$14544 ( \14887 , RI98716e0_125, \2462 );
nor \U$14545 ( \14888 , \14886 , \14887 );
and \U$14546 ( \14889 , \14888 , \2468 );
not \U$14547 ( \14890 , \14888 );
and \U$14548 ( \14891 , \14890 , \2263 );
nor \U$14549 ( \14892 , \14889 , \14891 );
and \U$14550 ( \14893 , \14885 , \14892 );
and \U$14551 ( \14894 , \14876 , \14884 );
or \U$14552 ( \14895 , \14893 , \14894 );
and \U$14553 ( \14896 , \14869 , \14895 );
and \U$14554 ( \14897 , \14842 , \14868 );
or \U$14555 ( \14898 , \14896 , \14897 );
and \U$14556 ( \14899 , \8486 , RI986e620_21);
and \U$14557 ( \14900 , RI986f7f0_59, \8484 );
nor \U$14558 ( \14901 , \14899 , \14900 );
and \U$14559 ( \14902 , \14901 , \8050 );
not \U$14560 ( \14903 , \14901 );
and \U$14561 ( \14904 , \14903 , \8051 );
nor \U$14562 ( \14905 , \14902 , \14904 );
and \U$14563 ( \14906 , \9237 , RI986f700_57);
and \U$14564 ( \14907 , RI986f9d0_63, \9235 );
nor \U$14565 ( \14908 , \14906 , \14907 );
and \U$14566 ( \14909 , \14908 , \9241 );
not \U$14567 ( \14910 , \14908 );
and \U$14568 ( \14911 , \14910 , \8836 );
nor \U$14569 ( \14912 , \14909 , \14911 );
xor \U$14570 ( \14913 , \14905 , \14912 );
and \U$14571 ( \14914 , \9505 , RI986f8e0_61);
and \U$14572 ( \14915 , RI986f430_51, \9503 );
nor \U$14573 ( \14916 , \14914 , \14915 );
and \U$14574 ( \14917 , \14916 , \9510 );
not \U$14575 ( \14918 , \14916 );
and \U$14576 ( \14919 , \14918 , \9513 );
nor \U$14577 ( \14920 , \14917 , \14919 );
and \U$14578 ( \14921 , \14913 , \14920 );
and \U$14579 ( \14922 , \14905 , \14912 );
or \U$14580 ( \14923 , \14921 , \14922 );
and \U$14581 ( \14924 , \13045 , RI986dcc0_1);
and \U$14582 ( \14925 , RI986e170_11, \13043 );
nor \U$14583 ( \14926 , \14924 , \14925 );
and \U$14584 ( \14927 , \14926 , \13047 );
not \U$14585 ( \14928 , \14926 );
and \U$14586 ( \14929 , \14928 , \12619 );
nor \U$14587 ( \14930 , \14927 , \14929 );
and \U$14588 ( \14931 , RI98734e0_189, RI98735d0_191);
not \U$14589 ( \14932 , RI9873558_190);
and \U$14590 ( \14933 , \14932 , RI98735d0_191);
nor \U$14591 ( \14934 , \14932 , RI98735d0_191);
or \U$14592 ( \14935 , \14933 , \14934 );
nor \U$14593 ( \14936 , RI98734e0_189, RI98735d0_191);
nor \U$14594 ( \14937 , \14931 , \14935 , \14936 );
nand \U$14595 ( \14938 , RI986e350_15, \14937 );
and \U$14596 ( \14939 , \14938 , \14539 );
not \U$14597 ( \14940 , \14938 );
and \U$14598 ( \14941 , \14940 , \14538 );
nor \U$14599 ( \14942 , \14939 , \14941 );
xor \U$14600 ( \14943 , \14930 , \14942 );
and \U$14601 ( \14944 , \13882 , RI986e080_9);
and \U$14602 ( \14945 , RI986e260_13, \13880 );
nor \U$14603 ( \14946 , \14944 , \14945 );
and \U$14604 ( \14947 , \14946 , \13358 );
not \U$14605 ( \14948 , \14946 );
and \U$14606 ( \14949 , \14948 , \13359 );
nor \U$14607 ( \14950 , \14947 , \14949 );
and \U$14608 ( \14951 , \14943 , \14950 );
and \U$14609 ( \14952 , \14930 , \14942 );
or \U$14610 ( \14953 , \14951 , \14952 );
xor \U$14611 ( \14954 , \14923 , \14953 );
and \U$14612 ( \14955 , \10424 , RI986f340_49);
and \U$14613 ( \14956 , RI986f520_53, \10422 );
nor \U$14614 ( \14957 , \14955 , \14956 );
and \U$14615 ( \14958 , \14957 , \9840 );
not \U$14616 ( \14959 , \14957 );
and \U$14617 ( \14960 , \14959 , \10428 );
nor \U$14618 ( \14961 , \14958 , \14960 );
and \U$14619 ( \14962 , \11696 , RI986f610_55);
and \U$14620 ( \14963 , RI986df90_7, \11694 );
nor \U$14621 ( \14964 , \14962 , \14963 );
and \U$14622 ( \14965 , \14964 , \10965 );
not \U$14623 ( \14966 , \14964 );
and \U$14624 ( \14967 , \14966 , \11702 );
nor \U$14625 ( \14968 , \14965 , \14967 );
xor \U$14626 ( \14969 , \14961 , \14968 );
and \U$14627 ( \14970 , \12293 , RI986dea0_5);
and \U$14628 ( \14971 , RI986ddb0_3, \12291 );
nor \U$14629 ( \14972 , \14970 , \14971 );
and \U$14630 ( \14973 , \14972 , \11687 );
not \U$14631 ( \14974 , \14972 );
and \U$14632 ( \14975 , \14974 , \11686 );
nor \U$14633 ( \14976 , \14973 , \14975 );
and \U$14634 ( \14977 , \14969 , \14976 );
and \U$14635 ( \14978 , \14961 , \14968 );
or \U$14636 ( \14979 , \14977 , \14978 );
and \U$14637 ( \14980 , \14954 , \14979 );
and \U$14638 ( \14981 , \14923 , \14953 );
or \U$14639 ( \14982 , \14980 , \14981 );
xor \U$14640 ( \14983 , \14898 , \14982 );
and \U$14641 ( \14984 , \7729 , RI986e440_17);
and \U$14642 ( \14985 , RI986e710_23, \7727 );
nor \U$14643 ( \14986 , \14984 , \14985 );
and \U$14644 ( \14987 , \14986 , \7480 );
not \U$14645 ( \14988 , \14986 );
and \U$14646 ( \14989 , \14988 , \7733 );
nor \U$14647 ( \14990 , \14987 , \14989 );
and \U$14648 ( \14991 , \6453 , RI986ef80_41);
and \U$14649 ( \14992 , RI986f250_47, \6451 );
nor \U$14650 ( \14993 , \14991 , \14992 );
and \U$14651 ( \14994 , \14993 , \6190 );
not \U$14652 ( \14995 , \14993 );
and \U$14653 ( \14996 , \14995 , \6180 );
nor \U$14654 ( \14997 , \14994 , \14996 );
xor \U$14655 ( \14998 , \14990 , \14997 );
and \U$14656 ( \14999 , \7079 , RI986f160_45);
and \U$14657 ( \15000 , RI986e530_19, \7077 );
nor \U$14658 ( \15001 , \14999 , \15000 );
and \U$14659 ( \15002 , \15001 , \6710 );
not \U$14660 ( \15003 , \15001 );
and \U$14661 ( \15004 , \15003 , \6709 );
nor \U$14662 ( \15005 , \15002 , \15004 );
and \U$14663 ( \15006 , \14998 , \15005 );
and \U$14664 ( \15007 , \14990 , \14997 );
or \U$14665 ( \15008 , \15006 , \15007 );
not \U$14666 ( \15009 , \3412 );
and \U$14667 ( \15010 , \3683 , RI98715f0_123);
and \U$14668 ( \15011 , RI986ead0_31, \3681 );
nor \U$14669 ( \15012 , \15010 , \15011 );
not \U$14670 ( \15013 , \15012 );
or \U$14671 ( \15014 , \15009 , \15013 );
or \U$14672 ( \15015 , \15012 , \3918 );
nand \U$14673 ( \15016 , \15014 , \15015 );
not \U$14674 ( \15017 , \3406 );
and \U$14675 ( \15018 , \3254 , RI98717d0_127);
and \U$14676 ( \15019 , RI9871500_121, \3252 );
nor \U$14677 ( \15020 , \15018 , \15019 );
not \U$14678 ( \15021 , \15020 );
or \U$14679 ( \15022 , \15017 , \15021 );
or \U$14680 ( \15023 , \15020 , \2935 );
nand \U$14681 ( \15024 , \15022 , \15023 );
xor \U$14682 ( \15025 , \15016 , \15024 );
and \U$14683 ( \15026 , \4203 , RI986e9e0_29);
and \U$14684 ( \15027 , RI986e8f0_27, \4201 );
nor \U$14685 ( \15028 , \15026 , \15027 );
and \U$14686 ( \15029 , \15028 , \4207 );
not \U$14687 ( \15030 , \15028 );
and \U$14688 ( \15031 , \15030 , \3922 );
nor \U$14689 ( \15032 , \15029 , \15031 );
and \U$14690 ( \15033 , \15025 , \15032 );
and \U$14691 ( \15034 , \15016 , \15024 );
or \U$14692 ( \15035 , \15033 , \15034 );
xor \U$14693 ( \15036 , \15008 , \15035 );
and \U$14694 ( \15037 , \5881 , RI986ecb0_35);
and \U$14695 ( \15038 , RI986f070_43, \5879 );
nor \U$14696 ( \15039 , \15037 , \15038 );
and \U$14697 ( \15040 , \15039 , \5594 );
not \U$14698 ( \15041 , \15039 );
and \U$14699 ( \15042 , \15041 , \5885 );
nor \U$14700 ( \15043 , \15040 , \15042 );
not \U$14701 ( \15044 , \4521 );
and \U$14702 ( \15045 , \4710 , RI986e800_25);
and \U$14703 ( \15046 , RI986ee90_39, \4708 );
nor \U$14704 ( \15047 , \15045 , \15046 );
not \U$14705 ( \15048 , \15047 );
or \U$14706 ( \15049 , \15044 , \15048 );
or \U$14707 ( \15050 , \15047 , \4521 );
nand \U$14708 ( \15051 , \15049 , \15050 );
xor \U$14709 ( \15052 , \15043 , \15051 );
and \U$14710 ( \15053 , \5318 , RI986eda0_37);
and \U$14711 ( \15054 , RI986ebc0_33, \5316 );
nor \U$14712 ( \15055 , \15053 , \15054 );
and \U$14713 ( \15056 , \15055 , \5052 );
not \U$14714 ( \15057 , \15055 );
and \U$14715 ( \15058 , \15057 , \5322 );
nor \U$14716 ( \15059 , \15056 , \15058 );
and \U$14717 ( \15060 , \15052 , \15059 );
and \U$14718 ( \15061 , \15043 , \15051 );
or \U$14719 ( \15062 , \15060 , \15061 );
and \U$14720 ( \15063 , \15036 , \15062 );
and \U$14721 ( \15064 , \15008 , \15035 );
or \U$14722 ( \15065 , \15063 , \15064 );
and \U$14723 ( \15066 , \14983 , \15065 );
and \U$14724 ( \15067 , \14898 , \14982 );
or \U$14725 ( \15068 , \15066 , \15067 );
xor \U$14726 ( \15069 , \14816 , \15068 );
xor \U$14727 ( \15070 , \14399 , \14407 );
xor \U$14728 ( \15071 , \15070 , \14415 );
xor \U$14729 ( \15072 , \14346 , \14353 );
xor \U$14730 ( \15073 , \15072 , \14361 );
and \U$14731 ( \15074 , \15071 , \15073 );
xor \U$14732 ( \15075 , \14511 , \14518 );
xor \U$14733 ( \15076 , \15075 , \14526 );
xor \U$14734 ( \15077 , \14346 , \14353 );
xor \U$14735 ( \15078 , \15077 , \14361 );
and \U$14736 ( \15079 , \15076 , \15078 );
and \U$14737 ( \15080 , \15071 , \15076 );
or \U$14738 ( \15081 , \15074 , \15079 , \15080 );
xor \U$14739 ( \15082 , \14558 , \14565 );
xor \U$14740 ( \15083 , \15082 , \14573 );
xor \U$14741 ( \15084 , \14536 , \14539 );
xor \U$14742 ( \15085 , \15084 , \14547 );
and \U$14743 ( \15086 , \15083 , \15085 );
xor \U$14744 ( \15087 , \15081 , \15086 );
xor \U$14745 ( \15088 , \13875 , \13887 );
xor \U$14746 ( \15089 , \15088 , \13895 );
xor \U$14747 ( \15090 , \14600 , \14605 );
xor \U$14748 ( \15091 , \15089 , \15090 );
and \U$14749 ( \15092 , \15087 , \15091 );
and \U$14750 ( \15093 , \15081 , \15086 );
or \U$14751 ( \15094 , \15092 , \15093 );
and \U$14752 ( \15095 , \15069 , \15094 );
and \U$14753 ( \15096 , \14816 , \15068 );
or \U$14754 ( \15097 , \15095 , \15096 );
and \U$14755 ( \15098 , \14742 , \15097 );
not \U$14756 ( \15099 , \14742 );
not \U$14757 ( \15100 , \15097 );
and \U$14758 ( \15101 , \15099 , \15100 );
xor \U$14759 ( \15102 , \14291 , \14325 );
xor \U$14760 ( \15103 , \15102 , \14336 );
not \U$14761 ( \15104 , \14594 );
not \U$14762 ( \15105 , \14610 );
or \U$14763 ( \15106 , \15104 , \15105 );
or \U$14764 ( \15107 , \14610 , \14594 );
nand \U$14765 ( \15108 , \15106 , \15107 );
not \U$14766 ( \15109 , \15108 );
not \U$14767 ( \15110 , \14585 );
and \U$14768 ( \15111 , \15109 , \15110 );
and \U$14769 ( \15112 , \15108 , \14585 );
nor \U$14770 ( \15113 , \15111 , \15112 );
not \U$14771 ( \15114 , \15113 );
and \U$14772 ( \15115 , \15103 , \15114 );
not \U$14773 ( \15116 , \15103 );
not \U$14774 ( \15117 , \15114 );
and \U$14775 ( \15118 , \15116 , \15117 );
xor \U$14776 ( \15119 , \14252 , \14262 );
xor \U$14777 ( \15120 , \15119 , \14273 );
nor \U$14778 ( \15121 , \15118 , \15120 );
nor \U$14779 ( \15122 , \15115 , \15121 );
nor \U$14780 ( \15123 , \15101 , \15122 );
nor \U$14781 ( \15124 , \15098 , \15123 );
nor \U$14782 ( \15125 , \14708 , \15124 );
nor \U$14783 ( \15126 , \14707 , \15125 );
not \U$14784 ( \15127 , \15126 );
nand \U$14785 ( \15128 , \14686 , \15127 );
nand \U$14786 ( \15129 , \14685 , \15128 );
xor \U$14787 ( \15130 , \14180 , \14192 );
xor \U$14788 ( \15131 , \15130 , \14197 );
xor \U$14789 ( \15132 , \15129 , \15131 );
xor \U$14790 ( \15133 , \14214 , \14226 );
xor \U$14791 ( \15134 , \15133 , \14663 );
and \U$14792 ( \15135 , \15132 , \15134 );
and \U$14793 ( \15136 , \15129 , \15131 );
or \U$14794 ( \15137 , \15135 , \15136 );
not \U$14795 ( \15138 , \14666 );
not \U$14796 ( \15139 , \14669 );
or \U$14797 ( \15140 , \15138 , \15139 );
or \U$14798 ( \15141 , \14669 , \14666 );
nand \U$14799 ( \15142 , \15140 , \15141 );
and \U$14800 ( \15143 , \15137 , \15142 );
xor \U$14801 ( \15144 , \15142 , \15137 );
xor \U$14802 ( \15145 , \15129 , \15131 );
xor \U$14803 ( \15146 , \15145 , \15134 );
not \U$14804 ( \15147 , \15146 );
not \U$14805 ( \15148 , \14683 );
not \U$14806 ( \15149 , \15126 );
and \U$14807 ( \15150 , \15148 , \15149 );
and \U$14808 ( \15151 , \14683 , \15126 );
nor \U$14809 ( \15152 , \15150 , \15151 );
not \U$14810 ( \15153 , \15152 );
not \U$14811 ( \15154 , \14680 );
and \U$14812 ( \15155 , \15153 , \15154 );
and \U$14813 ( \15156 , \15152 , \14680 );
nor \U$14814 ( \15157 , \15155 , \15156 );
not \U$14815 ( \15158 , \15157 );
xor \U$14816 ( \15159 , \14754 , \14802 );
xor \U$14817 ( \15160 , \15159 , \14813 );
xor \U$14818 ( \15161 , \15081 , \15086 );
xor \U$14819 ( \15162 , \15161 , \15091 );
and \U$14820 ( \15163 , \15160 , \15162 );
xor \U$14821 ( \15164 , \14328 , \14330 );
xor \U$14822 ( \15165 , \15164 , \14333 );
xor \U$14823 ( \15166 , \14710 , \14717 );
xor \U$14824 ( \15167 , \15165 , \15166 );
xor \U$14825 ( \15168 , \15081 , \15086 );
xor \U$14826 ( \15169 , \15168 , \15091 );
and \U$14827 ( \15170 , \15167 , \15169 );
and \U$14828 ( \15171 , \15160 , \15167 );
or \U$14829 ( \15172 , \15163 , \15170 , \15171 );
xor \U$14830 ( \15173 , \14849 , \14856 );
xor \U$14831 ( \15174 , \15173 , \14865 );
xor \U$14832 ( \15175 , \14779 , \14787 );
xor \U$14833 ( \15176 , \15175 , \14796 );
xor \U$14834 ( \15177 , \15174 , \15176 );
xor \U$14835 ( \15178 , \14823 , \14831 );
xor \U$14836 ( \15179 , \15178 , \14839 );
and \U$14837 ( \15180 , \15177 , \15179 );
and \U$14838 ( \15181 , \15174 , \15176 );
or \U$14839 ( \15182 , \15180 , \15181 );
not \U$14840 ( \15183 , \345 );
and \U$14841 ( \15184 , \354 , RI98706f0_91);
and \U$14842 ( \15185 , RI9870600_89, \352 );
nor \U$14843 ( \15186 , \15184 , \15185 );
not \U$14844 ( \15187 , \15186 );
or \U$14845 ( \15188 , \15183 , \15187 );
or \U$14846 ( \15189 , \15186 , \361 );
nand \U$14847 ( \15190 , \15188 , \15189 );
not \U$14848 ( \15191 , RI9870510_87);
nor \U$14849 ( \15192 , \15191 , \407 );
xor \U$14850 ( \15193 , \15190 , \15192 );
and \U$14851 ( \15194 , \416 , RI9870330_83);
and \U$14852 ( \15195 , RI9870240_81, \414 );
nor \U$14853 ( \15196 , \15194 , \15195 );
and \U$14854 ( \15197 , \15196 , \422 );
not \U$14855 ( \15198 , \15196 );
and \U$14856 ( \15199 , \15198 , \421 );
nor \U$14857 ( \15200 , \15197 , \15199 );
and \U$14858 ( \15201 , \15193 , \15200 );
and \U$14859 ( \15202 , \15190 , \15192 );
or \U$14860 ( \15203 , \15201 , \15202 );
or \U$14861 ( \15204 , \14762 , \14755 );
nand \U$14862 ( \15205 , \15204 , \14763 );
xor \U$14863 ( \15206 , \15203 , \15205 );
not \U$14864 ( \15207 , \386 );
and \U$14865 ( \15208 , \395 , RI98708d0_95);
and \U$14866 ( \15209 , RI98707e0_93, \393 );
nor \U$14867 ( \15210 , \15208 , \15209 );
not \U$14868 ( \15211 , \15210 );
or \U$14869 ( \15212 , \15207 , \15211 );
or \U$14870 ( \15213 , \15210 , \487 );
nand \U$14871 ( \15214 , \15212 , \15213 );
not \U$14872 ( \15215 , \456 );
and \U$14873 ( \15216 , \465 , RI986fd90_71);
and \U$14874 ( \15217 , RI986fca0_69, \463 );
nor \U$14875 ( \15218 , \15216 , \15217 );
not \U$14876 ( \15219 , \15218 );
or \U$14877 ( \15220 , \15215 , \15219 );
or \U$14878 ( \15221 , \15218 , \456 );
nand \U$14879 ( \15222 , \15220 , \15221 );
xor \U$14880 ( \15223 , \15214 , \15222 );
not \U$14881 ( \15224 , \365 );
and \U$14882 ( \15225 , \376 , RI986fac0_65);
and \U$14883 ( \15226 , RI986fbb0_67, \374 );
nor \U$14884 ( \15227 , \15225 , \15226 );
not \U$14885 ( \15228 , \15227 );
or \U$14886 ( \15229 , \15224 , \15228 );
or \U$14887 ( \15230 , \15227 , \367 );
nand \U$14888 ( \15231 , \15229 , \15230 );
and \U$14889 ( \15232 , \15223 , \15231 );
and \U$14890 ( \15233 , \15214 , \15222 );
or \U$14891 ( \15234 , \15232 , \15233 );
and \U$14892 ( \15235 , \15206 , \15234 );
and \U$14893 ( \15236 , \15203 , \15205 );
or \U$14894 ( \15237 , \15235 , \15236 );
xor \U$14895 ( \15238 , \15182 , \15237 );
xor \U$14896 ( \15239 , \15016 , \15024 );
xor \U$14897 ( \15240 , \15239 , \15032 );
xor \U$14898 ( \15241 , \14876 , \14884 );
xor \U$14899 ( \15242 , \15241 , \14892 );
and \U$14900 ( \15243 , \15240 , \15242 );
xor \U$14901 ( \15244 , \15043 , \15051 );
xor \U$14902 ( \15245 , \15244 , \15059 );
xor \U$14903 ( \15246 , \14876 , \14884 );
xor \U$14904 ( \15247 , \15246 , \14892 );
and \U$14905 ( \15248 , \15245 , \15247 );
and \U$14906 ( \15249 , \15240 , \15245 );
or \U$14907 ( \15250 , \15243 , \15248 , \15249 );
and \U$14908 ( \15251 , \15238 , \15250 );
and \U$14909 ( \15252 , \15182 , \15237 );
or \U$14910 ( \15253 , \15251 , \15252 );
and \U$14911 ( \15254 , \5318 , RI986ee90_39);
and \U$14912 ( \15255 , RI986eda0_37, \5316 );
nor \U$14913 ( \15256 , \15254 , \15255 );
and \U$14914 ( \15257 , \15256 , \5322 );
not \U$14915 ( \15258 , \15256 );
and \U$14916 ( \15259 , \15258 , \5052 );
nor \U$14917 ( \15260 , \15257 , \15259 );
and \U$14918 ( \15261 , \5881 , RI986ebc0_33);
and \U$14919 ( \15262 , RI986ecb0_35, \5879 );
nor \U$14920 ( \15263 , \15261 , \15262 );
and \U$14921 ( \15264 , \15263 , \5885 );
not \U$14922 ( \15265 , \15263 );
and \U$14923 ( \15266 , \15265 , \5594 );
nor \U$14924 ( \15267 , \15264 , \15266 );
or \U$14925 ( \15268 , \15260 , \15267 );
not \U$14926 ( \15269 , \15267 );
not \U$14927 ( \15270 , \15260 );
or \U$14928 ( \15271 , \15269 , \15270 );
and \U$14929 ( \15272 , \6453 , RI986f070_43);
and \U$14930 ( \15273 , RI986ef80_41, \6451 );
nor \U$14931 ( \15274 , \15272 , \15273 );
and \U$14932 ( \15275 , \15274 , \6190 );
not \U$14933 ( \15276 , \15274 );
and \U$14934 ( \15277 , \15276 , \6705 );
nor \U$14935 ( \15278 , \15275 , \15277 );
nand \U$14936 ( \15279 , \15271 , \15278 );
nand \U$14937 ( \15280 , \15268 , \15279 );
and \U$14938 ( \15281 , \3683 , RI9871500_121);
and \U$14939 ( \15282 , RI98715f0_123, \3681 );
nor \U$14940 ( \15283 , \15281 , \15282 );
not \U$14941 ( \15284 , \15283 );
not \U$14942 ( \15285 , \3412 );
and \U$14943 ( \15286 , \15284 , \15285 );
and \U$14944 ( \15287 , \15283 , \3918 );
nor \U$14945 ( \15288 , \15286 , \15287 );
and \U$14946 ( \15289 , \4203 , RI986ead0_31);
and \U$14947 ( \15290 , RI986e9e0_29, \4201 );
nor \U$14948 ( \15291 , \15289 , \15290 );
and \U$14949 ( \15292 , \15291 , \3923 );
not \U$14950 ( \15293 , \15291 );
and \U$14951 ( \15294 , \15293 , \4207 );
nor \U$14952 ( \15295 , \15292 , \15294 );
or \U$14953 ( \15296 , \15288 , \15295 );
not \U$14954 ( \15297 , \15295 );
not \U$14955 ( \15298 , \15288 );
or \U$14956 ( \15299 , \15297 , \15298 );
not \U$14957 ( \15300 , \4519 );
and \U$14958 ( \15301 , \4710 , RI986e8f0_27);
and \U$14959 ( \15302 , RI986e800_25, \4708 );
nor \U$14960 ( \15303 , \15301 , \15302 );
not \U$14961 ( \15304 , \15303 );
or \U$14962 ( \15305 , \15300 , \15304 );
or \U$14963 ( \15306 , \15303 , \4521 );
nand \U$14964 ( \15307 , \15305 , \15306 );
nand \U$14965 ( \15308 , \15299 , \15307 );
nand \U$14966 ( \15309 , \15296 , \15308 );
xor \U$14967 ( \15310 , \15280 , \15309 );
and \U$14968 ( \15311 , \7079 , RI986f250_47);
and \U$14969 ( \15312 , RI986f160_45, \7077 );
nor \U$14970 ( \15313 , \15311 , \15312 );
and \U$14971 ( \15314 , \15313 , \6709 );
not \U$14972 ( \15315 , \15313 );
and \U$14973 ( \15316 , \15315 , \6710 );
nor \U$14974 ( \15317 , \15314 , \15316 );
and \U$14975 ( \15318 , \7729 , RI986e530_19);
and \U$14976 ( \15319 , RI986e440_17, \7727 );
nor \U$14977 ( \15320 , \15318 , \15319 );
and \U$14978 ( \15321 , \15320 , \7733 );
not \U$14979 ( \15322 , \15320 );
and \U$14980 ( \15323 , \15322 , \7480 );
nor \U$14981 ( \15324 , \15321 , \15323 );
or \U$14982 ( \15325 , \15317 , \15324 );
not \U$14983 ( \15326 , \15324 );
not \U$14984 ( \15327 , \15317 );
or \U$14985 ( \15328 , \15326 , \15327 );
and \U$14986 ( \15329 , \8486 , RI986e710_23);
and \U$14987 ( \15330 , RI986e620_21, \8484 );
nor \U$14988 ( \15331 , \15329 , \15330 );
and \U$14989 ( \15332 , \15331 , \8050 );
not \U$14990 ( \15333 , \15331 );
and \U$14991 ( \15334 , \15333 , \8051 );
nor \U$14992 ( \15335 , \15332 , \15334 );
nand \U$14993 ( \15336 , \15328 , \15335 );
nand \U$14994 ( \15337 , \15325 , \15336 );
and \U$14995 ( \15338 , \15310 , \15337 );
and \U$14996 ( \15339 , \15280 , \15309 );
or \U$14997 ( \15340 , \15338 , \15339 );
and \U$14998 ( \15341 , \14937 , RI986e260_13);
and \U$14999 ( \15342 , RI986e350_15, \14935 );
nor \U$15000 ( \15343 , \15341 , \15342 );
and \U$15001 ( \15344 , \15343 , \14538 );
not \U$15002 ( \15345 , \15343 );
and \U$15003 ( \15346 , \15345 , \14539 );
nor \U$15004 ( \15347 , \15344 , \15346 );
xor \U$15005 ( \15348 , \15347 , RI9873558_190);
and \U$15006 ( \15349 , \13882 , RI986e170_11);
and \U$15007 ( \15350 , RI986e080_9, \13880 );
nor \U$15008 ( \15351 , \15349 , \15350 );
and \U$15009 ( \15352 , \15351 , \13359 );
not \U$15010 ( \15353 , \15351 );
and \U$15011 ( \15354 , \15353 , \13358 );
nor \U$15012 ( \15355 , \15352 , \15354 );
and \U$15013 ( \15356 , \15348 , \15355 );
and \U$15014 ( \15357 , \15347 , RI9873558_190);
or \U$15015 ( \15358 , \15356 , \15357 );
and \U$15016 ( \15359 , \11696 , RI986f520_53);
and \U$15017 ( \15360 , RI986f610_55, \11694 );
nor \U$15018 ( \15361 , \15359 , \15360 );
and \U$15019 ( \15362 , \15361 , \11702 );
not \U$15020 ( \15363 , \15361 );
and \U$15021 ( \15364 , \15363 , \10965 );
nor \U$15022 ( \15365 , \15362 , \15364 );
not \U$15023 ( \15366 , \15365 );
and \U$15024 ( \15367 , \12293 , RI986df90_7);
and \U$15025 ( \15368 , RI986dea0_5, \12291 );
nor \U$15026 ( \15369 , \15367 , \15368 );
and \U$15027 ( \15370 , \15369 , \11686 );
not \U$15028 ( \15371 , \15369 );
and \U$15029 ( \15372 , \15371 , \11687 );
nor \U$15030 ( \15373 , \15370 , \15372 );
not \U$15031 ( \15374 , \15373 );
and \U$15032 ( \15375 , \15366 , \15374 );
and \U$15033 ( \15376 , \15373 , \15365 );
and \U$15034 ( \15377 , \13045 , RI986ddb0_3);
and \U$15035 ( \15378 , RI986dcc0_1, \13043 );
nor \U$15036 ( \15379 , \15377 , \15378 );
and \U$15037 ( \15380 , \15379 , \12619 );
not \U$15038 ( \15381 , \15379 );
and \U$15039 ( \15382 , \15381 , \13047 );
nor \U$15040 ( \15383 , \15380 , \15382 );
nor \U$15041 ( \15384 , \15376 , \15383 );
nor \U$15042 ( \15385 , \15375 , \15384 );
xor \U$15043 ( \15386 , \15358 , \15385 );
and \U$15044 ( \15387 , \9237 , RI986f7f0_59);
and \U$15045 ( \15388 , RI986f700_57, \9235 );
nor \U$15046 ( \15389 , \15387 , \15388 );
and \U$15047 ( \15390 , \15389 , \8836 );
not \U$15048 ( \15391 , \15389 );
and \U$15049 ( \15392 , \15391 , \9241 );
nor \U$15050 ( \15393 , \15390 , \15392 );
and \U$15051 ( \15394 , \9505 , RI986f9d0_63);
and \U$15052 ( \15395 , RI986f8e0_61, \9503 );
nor \U$15053 ( \15396 , \15394 , \15395 );
and \U$15054 ( \15397 , \15396 , \9513 );
not \U$15055 ( \15398 , \15396 );
and \U$15056 ( \15399 , \15398 , \9510 );
nor \U$15057 ( \15400 , \15397 , \15399 );
xor \U$15058 ( \15401 , \15393 , \15400 );
and \U$15059 ( \15402 , \10424 , RI986f430_51);
and \U$15060 ( \15403 , RI986f340_49, \10422 );
nor \U$15061 ( \15404 , \15402 , \15403 );
and \U$15062 ( \15405 , \15404 , \10428 );
not \U$15063 ( \15406 , \15404 );
and \U$15064 ( \15407 , \15406 , \9840 );
nor \U$15065 ( \15408 , \15405 , \15407 );
and \U$15066 ( \15409 , \15401 , \15408 );
and \U$15067 ( \15410 , \15393 , \15400 );
or \U$15068 ( \15411 , \15409 , \15410 );
and \U$15069 ( \15412 , \15386 , \15411 );
and \U$15070 ( \15413 , \15358 , \15385 );
nor \U$15071 ( \15414 , \15412 , \15413 );
xor \U$15072 ( \15415 , \15340 , \15414 );
and \U$15073 ( \15416 , \2274 , RI9871230_115);
and \U$15074 ( \15417 , RI9871140_113, \2272 );
nor \U$15075 ( \15418 , \15416 , \15417 );
and \U$15076 ( \15419 , \15418 , \2031 );
not \U$15077 ( \15420 , \15418 );
and \U$15078 ( \15421 , \15420 , \2030 );
nor \U$15079 ( \15422 , \15419 , \15421 );
and \U$15080 ( \15423 , \3254 , RI98716e0_125);
and \U$15081 ( \15424 , RI98717d0_127, \3252 );
nor \U$15082 ( \15425 , \15423 , \15424 );
not \U$15083 ( \15426 , \15425 );
not \U$15084 ( \15427 , \2935 );
and \U$15085 ( \15428 , \15426 , \15427 );
and \U$15086 ( \15429 , \15425 , \3406 );
nor \U$15087 ( \15430 , \15428 , \15429 );
or \U$15088 ( \15431 , \15422 , \15430 );
not \U$15089 ( \15432 , \15430 );
not \U$15090 ( \15433 , \15422 );
or \U$15091 ( \15434 , \15432 , \15433 );
and \U$15092 ( \15435 , \2464 , RI9871320_117);
and \U$15093 ( \15436 , RI9871410_119, \2462 );
nor \U$15094 ( \15437 , \15435 , \15436 );
and \U$15095 ( \15438 , \15437 , \2468 );
not \U$15096 ( \15439 , \15437 );
and \U$15097 ( \15440 , \15439 , \2263 );
nor \U$15098 ( \15441 , \15438 , \15440 );
nand \U$15099 ( \15442 , \15434 , \15441 );
nand \U$15100 ( \15443 , \15431 , \15442 );
and \U$15101 ( \15444 , \776 , RI9870060_77);
and \U$15102 ( \15445 , RI9870150_79, \774 );
nor \U$15103 ( \15446 , \15444 , \15445 );
and \U$15104 ( \15447 , \15446 , \474 );
not \U$15105 ( \15448 , \15446 );
and \U$15106 ( \15449 , \15448 , \451 );
nor \U$15107 ( \15450 , \15447 , \15449 );
and \U$15108 ( \15451 , \438 , RI986ff70_75);
and \U$15109 ( \15452 , RI986fe80_73, \436 );
nor \U$15110 ( \15453 , \15451 , \15452 );
and \U$15111 ( \15454 , \15453 , \444 );
not \U$15112 ( \15455 , \15453 );
and \U$15113 ( \15456 , \15455 , \443 );
nor \U$15114 ( \15457 , \15454 , \15456 );
xor \U$15115 ( \15458 , \15450 , \15457 );
not \U$15116 ( \15459 , \1128 );
and \U$15117 ( \15460 , \1293 , RI9870f60_109);
and \U$15118 ( \15461 , RI9870ab0_99, \1291 );
nor \U$15119 ( \15462 , \15460 , \15461 );
not \U$15120 ( \15463 , \15462 );
or \U$15121 ( \15464 , \15459 , \15463 );
or \U$15122 ( \15465 , \15462 , \1128 );
nand \U$15123 ( \15466 , \15464 , \15465 );
and \U$15124 ( \15467 , \15458 , \15466 );
and \U$15125 ( \15468 , \15450 , \15457 );
or \U$15126 ( \15469 , \15467 , \15468 );
xor \U$15127 ( \15470 , \15443 , \15469 );
and \U$15128 ( \15471 , \1329 , RI9870d80_105);
and \U$15129 ( \15472 , RI98709c0_97, \1327 );
nor \U$15130 ( \15473 , \15471 , \15472 );
and \U$15131 ( \15474 , \15473 , \1337 );
not \U$15132 ( \15475 , \15473 );
and \U$15133 ( \15476 , \15475 , \1336 );
nor \U$15134 ( \15477 , \15474 , \15476 );
and \U$15135 ( \15478 , \1311 , RI9870e70_107);
and \U$15136 ( \15479 , RI9870ba0_101, \1309 );
nor \U$15137 ( \15480 , \15478 , \15479 );
and \U$15138 ( \15481 , \15480 , \1315 );
not \U$15139 ( \15482 , \15480 );
and \U$15140 ( \15483 , \15482 , \1458 );
nor \U$15141 ( \15484 , \15481 , \15483 );
or \U$15142 ( \15485 , \15477 , \15484 );
not \U$15143 ( \15486 , \15484 );
not \U$15144 ( \15487 , \15477 );
or \U$15145 ( \15488 , \15486 , \15487 );
not \U$15146 ( \15489 , \1462 );
and \U$15147 ( \15490 , \2042 , RI9871050_111);
and \U$15148 ( \15491 , RI9870c90_103, \2040 );
nor \U$15149 ( \15492 , \15490 , \15491 );
not \U$15150 ( \15493 , \15492 );
or \U$15151 ( \15494 , \15489 , \15493 );
or \U$15152 ( \15495 , \15492 , \2034 );
nand \U$15153 ( \15496 , \15494 , \15495 );
nand \U$15154 ( \15497 , \15488 , \15496 );
nand \U$15155 ( \15498 , \15485 , \15497 );
and \U$15156 ( \15499 , \15470 , \15498 );
and \U$15157 ( \15500 , \15443 , \15469 );
or \U$15158 ( \15501 , \15499 , \15500 );
and \U$15159 ( \15502 , \15415 , \15501 );
and \U$15160 ( \15503 , \15340 , \15414 );
or \U$15161 ( \15504 , \15502 , \15503 );
xor \U$15162 ( \15505 , \15253 , \15504 );
xor \U$15163 ( \15506 , \14905 , \14912 );
xor \U$15164 ( \15507 , \15506 , \14920 );
xor \U$15165 ( \15508 , \14990 , \14997 );
xor \U$15166 ( \15509 , \15508 , \15005 );
and \U$15167 ( \15510 , \15507 , \15509 );
xor \U$15168 ( \15511 , \14961 , \14968 );
xor \U$15169 ( \15512 , \15511 , \14976 );
xor \U$15170 ( \15513 , \14990 , \14997 );
xor \U$15171 ( \15514 , \15513 , \15005 );
and \U$15172 ( \15515 , \15512 , \15514 );
and \U$15173 ( \15516 , \15507 , \15512 );
or \U$15174 ( \15517 , \15510 , \15515 , \15516 );
xor \U$15175 ( \15518 , \15083 , \15085 );
xor \U$15176 ( \15519 , \15517 , \15518 );
xor \U$15177 ( \15520 , \14346 , \14353 );
xor \U$15178 ( \15521 , \15520 , \14361 );
xor \U$15179 ( \15522 , \15071 , \15076 );
xor \U$15180 ( \15523 , \15521 , \15522 );
and \U$15181 ( \15524 , \15519 , \15523 );
and \U$15182 ( \15525 , \15517 , \15518 );
or \U$15183 ( \15526 , \15524 , \15525 );
and \U$15184 ( \15527 , \15505 , \15526 );
and \U$15185 ( \15528 , \15253 , \15504 );
or \U$15186 ( \15529 , \15527 , \15528 );
xor \U$15187 ( \15530 , \15172 , \15529 );
xor \U$15188 ( \15531 , \14763 , \14770 );
xor \U$15189 ( \15532 , \15531 , \14799 );
xor \U$15190 ( \15533 , \14805 , \14807 );
xor \U$15191 ( \15534 , \15533 , \14810 );
and \U$15192 ( \15535 , \15532 , \15534 );
xor \U$15193 ( \15536 , \14299 , \14307 );
xor \U$15194 ( \15537 , \15536 , \14316 );
xor \U$15195 ( \15538 , \14744 , \14749 );
xor \U$15196 ( \15539 , \15537 , \15538 );
xor \U$15197 ( \15540 , \14805 , \14807 );
xor \U$15198 ( \15541 , \15540 , \14810 );
and \U$15199 ( \15542 , \15539 , \15541 );
and \U$15200 ( \15543 , \15532 , \15539 );
or \U$15201 ( \15544 , \15535 , \15542 , \15543 );
xor \U$15202 ( \15545 , \14923 , \14953 );
xor \U$15203 ( \15546 , \15545 , \14979 );
xor \U$15204 ( \15547 , \14842 , \14868 );
xor \U$15205 ( \15548 , \15547 , \14895 );
and \U$15206 ( \15549 , \15546 , \15548 );
xor \U$15207 ( \15550 , \15008 , \15035 );
xor \U$15208 ( \15551 , \15550 , \15062 );
xor \U$15209 ( \15552 , \14842 , \14868 );
xor \U$15210 ( \15553 , \15552 , \14895 );
and \U$15211 ( \15554 , \15551 , \15553 );
and \U$15212 ( \15555 , \15546 , \15551 );
or \U$15213 ( \15556 , \15549 , \15554 , \15555 );
xor \U$15214 ( \15557 , \15544 , \15556 );
xor \U$15215 ( \15558 , \14529 , \14550 );
xor \U$15216 ( \15559 , \15558 , \14576 );
xor \U$15217 ( \15560 , \14724 , \14729 );
xor \U$15218 ( \15561 , \15559 , \15560 );
and \U$15219 ( \15562 , \15557 , \15561 );
and \U$15220 ( \15563 , \15544 , \15556 );
or \U$15221 ( \15564 , \15562 , \15563 );
and \U$15222 ( \15565 , \15530 , \15564 );
and \U$15223 ( \15566 , \15172 , \15529 );
or \U$15224 ( \15567 , \15565 , \15566 );
xor \U$15225 ( \15568 , \14239 , \14241 );
xor \U$15226 ( \15569 , \15568 , \14276 );
xor \U$15227 ( \15570 , \15567 , \15569 );
xor \U$15228 ( \15571 , \14421 , \14503 );
xor \U$15229 ( \15572 , \15571 , \14579 );
xor \U$15230 ( \15573 , \14722 , \14734 );
xor \U$15231 ( \15574 , \15573 , \14739 );
and \U$15232 ( \15575 , \15572 , \15574 );
not \U$15233 ( \15576 , \15113 );
not \U$15234 ( \15577 , \15103 );
not \U$15235 ( \15578 , \15120 );
or \U$15236 ( \15579 , \15577 , \15578 );
or \U$15237 ( \15580 , \15120 , \15103 );
nand \U$15238 ( \15581 , \15579 , \15580 );
not \U$15239 ( \15582 , \15581 );
or \U$15240 ( \15583 , \15576 , \15582 );
or \U$15241 ( \15584 , \15581 , \15113 );
nand \U$15242 ( \15585 , \15583 , \15584 );
xor \U$15243 ( \15586 , \14722 , \14734 );
xor \U$15244 ( \15587 , \15586 , \14739 );
and \U$15245 ( \15588 , \15585 , \15587 );
and \U$15246 ( \15589 , \15572 , \15585 );
or \U$15247 ( \15590 , \15575 , \15588 , \15589 );
and \U$15248 ( \15591 , \15570 , \15590 );
and \U$15249 ( \15592 , \15567 , \15569 );
or \U$15250 ( \15593 , \15591 , \15592 );
xor \U$15251 ( \15594 , \14279 , \14615 );
xor \U$15252 ( \15595 , \15594 , \14632 );
xor \U$15253 ( \15596 , \15593 , \15595 );
xor \U$15254 ( \15597 , \14695 , \14697 );
xor \U$15255 ( \15598 , \15597 , \14702 );
xor \U$15256 ( \15599 , \14339 , \14582 );
xor \U$15257 ( \15600 , \15599 , \14612 );
xor \U$15258 ( \15601 , \15598 , \15600 );
not \U$15259 ( \15602 , \15122 );
xor \U$15260 ( \15603 , \15097 , \14742 );
not \U$15261 ( \15604 , \15603 );
or \U$15262 ( \15605 , \15602 , \15604 );
or \U$15263 ( \15606 , \15603 , \15122 );
nand \U$15264 ( \15607 , \15605 , \15606 );
and \U$15265 ( \15608 , \15601 , \15607 );
and \U$15266 ( \15609 , \15598 , \15600 );
or \U$15267 ( \15610 , \15608 , \15609 );
and \U$15268 ( \15611 , \15596 , \15610 );
and \U$15269 ( \15612 , \15593 , \15595 );
or \U$15270 ( \15613 , \15611 , \15612 );
nand \U$15271 ( \15614 , \15158 , \15613 );
or \U$15272 ( \15615 , \15147 , \15614 );
not \U$15273 ( \15616 , \15146 );
not \U$15274 ( \15617 , \15614 );
and \U$15275 ( \15618 , \15616 , \15617 );
and \U$15276 ( \15619 , \15146 , \15614 );
nor \U$15277 ( \15620 , \15618 , \15619 );
xor \U$15278 ( \15621 , \15172 , \15529 );
xor \U$15279 ( \15622 , \15621 , \15564 );
xor \U$15280 ( \15623 , \14876 , \14884 );
xor \U$15281 ( \15624 , \15623 , \14892 );
xor \U$15282 ( \15625 , \15240 , \15245 );
xor \U$15283 ( \15626 , \15624 , \15625 );
xor \U$15284 ( \15627 , \15174 , \15176 );
xor \U$15285 ( \15628 , \15627 , \15179 );
and \U$15286 ( \15629 , \15626 , \15628 );
xor \U$15287 ( \15630 , \14990 , \14997 );
xor \U$15288 ( \15631 , \15630 , \15005 );
xor \U$15289 ( \15632 , \15507 , \15512 );
xor \U$15290 ( \15633 , \15631 , \15632 );
xor \U$15291 ( \15634 , \15174 , \15176 );
xor \U$15292 ( \15635 , \15634 , \15179 );
and \U$15293 ( \15636 , \15633 , \15635 );
and \U$15294 ( \15637 , \15626 , \15633 );
or \U$15295 ( \15638 , \15629 , \15636 , \15637 );
xor \U$15296 ( \15639 , \15203 , \15205 );
xor \U$15297 ( \15640 , \15639 , \15234 );
xor \U$15298 ( \15641 , \15280 , \15309 );
xor \U$15299 ( \15642 , \15641 , \15337 );
xor \U$15300 ( \15643 , \15640 , \15642 );
xor \U$15301 ( \15644 , \15443 , \15469 );
xor \U$15302 ( \15645 , \15644 , \15498 );
and \U$15303 ( \15646 , \15643 , \15645 );
and \U$15304 ( \15647 , \15640 , \15642 );
or \U$15305 ( \15648 , \15646 , \15647 );
xor \U$15306 ( \15649 , \15638 , \15648 );
xor \U$15307 ( \15650 , \14842 , \14868 );
xor \U$15308 ( \15651 , \15650 , \14895 );
xor \U$15309 ( \15652 , \15546 , \15551 );
xor \U$15310 ( \15653 , \15651 , \15652 );
and \U$15311 ( \15654 , \15649 , \15653 );
and \U$15312 ( \15655 , \15638 , \15648 );
or \U$15313 ( \15656 , \15654 , \15655 );
and \U$15314 ( \15657 , \1311 , RI98709c0_97);
and \U$15315 ( \15658 , RI9870e70_107, \1309 );
nor \U$15316 ( \15659 , \15657 , \15658 );
and \U$15317 ( \15660 , \15659 , \1318 );
not \U$15318 ( \15661 , \15659 );
and \U$15319 ( \15662 , \15661 , \1458 );
nor \U$15320 ( \15663 , \15660 , \15662 );
and \U$15321 ( \15664 , \2042 , RI9870ba0_101);
and \U$15322 ( \15665 , RI9871050_111, \2040 );
nor \U$15323 ( \15666 , \15664 , \15665 );
not \U$15324 ( \15667 , \15666 );
not \U$15325 ( \15668 , \1462 );
and \U$15326 ( \15669 , \15667 , \15668 );
and \U$15327 ( \15670 , \15666 , \1462 );
nor \U$15328 ( \15671 , \15669 , \15670 );
or \U$15329 ( \15672 , \15663 , \15671 );
not \U$15330 ( \15673 , \15671 );
not \U$15331 ( \15674 , \15663 );
or \U$15332 ( \15675 , \15673 , \15674 );
and \U$15333 ( \15676 , \2274 , RI9870c90_103);
and \U$15334 ( \15677 , RI9871230_115, \2272 );
nor \U$15335 ( \15678 , \15676 , \15677 );
and \U$15336 ( \15679 , \15678 , \2030 );
not \U$15337 ( \15680 , \15678 );
and \U$15338 ( \15681 , \15680 , \2031 );
nor \U$15339 ( \15682 , \15679 , \15681 );
nand \U$15340 ( \15683 , \15675 , \15682 );
nand \U$15341 ( \15684 , \15672 , \15683 );
and \U$15342 ( \15685 , \776 , RI986fe80_73);
and \U$15343 ( \15686 , RI9870060_77, \774 );
nor \U$15344 ( \15687 , \15685 , \15686 );
and \U$15345 ( \15688 , \15687 , \451 );
not \U$15346 ( \15689 , \15687 );
and \U$15347 ( \15690 , \15689 , \474 );
nor \U$15348 ( \15691 , \15688 , \15690 );
and \U$15349 ( \15692 , \1329 , RI9870ab0_99);
and \U$15350 ( \15693 , RI9870d80_105, \1327 );
nor \U$15351 ( \15694 , \15692 , \15693 );
and \U$15352 ( \15695 , \15694 , \1337 );
not \U$15353 ( \15696 , \15694 );
and \U$15354 ( \15697 , \15696 , \1336 );
nor \U$15355 ( \15698 , \15695 , \15697 );
or \U$15356 ( \15699 , \15691 , \15698 );
not \U$15357 ( \15700 , \15698 );
not \U$15358 ( \15701 , \15691 );
or \U$15359 ( \15702 , \15700 , \15701 );
not \U$15360 ( \15703 , \1128 );
and \U$15361 ( \15704 , \1293 , RI9870150_79);
and \U$15362 ( \15705 , RI9870f60_109, \1291 );
nor \U$15363 ( \15706 , \15704 , \15705 );
not \U$15364 ( \15707 , \15706 );
or \U$15365 ( \15708 , \15703 , \15707 );
or \U$15366 ( \15709 , \15706 , \1128 );
nand \U$15367 ( \15710 , \15708 , \15709 );
nand \U$15368 ( \15711 , \15702 , \15710 );
nand \U$15369 ( \15712 , \15699 , \15711 );
xor \U$15370 ( \15713 , \15684 , \15712 );
and \U$15371 ( \15714 , \2464 , RI9871140_113);
and \U$15372 ( \15715 , RI9871320_117, \2462 );
nor \U$15373 ( \15716 , \15714 , \15715 );
and \U$15374 ( \15717 , \15716 , \2263 );
not \U$15375 ( \15718 , \15716 );
and \U$15376 ( \15719 , \15718 , \2468 );
nor \U$15377 ( \15720 , \15717 , \15719 );
and \U$15378 ( \15721 , \3683 , RI98717d0_127);
and \U$15379 ( \15722 , RI9871500_121, \3681 );
nor \U$15380 ( \15723 , \15721 , \15722 );
not \U$15381 ( \15724 , \15723 );
not \U$15382 ( \15725 , \3412 );
and \U$15383 ( \15726 , \15724 , \15725 );
and \U$15384 ( \15727 , \15723 , \3918 );
nor \U$15385 ( \15728 , \15726 , \15727 );
or \U$15386 ( \15729 , \15720 , \15728 );
not \U$15387 ( \15730 , \15728 );
not \U$15388 ( \15731 , \15720 );
or \U$15389 ( \15732 , \15730 , \15731 );
not \U$15390 ( \15733 , \2935 );
and \U$15391 ( \15734 , \3254 , RI9871410_119);
and \U$15392 ( \15735 , RI98716e0_125, \3252 );
nor \U$15393 ( \15736 , \15734 , \15735 );
not \U$15394 ( \15737 , \15736 );
or \U$15395 ( \15738 , \15733 , \15737 );
or \U$15396 ( \15739 , \15736 , \2935 );
nand \U$15397 ( \15740 , \15738 , \15739 );
nand \U$15398 ( \15741 , \15732 , \15740 );
nand \U$15399 ( \15742 , \15729 , \15741 );
and \U$15400 ( \15743 , \15713 , \15742 );
and \U$15401 ( \15744 , \15684 , \15712 );
or \U$15402 ( \15745 , \15743 , \15744 );
and \U$15403 ( \15746 , \13882 , RI986dcc0_1);
and \U$15404 ( \15747 , RI986e170_11, \13880 );
nor \U$15405 ( \15748 , \15746 , \15747 );
and \U$15406 ( \15749 , \15748 , \13359 );
not \U$15407 ( \15750 , \15748 );
and \U$15408 ( \15751 , \15750 , \13358 );
nor \U$15409 ( \15752 , \15749 , \15751 );
and \U$15410 ( \15753 , \12293 , RI986f610_55);
and \U$15411 ( \15754 , RI986df90_7, \12291 );
nor \U$15412 ( \15755 , \15753 , \15754 );
and \U$15413 ( \15756 , \15755 , \11686 );
not \U$15414 ( \15757 , \15755 );
and \U$15415 ( \15758 , \15757 , \11687 );
nor \U$15416 ( \15759 , \15756 , \15758 );
xor \U$15417 ( \15760 , \15752 , \15759 );
and \U$15418 ( \15761 , \13045 , RI986dea0_5);
and \U$15419 ( \15762 , RI986ddb0_3, \13043 );
nor \U$15420 ( \15763 , \15761 , \15762 );
and \U$15421 ( \15764 , \15763 , \12619 );
not \U$15422 ( \15765 , \15763 );
and \U$15423 ( \15766 , \15765 , \13047 );
nor \U$15424 ( \15767 , \15764 , \15766 );
and \U$15425 ( \15768 , \15760 , \15767 );
and \U$15426 ( \15769 , \15752 , \15759 );
or \U$15427 ( \15770 , \15768 , \15769 );
and \U$15428 ( \15771 , \14937 , RI986e080_9);
and \U$15429 ( \15772 , RI986e260_13, \14935 );
nor \U$15430 ( \15773 , \15771 , \15772 );
and \U$15431 ( \15774 , \15773 , \14538 );
not \U$15432 ( \15775 , \15773 );
and \U$15433 ( \15776 , \15775 , \14539 );
nor \U$15434 ( \15777 , \15774 , \15776 );
not \U$15435 ( \15778 , \15777 );
not \U$15436 ( \15779 , RI9873648_192);
and \U$15437 ( \15780 , \15779 , RI9873558_190);
and \U$15438 ( \15781 , \15780 , RI986e350_15);
nor \U$15439 ( \15782 , \15781 , \14932 );
nand \U$15440 ( \15783 , \15778 , \15782 );
or \U$15441 ( \15784 , \15770 , \15783 );
not \U$15442 ( \15785 , \15783 );
not \U$15443 ( \15786 , \15770 );
or \U$15444 ( \15787 , \15785 , \15786 );
and \U$15445 ( \15788 , \9505 , RI986f700_57);
and \U$15446 ( \15789 , RI986f9d0_63, \9503 );
nor \U$15447 ( \15790 , \15788 , \15789 );
and \U$15448 ( \15791 , \15790 , \9513 );
not \U$15449 ( \15792 , \15790 );
and \U$15450 ( \15793 , \15792 , \9510 );
nor \U$15451 ( \15794 , \15791 , \15793 );
and \U$15452 ( \15795 , \10424 , RI986f8e0_61);
and \U$15453 ( \15796 , RI986f430_51, \10422 );
nor \U$15454 ( \15797 , \15795 , \15796 );
and \U$15455 ( \15798 , \15797 , \10428 );
not \U$15456 ( \15799 , \15797 );
and \U$15457 ( \15800 , \15799 , \9840 );
nor \U$15458 ( \15801 , \15798 , \15800 );
or \U$15459 ( \15802 , \15794 , \15801 );
not \U$15460 ( \15803 , \15801 );
not \U$15461 ( \15804 , \15794 );
or \U$15462 ( \15805 , \15803 , \15804 );
and \U$15463 ( \15806 , \11696 , RI986f340_49);
and \U$15464 ( \15807 , RI986f520_53, \11694 );
nor \U$15465 ( \15808 , \15806 , \15807 );
and \U$15466 ( \15809 , \15808 , \10965 );
not \U$15467 ( \15810 , \15808 );
and \U$15468 ( \15811 , \15810 , \11702 );
nor \U$15469 ( \15812 , \15809 , \15811 );
nand \U$15470 ( \15813 , \15805 , \15812 );
nand \U$15471 ( \15814 , \15802 , \15813 );
nand \U$15472 ( \15815 , \15787 , \15814 );
nand \U$15473 ( \15816 , \15784 , \15815 );
xor \U$15474 ( \15817 , \15745 , \15816 );
and \U$15475 ( \15818 , \6453 , RI986ecb0_35);
and \U$15476 ( \15819 , RI986f070_43, \6451 );
nor \U$15477 ( \15820 , \15818 , \15819 );
and \U$15478 ( \15821 , \15820 , \6180 );
not \U$15479 ( \15822 , \15820 );
and \U$15480 ( \15823 , \15822 , \6190 );
nor \U$15481 ( \15824 , \15821 , \15823 );
and \U$15482 ( \15825 , \7079 , RI986ef80_41);
and \U$15483 ( \15826 , RI986f250_47, \7077 );
nor \U$15484 ( \15827 , \15825 , \15826 );
and \U$15485 ( \15828 , \15827 , \6709 );
not \U$15486 ( \15829 , \15827 );
and \U$15487 ( \15830 , \15829 , \6710 );
nor \U$15488 ( \15831 , \15828 , \15830 );
xor \U$15489 ( \15832 , \15824 , \15831 );
and \U$15490 ( \15833 , \5881 , RI986eda0_37);
and \U$15491 ( \15834 , RI986ebc0_33, \5879 );
nor \U$15492 ( \15835 , \15833 , \15834 );
and \U$15493 ( \15836 , \15835 , \5885 );
not \U$15494 ( \15837 , \15835 );
and \U$15495 ( \15838 , \15837 , \5594 );
nor \U$15496 ( \15839 , \15836 , \15838 );
and \U$15497 ( \15840 , \15832 , \15839 );
and \U$15498 ( \15841 , \15824 , \15831 );
nor \U$15499 ( \15842 , \15840 , \15841 );
and \U$15500 ( \15843 , \4203 , RI98715f0_123);
and \U$15501 ( \15844 , RI986ead0_31, \4201 );
nor \U$15502 ( \15845 , \15843 , \15844 );
and \U$15503 ( \15846 , \15845 , \3922 );
not \U$15504 ( \15847 , \15845 );
and \U$15505 ( \15848 , \15847 , \4207 );
nor \U$15506 ( \15849 , \15846 , \15848 );
and \U$15507 ( \15850 , \4710 , RI986e9e0_29);
and \U$15508 ( \15851 , RI986e8f0_27, \4708 );
nor \U$15509 ( \15852 , \15850 , \15851 );
not \U$15510 ( \15853 , \15852 );
not \U$15511 ( \15854 , \4519 );
and \U$15512 ( \15855 , \15853 , \15854 );
and \U$15513 ( \15856 , \15852 , \4521 );
nor \U$15514 ( \15857 , \15855 , \15856 );
or \U$15515 ( \15858 , \15849 , \15857 );
not \U$15516 ( \15859 , \15857 );
not \U$15517 ( \15860 , \15849 );
or \U$15518 ( \15861 , \15859 , \15860 );
and \U$15519 ( \15862 , \5318 , RI986e800_25);
and \U$15520 ( \15863 , RI986ee90_39, \5316 );
nor \U$15521 ( \15864 , \15862 , \15863 );
and \U$15522 ( \15865 , \15864 , \5052 );
not \U$15523 ( \15866 , \15864 );
and \U$15524 ( \15867 , \15866 , \5322 );
nor \U$15525 ( \15868 , \15865 , \15867 );
nand \U$15526 ( \15869 , \15861 , \15868 );
nand \U$15527 ( \15870 , \15858 , \15869 );
xor \U$15528 ( \15871 , \15842 , \15870 );
and \U$15529 ( \15872 , \7729 , RI986f160_45);
and \U$15530 ( \15873 , RI986e530_19, \7727 );
nor \U$15531 ( \15874 , \15872 , \15873 );
and \U$15532 ( \15875 , \15874 , \7733 );
not \U$15533 ( \15876 , \15874 );
and \U$15534 ( \15877 , \15876 , \7480 );
nor \U$15535 ( \15878 , \15875 , \15877 );
and \U$15536 ( \15879 , \9237 , RI986e620_21);
and \U$15537 ( \15880 , RI986f7f0_59, \9235 );
nor \U$15538 ( \15881 , \15879 , \15880 );
and \U$15539 ( \15882 , \15881 , \8836 );
not \U$15540 ( \15883 , \15881 );
and \U$15541 ( \15884 , \15883 , \9241 );
nor \U$15542 ( \15885 , \15882 , \15884 );
or \U$15543 ( \15886 , \15878 , \15885 );
not \U$15544 ( \15887 , \15885 );
not \U$15545 ( \15888 , \15878 );
or \U$15546 ( \15889 , \15887 , \15888 );
and \U$15547 ( \15890 , \8486 , RI986e440_17);
and \U$15548 ( \15891 , RI986e710_23, \8484 );
nor \U$15549 ( \15892 , \15890 , \15891 );
and \U$15550 ( \15893 , \15892 , \8050 );
not \U$15551 ( \15894 , \15892 );
and \U$15552 ( \15895 , \15894 , \8051 );
nor \U$15553 ( \15896 , \15893 , \15895 );
nand \U$15554 ( \15897 , \15889 , \15896 );
nand \U$15555 ( \15898 , \15886 , \15897 );
and \U$15556 ( \15899 , \15871 , \15898 );
and \U$15557 ( \15900 , \15842 , \15870 );
or \U$15558 ( \15901 , \15899 , \15900 );
and \U$15559 ( \15902 , \15817 , \15901 );
and \U$15560 ( \15903 , \15745 , \15816 );
or \U$15561 ( \15904 , \15902 , \15903 );
not \U$15562 ( \15905 , \15365 );
xor \U$15563 ( \15906 , \15373 , \15383 );
not \U$15564 ( \15907 , \15906 );
or \U$15565 ( \15908 , \15905 , \15907 );
or \U$15566 ( \15909 , \15906 , \15365 );
nand \U$15567 ( \15910 , \15908 , \15909 );
not \U$15568 ( \15911 , \15910 );
xor \U$15569 ( \15912 , \15347 , RI9873558_190);
xor \U$15570 ( \15913 , \15912 , \15355 );
nor \U$15571 ( \15914 , \15911 , \15913 );
xor \U$15572 ( \15915 , \14930 , \14942 );
xor \U$15573 ( \15916 , \15915 , \14950 );
xor \U$15574 ( \15917 , \15914 , \15916 );
not \U$15575 ( \15918 , \15267 );
not \U$15576 ( \15919 , \15278 );
or \U$15577 ( \15920 , \15918 , \15919 );
or \U$15578 ( \15921 , \15267 , \15278 );
nand \U$15579 ( \15922 , \15920 , \15921 );
not \U$15580 ( \15923 , \15922 );
not \U$15581 ( \15924 , \15260 );
and \U$15582 ( \15925 , \15923 , \15924 );
and \U$15583 ( \15926 , \15922 , \15260 );
nor \U$15584 ( \15927 , \15925 , \15926 );
xor \U$15585 ( \15928 , \15393 , \15400 );
xor \U$15586 ( \15929 , \15928 , \15408 );
xor \U$15587 ( \15930 , \15927 , \15929 );
not \U$15588 ( \15931 , \15324 );
not \U$15589 ( \15932 , \15335 );
or \U$15590 ( \15933 , \15931 , \15932 );
or \U$15591 ( \15934 , \15324 , \15335 );
nand \U$15592 ( \15935 , \15933 , \15934 );
not \U$15593 ( \15936 , \15935 );
not \U$15594 ( \15937 , \15317 );
and \U$15595 ( \15938 , \15936 , \15937 );
and \U$15596 ( \15939 , \15935 , \15317 );
nor \U$15597 ( \15940 , \15938 , \15939 );
and \U$15598 ( \15941 , \15930 , \15940 );
and \U$15599 ( \15942 , \15927 , \15929 );
nor \U$15600 ( \15943 , \15941 , \15942 );
and \U$15601 ( \15944 , \15917 , \15943 );
and \U$15602 ( \15945 , \15914 , \15916 );
or \U$15603 ( \15946 , \15944 , \15945 );
xor \U$15604 ( \15947 , \15904 , \15946 );
xor \U$15605 ( \15948 , \15214 , \15222 );
xor \U$15606 ( \15949 , \15948 , \15231 );
xor \U$15607 ( \15950 , \15190 , \15192 );
xor \U$15608 ( \15951 , \15950 , \15200 );
and \U$15609 ( \15952 , \15949 , \15951 );
xor \U$15610 ( \15953 , \15450 , \15457 );
xor \U$15611 ( \15954 , \15953 , \15466 );
xor \U$15612 ( \15955 , \15190 , \15192 );
xor \U$15613 ( \15956 , \15955 , \15200 );
and \U$15614 ( \15957 , \15954 , \15956 );
and \U$15615 ( \15958 , \15949 , \15954 );
or \U$15616 ( \15959 , \15952 , \15957 , \15958 );
and \U$15617 ( \15960 , \465 , RI986fbb0_67);
and \U$15618 ( \15961 , RI986fd90_71, \463 );
nor \U$15619 ( \15962 , \15960 , \15961 );
not \U$15620 ( \15963 , \15962 );
not \U$15621 ( \15964 , \454 );
and \U$15622 ( \15965 , \15963 , \15964 );
and \U$15623 ( \15966 , \15962 , \454 );
nor \U$15624 ( \15967 , \15965 , \15966 );
and \U$15625 ( \15968 , \376 , RI98707e0_93);
and \U$15626 ( \15969 , RI986fac0_65, \374 );
nor \U$15627 ( \15970 , \15968 , \15969 );
not \U$15628 ( \15971 , \15970 );
not \U$15629 ( \15972 , \365 );
and \U$15630 ( \15973 , \15971 , \15972 );
and \U$15631 ( \15974 , \15970 , \365 );
nor \U$15632 ( \15975 , \15973 , \15974 );
or \U$15633 ( \15976 , \15967 , \15975 );
not \U$15634 ( \15977 , \15975 );
not \U$15635 ( \15978 , \15967 );
or \U$15636 ( \15979 , \15977 , \15978 );
and \U$15637 ( \15980 , \438 , RI986fca0_69);
and \U$15638 ( \15981 , RI986ff70_75, \436 );
nor \U$15639 ( \15982 , \15980 , \15981 );
and \U$15640 ( \15983 , \15982 , \444 );
not \U$15641 ( \15984 , \15982 );
and \U$15642 ( \15985 , \15984 , \443 );
nor \U$15643 ( \15986 , \15983 , \15985 );
nand \U$15644 ( \15987 , \15979 , \15986 );
nand \U$15645 ( \15988 , \15976 , \15987 );
and \U$15646 ( \15989 , \354 , RI9870240_81);
and \U$15647 ( \15990 , RI98706f0_91, \352 );
nor \U$15648 ( \15991 , \15989 , \15990 );
not \U$15649 ( \15992 , \15991 );
not \U$15650 ( \15993 , \345 );
and \U$15651 ( \15994 , \15992 , \15993 );
and \U$15652 ( \15995 , \15991 , \345 );
nor \U$15653 ( \15996 , \15994 , \15995 );
and \U$15654 ( \15997 , \416 , RI9870510_87);
and \U$15655 ( \15998 , RI9870330_83, \414 );
nor \U$15656 ( \15999 , \15997 , \15998 );
and \U$15657 ( \16000 , \15999 , \421 );
not \U$15658 ( \16001 , \15999 );
and \U$15659 ( \16002 , \16001 , \422 );
nor \U$15660 ( \16003 , \16000 , \16002 );
or \U$15661 ( \16004 , \15996 , \16003 );
not \U$15662 ( \16005 , \16003 );
not \U$15663 ( \16006 , \15996 );
or \U$15664 ( \16007 , \16005 , \16006 );
not \U$15665 ( \16008 , \386 );
and \U$15666 ( \16009 , \395 , RI9870600_89);
and \U$15667 ( \16010 , RI98708d0_95, \393 );
nor \U$15668 ( \16011 , \16009 , \16010 );
not \U$15669 ( \16012 , \16011 );
or \U$15670 ( \16013 , \16008 , \16012 );
or \U$15671 ( \16014 , \16011 , \487 );
nand \U$15672 ( \16015 , \16013 , \16014 );
nand \U$15673 ( \16016 , \16007 , \16015 );
nand \U$15674 ( \16017 , \16004 , \16016 );
nor \U$15675 ( \16018 , \15988 , \16017 );
not \U$15676 ( \16019 , \16018 );
xor \U$15677 ( \16020 , \15959 , \16019 );
not \U$15678 ( \16021 , \15484 );
not \U$15679 ( \16022 , \15496 );
or \U$15680 ( \16023 , \16021 , \16022 );
or \U$15681 ( \16024 , \15484 , \15496 );
nand \U$15682 ( \16025 , \16023 , \16024 );
not \U$15683 ( \16026 , \16025 );
not \U$15684 ( \16027 , \15477 );
and \U$15685 ( \16028 , \16026 , \16027 );
and \U$15686 ( \16029 , \16025 , \15477 );
nor \U$15687 ( \16030 , \16028 , \16029 );
not \U$15688 ( \16031 , \15430 );
not \U$15689 ( \16032 , \15441 );
or \U$15690 ( \16033 , \16031 , \16032 );
or \U$15691 ( \16034 , \15430 , \15441 );
nand \U$15692 ( \16035 , \16033 , \16034 );
not \U$15693 ( \16036 , \16035 );
not \U$15694 ( \16037 , \15422 );
and \U$15695 ( \16038 , \16036 , \16037 );
and \U$15696 ( \16039 , \16035 , \15422 );
nor \U$15697 ( \16040 , \16038 , \16039 );
xor \U$15698 ( \16041 , \16030 , \16040 );
not \U$15699 ( \16042 , \15295 );
not \U$15700 ( \16043 , \15307 );
or \U$15701 ( \16044 , \16042 , \16043 );
or \U$15702 ( \16045 , \15295 , \15307 );
nand \U$15703 ( \16046 , \16044 , \16045 );
not \U$15704 ( \16047 , \16046 );
not \U$15705 ( \16048 , \15288 );
and \U$15706 ( \16049 , \16047 , \16048 );
and \U$15707 ( \16050 , \16046 , \15288 );
nor \U$15708 ( \16051 , \16049 , \16050 );
and \U$15709 ( \16052 , \16041 , \16051 );
and \U$15710 ( \16053 , \16030 , \16040 );
nor \U$15711 ( \16054 , \16052 , \16053 );
and \U$15712 ( \16055 , \16020 , \16054 );
and \U$15713 ( \16056 , \15959 , \16019 );
or \U$15714 ( \16057 , \16055 , \16056 );
and \U$15715 ( \16058 , \15947 , \16057 );
and \U$15716 ( \16059 , \15904 , \15946 );
or \U$15717 ( \16060 , \16058 , \16059 );
xor \U$15718 ( \16061 , \15656 , \16060 );
xor \U$15719 ( \16062 , \15182 , \15237 );
xor \U$15720 ( \16063 , \16062 , \15250 );
xor \U$15721 ( \16064 , \15517 , \15518 );
xor \U$15722 ( \16065 , \16064 , \15523 );
and \U$15723 ( \16066 , \16063 , \16065 );
xor \U$15724 ( \16067 , \14805 , \14807 );
xor \U$15725 ( \16068 , \16067 , \14810 );
xor \U$15726 ( \16069 , \15532 , \15539 );
xor \U$15727 ( \16070 , \16068 , \16069 );
xor \U$15728 ( \16071 , \15517 , \15518 );
xor \U$15729 ( \16072 , \16071 , \15523 );
and \U$15730 ( \16073 , \16070 , \16072 );
and \U$15731 ( \16074 , \16063 , \16070 );
or \U$15732 ( \16075 , \16066 , \16073 , \16074 );
and \U$15733 ( \16076 , \16061 , \16075 );
and \U$15734 ( \16077 , \15656 , \16060 );
or \U$15735 ( \16078 , \16076 , \16077 );
xor \U$15736 ( \16079 , \14816 , \15068 );
xor \U$15737 ( \16080 , \16079 , \15094 );
xor \U$15738 ( \16081 , \16078 , \16080 );
xor \U$15739 ( \16082 , \14898 , \14982 );
xor \U$15740 ( \16083 , \16082 , \15065 );
xor \U$15741 ( \16084 , \15544 , \15556 );
xor \U$15742 ( \16085 , \16084 , \15561 );
and \U$15743 ( \16086 , \16083 , \16085 );
xor \U$15744 ( \16087 , \15081 , \15086 );
xor \U$15745 ( \16088 , \16087 , \15091 );
xor \U$15746 ( \16089 , \15160 , \15167 );
xor \U$15747 ( \16090 , \16088 , \16089 );
xor \U$15748 ( \16091 , \15544 , \15556 );
xor \U$15749 ( \16092 , \16091 , \15561 );
and \U$15750 ( \16093 , \16090 , \16092 );
and \U$15751 ( \16094 , \16083 , \16090 );
or \U$15752 ( \16095 , \16086 , \16093 , \16094 );
xor \U$15753 ( \16096 , \16081 , \16095 );
and \U$15754 ( \16097 , \15622 , \16096 );
xor \U$15755 ( \16098 , \15842 , \15870 );
xor \U$15756 ( \16099 , \16098 , \15898 );
xor \U$15757 ( \16100 , \15684 , \15712 );
xor \U$15758 ( \16101 , \16100 , \15742 );
and \U$15759 ( \16102 , \16099 , \16101 );
not \U$15760 ( \16103 , \16101 );
not \U$15761 ( \16104 , \16099 );
and \U$15762 ( \16105 , \16103 , \16104 );
not \U$15763 ( \16106 , \15814 );
not \U$15764 ( \16107 , \15770 );
or \U$15765 ( \16108 , \16106 , \16107 );
or \U$15766 ( \16109 , \15770 , \15814 );
nand \U$15767 ( \16110 , \16108 , \16109 );
not \U$15768 ( \16111 , \16110 );
not \U$15769 ( \16112 , \15783 );
and \U$15770 ( \16113 , \16111 , \16112 );
and \U$15771 ( \16114 , \16110 , \15783 );
nor \U$15772 ( \16115 , \16113 , \16114 );
nor \U$15773 ( \16116 , \16105 , \16115 );
nor \U$15774 ( \16117 , \16102 , \16116 );
xor \U$15775 ( \16118 , \15358 , \15385 );
xor \U$15776 ( \16119 , \16118 , \15411 );
or \U$15777 ( \16120 , \16117 , \16119 );
not \U$15778 ( \16121 , \16119 );
not \U$15779 ( \16122 , \16117 );
or \U$15780 ( \16123 , \16121 , \16122 );
xor \U$15781 ( \16124 , \16030 , \16040 );
xor \U$15782 ( \16125 , \16124 , \16051 );
and \U$15783 ( \16126 , \15988 , \16017 );
nor \U$15784 ( \16127 , \16126 , \16018 );
or \U$15785 ( \16128 , \16125 , \16127 );
not \U$15786 ( \16129 , \16127 );
not \U$15787 ( \16130 , \16125 );
or \U$15788 ( \16131 , \16129 , \16130 );
xor \U$15789 ( \16132 , \15190 , \15192 );
xor \U$15790 ( \16133 , \16132 , \15200 );
xor \U$15791 ( \16134 , \15949 , \15954 );
xor \U$15792 ( \16135 , \16133 , \16134 );
nand \U$15793 ( \16136 , \16131 , \16135 );
nand \U$15794 ( \16137 , \16128 , \16136 );
nand \U$15795 ( \16138 , \16123 , \16137 );
nand \U$15796 ( \16139 , \16120 , \16138 );
and \U$15797 ( \16140 , \9505 , RI986f7f0_59);
and \U$15798 ( \16141 , RI986f700_57, \9503 );
nor \U$15799 ( \16142 , \16140 , \16141 );
and \U$15800 ( \16143 , \16142 , \9510 );
not \U$15801 ( \16144 , \16142 );
and \U$15802 ( \16145 , \16144 , \9513 );
nor \U$15803 ( \16146 , \16143 , \16145 );
and \U$15804 ( \16147 , \10424 , RI986f9d0_63);
and \U$15805 ( \16148 , RI986f8e0_61, \10422 );
nor \U$15806 ( \16149 , \16147 , \16148 );
and \U$15807 ( \16150 , \16149 , \9840 );
not \U$15808 ( \16151 , \16149 );
and \U$15809 ( \16152 , \16151 , \10428 );
nor \U$15810 ( \16153 , \16150 , \16152 );
xor \U$15811 ( \16154 , \16146 , \16153 );
and \U$15812 ( \16155 , \9237 , RI986e710_23);
and \U$15813 ( \16156 , RI986e620_21, \9235 );
nor \U$15814 ( \16157 , \16155 , \16156 );
and \U$15815 ( \16158 , \16157 , \9241 );
not \U$15816 ( \16159 , \16157 );
and \U$15817 ( \16160 , \16159 , \8836 );
nor \U$15818 ( \16161 , \16158 , \16160 );
and \U$15819 ( \16162 , \16154 , \16161 );
and \U$15820 ( \16163 , \16146 , \16153 );
nor \U$15821 ( \16164 , \16162 , \16163 );
and \U$15822 ( \16165 , \14937 , RI986e170_11);
and \U$15823 ( \16166 , RI986e080_9, \14935 );
nor \U$15824 ( \16167 , \16165 , \16166 );
and \U$15825 ( \16168 , \16167 , \14538 );
not \U$15826 ( \16169 , \16167 );
and \U$15827 ( \16170 , \16169 , \14539 );
nor \U$15828 ( \16171 , \16168 , \16170 );
and \U$15829 ( \16172 , \15780 , RI986e260_13);
and \U$15830 ( \16173 , RI9873648_192, RI986e350_15);
nor \U$15831 ( \16174 , \16172 , \16173 );
not \U$15832 ( \16175 , \16174 );
not \U$15833 ( \16176 , RI9873558_190);
and \U$15834 ( \16177 , \16175 , \16176 );
and \U$15835 ( \16178 , \16174 , RI9873558_190);
nor \U$15836 ( \16179 , \16177 , \16178 );
xor \U$15837 ( \16180 , \16171 , \16179 );
and \U$15838 ( \16181 , \13882 , RI986ddb0_3);
and \U$15839 ( \16182 , RI986dcc0_1, \13880 );
nor \U$15840 ( \16183 , \16181 , \16182 );
and \U$15841 ( \16184 , \16183 , \13359 );
not \U$15842 ( \16185 , \16183 );
and \U$15843 ( \16186 , \16185 , \13358 );
nor \U$15844 ( \16187 , \16184 , \16186 );
and \U$15845 ( \16188 , \16180 , \16187 );
and \U$15846 ( \16189 , \16171 , \16179 );
or \U$15847 ( \16190 , \16188 , \16189 );
xor \U$15848 ( \16191 , \16164 , \16190 );
and \U$15849 ( \16192 , \12293 , RI986f520_53);
and \U$15850 ( \16193 , RI986f610_55, \12291 );
nor \U$15851 ( \16194 , \16192 , \16193 );
and \U$15852 ( \16195 , \16194 , \11687 );
not \U$15853 ( \16196 , \16194 );
and \U$15854 ( \16197 , \16196 , \11686 );
nor \U$15855 ( \16198 , \16195 , \16197 );
and \U$15856 ( \16199 , \13045 , RI986df90_7);
and \U$15857 ( \16200 , RI986dea0_5, \13043 );
nor \U$15858 ( \16201 , \16199 , \16200 );
and \U$15859 ( \16202 , \16201 , \13047 );
not \U$15860 ( \16203 , \16201 );
and \U$15861 ( \16204 , \16203 , \12619 );
nor \U$15862 ( \16205 , \16202 , \16204 );
xor \U$15863 ( \16206 , \16198 , \16205 );
and \U$15864 ( \16207 , \11696 , RI986f430_51);
and \U$15865 ( \16208 , RI986f340_49, \11694 );
nor \U$15866 ( \16209 , \16207 , \16208 );
and \U$15867 ( \16210 , \16209 , \10965 );
not \U$15868 ( \16211 , \16209 );
and \U$15869 ( \16212 , \16211 , \11702 );
nor \U$15870 ( \16213 , \16210 , \16212 );
and \U$15871 ( \16214 , \16206 , \16213 );
and \U$15872 ( \16215 , \16198 , \16205 );
nor \U$15873 ( \16216 , \16214 , \16215 );
and \U$15874 ( \16217 , \16191 , \16216 );
and \U$15875 ( \16218 , \16164 , \16190 );
or \U$15876 ( \16219 , \16217 , \16218 );
not \U$15877 ( \16220 , \16219 );
and \U$15878 ( \16221 , \2274 , RI9871050_111);
and \U$15879 ( \16222 , RI9870c90_103, \2272 );
nor \U$15880 ( \16223 , \16221 , \16222 );
and \U$15881 ( \16224 , \16223 , \2031 );
not \U$15882 ( \16225 , \16223 );
and \U$15883 ( \16226 , \16225 , \2030 );
nor \U$15884 ( \16227 , \16224 , \16226 );
not \U$15885 ( \16228 , \16227 );
and \U$15886 ( \16229 , \2464 , RI9871230_115);
and \U$15887 ( \16230 , RI9871140_113, \2462 );
nor \U$15888 ( \16231 , \16229 , \16230 );
and \U$15889 ( \16232 , \16231 , \2263 );
not \U$15890 ( \16233 , \16231 );
and \U$15891 ( \16234 , \16233 , \2468 );
nor \U$15892 ( \16235 , \16232 , \16234 );
not \U$15893 ( \16236 , \16235 );
and \U$15894 ( \16237 , \16228 , \16236 );
and \U$15895 ( \16238 , \16235 , \16227 );
and \U$15896 ( \16239 , \3254 , RI9871320_117);
and \U$15897 ( \16240 , RI9871410_119, \3252 );
nor \U$15898 ( \16241 , \16239 , \16240 );
not \U$15899 ( \16242 , \16241 );
not \U$15900 ( \16243 , \3406 );
and \U$15901 ( \16244 , \16242 , \16243 );
and \U$15902 ( \16245 , \16241 , \3406 );
nor \U$15903 ( \16246 , \16244 , \16245 );
nor \U$15904 ( \16247 , \16238 , \16246 );
nor \U$15905 ( \16248 , \16237 , \16247 );
and \U$15906 ( \16249 , \1329 , RI9870f60_109);
and \U$15907 ( \16250 , RI9870ab0_99, \1327 );
nor \U$15908 ( \16251 , \16249 , \16250 );
and \U$15909 ( \16252 , \16251 , \1337 );
not \U$15910 ( \16253 , \16251 );
and \U$15911 ( \16254 , \16253 , \1336 );
nor \U$15912 ( \16255 , \16252 , \16254 );
not \U$15913 ( \16256 , \16255 );
and \U$15914 ( \16257 , \1311 , RI9870d80_105);
and \U$15915 ( \16258 , RI98709c0_97, \1309 );
nor \U$15916 ( \16259 , \16257 , \16258 );
and \U$15917 ( \16260 , \16259 , \1315 );
not \U$15918 ( \16261 , \16259 );
and \U$15919 ( \16262 , \16261 , \1458 );
nor \U$15920 ( \16263 , \16260 , \16262 );
not \U$15921 ( \16264 , \16263 );
and \U$15922 ( \16265 , \16256 , \16264 );
and \U$15923 ( \16266 , \16263 , \16255 );
and \U$15924 ( \16267 , \2042 , RI9870e70_107);
and \U$15925 ( \16268 , RI9870ba0_101, \2040 );
nor \U$15926 ( \16269 , \16267 , \16268 );
not \U$15927 ( \16270 , \16269 );
not \U$15928 ( \16271 , \2034 );
and \U$15929 ( \16272 , \16270 , \16271 );
and \U$15930 ( \16273 , \16269 , \2034 );
nor \U$15931 ( \16274 , \16272 , \16273 );
nor \U$15932 ( \16275 , \16266 , \16274 );
nor \U$15933 ( \16276 , \16265 , \16275 );
xor \U$15934 ( \16277 , \16248 , \16276 );
and \U$15935 ( \16278 , \776 , RI986ff70_75);
and \U$15936 ( \16279 , RI986fe80_73, \774 );
nor \U$15937 ( \16280 , \16278 , \16279 );
and \U$15938 ( \16281 , \16280 , \451 );
not \U$15939 ( \16282 , \16280 );
and \U$15940 ( \16283 , \16282 , \474 );
nor \U$15941 ( \16284 , \16281 , \16283 );
not \U$15942 ( \16285 , \16284 );
and \U$15943 ( \16286 , \438 , RI986fd90_71);
and \U$15944 ( \16287 , RI986fca0_69, \436 );
nor \U$15945 ( \16288 , \16286 , \16287 );
and \U$15946 ( \16289 , \16288 , \443 );
not \U$15947 ( \16290 , \16288 );
and \U$15948 ( \16291 , \16290 , \444 );
nor \U$15949 ( \16292 , \16289 , \16291 );
not \U$15950 ( \16293 , \16292 );
and \U$15951 ( \16294 , \16285 , \16293 );
and \U$15952 ( \16295 , \16292 , \16284 );
and \U$15953 ( \16296 , \1293 , RI9870060_77);
and \U$15954 ( \16297 , RI9870150_79, \1291 );
nor \U$15955 ( \16298 , \16296 , \16297 );
not \U$15956 ( \16299 , \16298 );
not \U$15957 ( \16300 , \1128 );
and \U$15958 ( \16301 , \16299 , \16300 );
and \U$15959 ( \16302 , \16298 , \1301 );
nor \U$15960 ( \16303 , \16301 , \16302 );
nor \U$15961 ( \16304 , \16295 , \16303 );
nor \U$15962 ( \16305 , \16294 , \16304 );
and \U$15963 ( \16306 , \16277 , \16305 );
and \U$15964 ( \16307 , \16248 , \16276 );
or \U$15965 ( \16308 , \16306 , \16307 );
not \U$15966 ( \16309 , \16308 );
and \U$15967 ( \16310 , \16220 , \16309 );
and \U$15968 ( \16311 , \16219 , \16308 );
and \U$15969 ( \16312 , \8486 , RI986e530_19);
and \U$15970 ( \16313 , RI986e440_17, \8484 );
nor \U$15971 ( \16314 , \16312 , \16313 );
and \U$15972 ( \16315 , \16314 , \8050 );
not \U$15973 ( \16316 , \16314 );
and \U$15974 ( \16317 , \16316 , \8051 );
nor \U$15975 ( \16318 , \16315 , \16317 );
and \U$15976 ( \16319 , \7079 , RI986f070_43);
and \U$15977 ( \16320 , RI986ef80_41, \7077 );
nor \U$15978 ( \16321 , \16319 , \16320 );
and \U$15979 ( \16322 , \16321 , \6710 );
not \U$15980 ( \16323 , \16321 );
and \U$15981 ( \16324 , \16323 , \6709 );
nor \U$15982 ( \16325 , \16322 , \16324 );
xor \U$15983 ( \16326 , \16318 , \16325 );
and \U$15984 ( \16327 , \7729 , RI986f250_47);
and \U$15985 ( \16328 , RI986f160_45, \7727 );
nor \U$15986 ( \16329 , \16327 , \16328 );
and \U$15987 ( \16330 , \16329 , \7480 );
not \U$15988 ( \16331 , \16329 );
and \U$15989 ( \16332 , \16331 , \7733 );
nor \U$15990 ( \16333 , \16330 , \16332 );
and \U$15991 ( \16334 , \16326 , \16333 );
and \U$15992 ( \16335 , \16318 , \16325 );
or \U$15993 ( \16336 , \16334 , \16335 );
and \U$15994 ( \16337 , \6453 , RI986ebc0_33);
and \U$15995 ( \16338 , RI986ecb0_35, \6451 );
nor \U$15996 ( \16339 , \16337 , \16338 );
and \U$15997 ( \16340 , \16339 , \6190 );
not \U$15998 ( \16341 , \16339 );
and \U$15999 ( \16342 , \16341 , \6180 );
nor \U$16000 ( \16343 , \16340 , \16342 );
and \U$16001 ( \16344 , \5318 , RI986e8f0_27);
and \U$16002 ( \16345 , RI986e800_25, \5316 );
nor \U$16003 ( \16346 , \16344 , \16345 );
and \U$16004 ( \16347 , \16346 , \5052 );
not \U$16005 ( \16348 , \16346 );
and \U$16006 ( \16349 , \16348 , \5322 );
nor \U$16007 ( \16350 , \16347 , \16349 );
xor \U$16008 ( \16351 , \16343 , \16350 );
and \U$16009 ( \16352 , \5881 , RI986ee90_39);
and \U$16010 ( \16353 , RI986eda0_37, \5879 );
nor \U$16011 ( \16354 , \16352 , \16353 );
and \U$16012 ( \16355 , \16354 , \5594 );
not \U$16013 ( \16356 , \16354 );
and \U$16014 ( \16357 , \16356 , \5885 );
nor \U$16015 ( \16358 , \16355 , \16357 );
and \U$16016 ( \16359 , \16351 , \16358 );
and \U$16017 ( \16360 , \16343 , \16350 );
or \U$16018 ( \16361 , \16359 , \16360 );
xor \U$16019 ( \16362 , \16336 , \16361 );
not \U$16020 ( \16363 , \4521 );
and \U$16021 ( \16364 , \4710 , RI986ead0_31);
and \U$16022 ( \16365 , RI986e9e0_29, \4708 );
nor \U$16023 ( \16366 , \16364 , \16365 );
not \U$16024 ( \16367 , \16366 );
or \U$16025 ( \16368 , \16363 , \16367 );
or \U$16026 ( \16369 , \16366 , \4521 );
nand \U$16027 ( \16370 , \16368 , \16369 );
not \U$16028 ( \16371 , \3412 );
and \U$16029 ( \16372 , \3683 , RI98716e0_125);
and \U$16030 ( \16373 , RI98717d0_127, \3681 );
nor \U$16031 ( \16374 , \16372 , \16373 );
not \U$16032 ( \16375 , \16374 );
or \U$16033 ( \16376 , \16371 , \16375 );
or \U$16034 ( \16377 , \16374 , \3918 );
nand \U$16035 ( \16378 , \16376 , \16377 );
xor \U$16036 ( \16379 , \16370 , \16378 );
and \U$16037 ( \16380 , \4203 , RI9871500_121);
and \U$16038 ( \16381 , RI98715f0_123, \4201 );
nor \U$16039 ( \16382 , \16380 , \16381 );
and \U$16040 ( \16383 , \16382 , \4207 );
not \U$16041 ( \16384 , \16382 );
and \U$16042 ( \16385 , \16384 , \3922 );
nor \U$16043 ( \16386 , \16383 , \16385 );
and \U$16044 ( \16387 , \16379 , \16386 );
and \U$16045 ( \16388 , \16370 , \16378 );
or \U$16046 ( \16389 , \16387 , \16388 );
and \U$16047 ( \16390 , \16362 , \16389 );
and \U$16048 ( \16391 , \16336 , \16361 );
nor \U$16049 ( \16392 , \16390 , \16391 );
nor \U$16050 ( \16393 , \16311 , \16392 );
nor \U$16051 ( \16394 , \16310 , \16393 );
not \U$16052 ( \16395 , \15728 );
not \U$16053 ( \16396 , \15740 );
or \U$16054 ( \16397 , \16395 , \16396 );
or \U$16055 ( \16398 , \15728 , \15740 );
nand \U$16056 ( \16399 , \16397 , \16398 );
not \U$16057 ( \16400 , \16399 );
not \U$16058 ( \16401 , \15720 );
and \U$16059 ( \16402 , \16400 , \16401 );
and \U$16060 ( \16403 , \16399 , \15720 );
nor \U$16061 ( \16404 , \16402 , \16403 );
not \U$16062 ( \16405 , \15857 );
not \U$16063 ( \16406 , \15868 );
or \U$16064 ( \16407 , \16405 , \16406 );
or \U$16065 ( \16408 , \15857 , \15868 );
nand \U$16066 ( \16409 , \16407 , \16408 );
not \U$16067 ( \16410 , \16409 );
not \U$16068 ( \16411 , \15849 );
and \U$16069 ( \16412 , \16410 , \16411 );
and \U$16070 ( \16413 , \16409 , \15849 );
nor \U$16071 ( \16414 , \16412 , \16413 );
xor \U$16072 ( \16415 , \16404 , \16414 );
xor \U$16073 ( \16416 , \15824 , \15831 );
xor \U$16074 ( \16417 , \16416 , \15839 );
and \U$16075 ( \16418 , \16415 , \16417 );
and \U$16076 ( \16419 , \16404 , \16414 );
or \U$16077 ( \16420 , \16418 , \16419 );
and \U$16078 ( \16421 , \465 , RI986fac0_65);
and \U$16079 ( \16422 , RI986fbb0_67, \463 );
nor \U$16080 ( \16423 , \16421 , \16422 );
not \U$16081 ( \16424 , \16423 );
not \U$16082 ( \16425 , \456 );
and \U$16083 ( \16426 , \16424 , \16425 );
and \U$16084 ( \16427 , \16423 , \454 );
nor \U$16085 ( \16428 , \16426 , \16427 );
not \U$16086 ( \16429 , \16428 );
and \U$16087 ( \16430 , \395 , RI98706f0_91);
and \U$16088 ( \16431 , RI9870600_89, \393 );
nor \U$16089 ( \16432 , \16430 , \16431 );
not \U$16090 ( \16433 , \16432 );
not \U$16091 ( \16434 , \386 );
and \U$16092 ( \16435 , \16433 , \16434 );
and \U$16093 ( \16436 , \16432 , \386 );
nor \U$16094 ( \16437 , \16435 , \16436 );
not \U$16095 ( \16438 , \16437 );
and \U$16096 ( \16439 , \16429 , \16438 );
and \U$16097 ( \16440 , \16428 , \16437 );
and \U$16098 ( \16441 , \376 , RI98708d0_95);
and \U$16099 ( \16442 , RI98707e0_93, \374 );
nor \U$16100 ( \16443 , \16441 , \16442 );
not \U$16101 ( \16444 , \16443 );
not \U$16102 ( \16445 , \365 );
and \U$16103 ( \16446 , \16444 , \16445 );
and \U$16104 ( \16447 , \16443 , \367 );
nor \U$16105 ( \16448 , \16446 , \16447 );
nor \U$16106 ( \16449 , \16440 , \16448 );
nor \U$16107 ( \16450 , \16439 , \16449 );
nand \U$16108 ( \16451 , RI9870420_85, RI9871fc8_144);
xor \U$16109 ( \16452 , \16450 , \16451 );
not \U$16110 ( \16453 , \15996 );
not \U$16111 ( \16454 , \16015 );
or \U$16112 ( \16455 , \16453 , \16454 );
or \U$16113 ( \16456 , \15996 , \16015 );
nand \U$16114 ( \16457 , \16455 , \16456 );
not \U$16115 ( \16458 , \16457 );
not \U$16116 ( \16459 , \16003 );
and \U$16117 ( \16460 , \16458 , \16459 );
and \U$16118 ( \16461 , \16457 , \16003 );
nor \U$16119 ( \16462 , \16460 , \16461 );
and \U$16120 ( \16463 , \16452 , \16462 );
and \U$16121 ( \16464 , \16450 , \16451 );
or \U$16122 ( \16465 , \16463 , \16464 );
xor \U$16123 ( \16466 , \16420 , \16465 );
not \U$16124 ( \16467 , \15671 );
not \U$16125 ( \16468 , \15682 );
or \U$16126 ( \16469 , \16467 , \16468 );
or \U$16127 ( \16470 , \15671 , \15682 );
nand \U$16128 ( \16471 , \16469 , \16470 );
not \U$16129 ( \16472 , \16471 );
not \U$16130 ( \16473 , \15663 );
and \U$16131 ( \16474 , \16472 , \16473 );
and \U$16132 ( \16475 , \16471 , \15663 );
nor \U$16133 ( \16476 , \16474 , \16475 );
not \U$16134 ( \16477 , \15967 );
not \U$16135 ( \16478 , \15986 );
or \U$16136 ( \16479 , \16477 , \16478 );
or \U$16137 ( \16480 , \15967 , \15986 );
nand \U$16138 ( \16481 , \16479 , \16480 );
not \U$16139 ( \16482 , \16481 );
not \U$16140 ( \16483 , \15975 );
and \U$16141 ( \16484 , \16482 , \16483 );
and \U$16142 ( \16485 , \16481 , \15975 );
nor \U$16143 ( \16486 , \16484 , \16485 );
xor \U$16144 ( \16487 , \16476 , \16486 );
not \U$16145 ( \16488 , \15698 );
not \U$16146 ( \16489 , \15710 );
or \U$16147 ( \16490 , \16488 , \16489 );
or \U$16148 ( \16491 , \15698 , \15710 );
nand \U$16149 ( \16492 , \16490 , \16491 );
not \U$16150 ( \16493 , \16492 );
not \U$16151 ( \16494 , \15691 );
and \U$16152 ( \16495 , \16493 , \16494 );
and \U$16153 ( \16496 , \16492 , \15691 );
nor \U$16154 ( \16497 , \16495 , \16496 );
and \U$16155 ( \16498 , \16487 , \16497 );
and \U$16156 ( \16499 , \16476 , \16486 );
or \U$16157 ( \16500 , \16498 , \16499 );
and \U$16158 ( \16501 , \16466 , \16500 );
and \U$16159 ( \16502 , \16420 , \16465 );
or \U$16160 ( \16503 , \16501 , \16502 );
xor \U$16161 ( \16504 , \16394 , \16503 );
not \U$16162 ( \16505 , \15885 );
not \U$16163 ( \16506 , \15896 );
or \U$16164 ( \16507 , \16505 , \16506 );
or \U$16165 ( \16508 , \15885 , \15896 );
nand \U$16166 ( \16509 , \16507 , \16508 );
not \U$16167 ( \16510 , \16509 );
not \U$16168 ( \16511 , \15878 );
and \U$16169 ( \16512 , \16510 , \16511 );
and \U$16170 ( \16513 , \16509 , \15878 );
nor \U$16171 ( \16514 , \16512 , \16513 );
not \U$16172 ( \16515 , \15801 );
not \U$16173 ( \16516 , \15812 );
or \U$16174 ( \16517 , \16515 , \16516 );
or \U$16175 ( \16518 , \15801 , \15812 );
nand \U$16176 ( \16519 , \16517 , \16518 );
not \U$16177 ( \16520 , \16519 );
not \U$16178 ( \16521 , \15794 );
and \U$16179 ( \16522 , \16520 , \16521 );
and \U$16180 ( \16523 , \16519 , \15794 );
nor \U$16181 ( \16524 , \16522 , \16523 );
xor \U$16182 ( \16525 , \16514 , \16524 );
xor \U$16183 ( \16526 , \15752 , \15759 );
xor \U$16184 ( \16527 , \16526 , \15767 );
and \U$16185 ( \16528 , \16525 , \16527 );
and \U$16186 ( \16529 , \16514 , \16524 );
or \U$16187 ( \16530 , \16528 , \16529 );
not \U$16188 ( \16531 , \15913 );
not \U$16189 ( \16532 , \15910 );
and \U$16190 ( \16533 , \16531 , \16532 );
and \U$16191 ( \16534 , \15913 , \15910 );
nor \U$16192 ( \16535 , \16533 , \16534 );
xor \U$16193 ( \16536 , \16530 , \16535 );
xor \U$16194 ( \16537 , \15927 , \15929 );
xor \U$16195 ( \16538 , \16537 , \15940 );
and \U$16196 ( \16539 , \16536 , \16538 );
and \U$16197 ( \16540 , \16530 , \16535 );
or \U$16198 ( \16541 , \16539 , \16540 );
and \U$16199 ( \16542 , \16504 , \16541 );
and \U$16200 ( \16543 , \16394 , \16503 );
nor \U$16201 ( \16544 , \16542 , \16543 );
xor \U$16202 ( \16545 , \16139 , \16544 );
xor \U$16203 ( \16546 , \15914 , \15916 );
xor \U$16204 ( \16547 , \16546 , \15943 );
xor \U$16205 ( \16548 , \15640 , \15642 );
xor \U$16206 ( \16549 , \16548 , \15645 );
and \U$16207 ( \16550 , \16547 , \16549 );
xor \U$16208 ( \16551 , \15174 , \15176 );
xor \U$16209 ( \16552 , \16551 , \15179 );
xor \U$16210 ( \16553 , \15626 , \15633 );
xor \U$16211 ( \16554 , \16552 , \16553 );
xor \U$16212 ( \16555 , \15640 , \15642 );
xor \U$16213 ( \16556 , \16555 , \15645 );
and \U$16214 ( \16557 , \16554 , \16556 );
and \U$16215 ( \16558 , \16547 , \16554 );
or \U$16216 ( \16559 , \16550 , \16557 , \16558 );
and \U$16217 ( \16560 , \16545 , \16559 );
and \U$16218 ( \16561 , \16139 , \16544 );
or \U$16219 ( \16562 , \16560 , \16561 );
xor \U$16220 ( \16563 , \15253 , \15504 );
xor \U$16221 ( \16564 , \16563 , \15526 );
xor \U$16222 ( \16565 , \16562 , \16564 );
xor \U$16223 ( \16566 , \15340 , \15414 );
xor \U$16224 ( \16567 , \16566 , \15501 );
xor \U$16225 ( \16568 , \15638 , \15648 );
xor \U$16226 ( \16569 , \16568 , \15653 );
and \U$16227 ( \16570 , \16567 , \16569 );
xor \U$16228 ( \16571 , \15517 , \15518 );
xor \U$16229 ( \16572 , \16571 , \15523 );
xor \U$16230 ( \16573 , \16063 , \16070 );
xor \U$16231 ( \16574 , \16572 , \16573 );
xor \U$16232 ( \16575 , \15638 , \15648 );
xor \U$16233 ( \16576 , \16575 , \15653 );
and \U$16234 ( \16577 , \16574 , \16576 );
and \U$16235 ( \16578 , \16567 , \16574 );
or \U$16236 ( \16579 , \16570 , \16577 , \16578 );
and \U$16237 ( \16580 , \16565 , \16579 );
and \U$16238 ( \16581 , \16562 , \16564 );
or \U$16239 ( \16582 , \16580 , \16581 );
xor \U$16240 ( \16583 , \14722 , \14734 );
xor \U$16241 ( \16584 , \16583 , \14739 );
xor \U$16242 ( \16585 , \15572 , \15585 );
xor \U$16243 ( \16586 , \16584 , \16585 );
xor \U$16244 ( \16587 , \16582 , \16586 );
xor \U$16245 ( \16588 , \15656 , \16060 );
xor \U$16246 ( \16589 , \16588 , \16075 );
xor \U$16247 ( \16590 , \15544 , \15556 );
xor \U$16248 ( \16591 , \16590 , \15561 );
xor \U$16249 ( \16592 , \16083 , \16090 );
xor \U$16250 ( \16593 , \16591 , \16592 );
and \U$16251 ( \16594 , \16589 , \16593 );
and \U$16252 ( \16595 , \16587 , \16594 );
and \U$16253 ( \16596 , \16582 , \16586 );
or \U$16254 ( \16597 , \16595 , \16596 );
xor \U$16255 ( \16598 , \16097 , \16597 );
xor \U$16256 ( \16599 , \15598 , \15600 );
xor \U$16257 ( \16600 , \16599 , \15607 );
xor \U$16258 ( \16601 , \16078 , \16080 );
and \U$16259 ( \16602 , \16601 , \16095 );
and \U$16260 ( \16603 , \16078 , \16080 );
or \U$16261 ( \16604 , \16602 , \16603 );
xor \U$16262 ( \16605 , \15567 , \15569 );
xor \U$16263 ( \16606 , \16605 , \15590 );
xor \U$16264 ( \16607 , \16604 , \16606 );
xor \U$16265 ( \16608 , \16600 , \16607 );
and \U$16266 ( \16609 , \16598 , \16608 );
and \U$16267 ( \16610 , \16097 , \16597 );
or \U$16268 ( \16611 , \16609 , \16610 );
not \U$16269 ( \16612 , \16611 );
xor \U$16270 ( \16613 , \15598 , \15600 );
xor \U$16271 ( \16614 , \16613 , \15607 );
and \U$16272 ( \16615 , \16604 , \16614 );
xor \U$16273 ( \16616 , \15598 , \15600 );
xor \U$16274 ( \16617 , \16616 , \15607 );
and \U$16275 ( \16618 , \16606 , \16617 );
and \U$16276 ( \16619 , \16604 , \16606 );
or \U$16277 ( \16620 , \16615 , \16618 , \16619 );
not \U$16278 ( \16621 , \14692 );
xor \U$16279 ( \16622 , \15124 , \14705 );
not \U$16280 ( \16623 , \16622 );
or \U$16281 ( \16624 , \16621 , \16623 );
or \U$16282 ( \16625 , \16622 , \14692 );
nand \U$16283 ( \16626 , \16624 , \16625 );
xor \U$16284 ( \16627 , \16620 , \16626 );
xor \U$16285 ( \16628 , \15593 , \15595 );
xor \U$16286 ( \16629 , \16628 , \15610 );
xor \U$16287 ( \16630 , \16627 , \16629 );
not \U$16288 ( \16631 , \16630 );
or \U$16289 ( \16632 , \16612 , \16631 );
xor \U$16290 ( \16633 , \15745 , \15816 );
xor \U$16291 ( \16634 , \16633 , \15901 );
xor \U$16292 ( \16635 , \15959 , \16019 );
xor \U$16293 ( \16636 , \16635 , \16054 );
and \U$16294 ( \16637 , \16634 , \16636 );
xor \U$16295 ( \16638 , \15640 , \15642 );
xor \U$16296 ( \16639 , \16638 , \15645 );
xor \U$16297 ( \16640 , \16547 , \16554 );
xor \U$16298 ( \16641 , \16639 , \16640 );
xor \U$16299 ( \16642 , \15959 , \16019 );
xor \U$16300 ( \16643 , \16642 , \16054 );
and \U$16301 ( \16644 , \16641 , \16643 );
and \U$16302 ( \16645 , \16634 , \16641 );
or \U$16303 ( \16646 , \16637 , \16644 , \16645 );
xor \U$16304 ( \16647 , \15904 , \15946 );
xor \U$16305 ( \16648 , \16647 , \16057 );
xor \U$16306 ( \16649 , \16646 , \16648 );
not \U$16307 ( \16650 , \2034 );
and \U$16308 ( \16651 , \2042 , RI98709c0_97);
and \U$16309 ( \16652 , RI9870e70_107, \2040 );
nor \U$16310 ( \16653 , \16651 , \16652 );
not \U$16311 ( \16654 , \16653 );
or \U$16312 ( \16655 , \16650 , \16654 );
or \U$16313 ( \16656 , \16653 , \1462 );
nand \U$16314 ( \16657 , \16655 , \16656 );
and \U$16315 ( \16658 , \2274 , RI9870ba0_101);
and \U$16316 ( \16659 , RI9871050_111, \2272 );
nor \U$16317 ( \16660 , \16658 , \16659 );
and \U$16318 ( \16661 , \16660 , \2030 );
not \U$16319 ( \16662 , \16660 );
and \U$16320 ( \16663 , \16662 , \2031 );
nor \U$16321 ( \16664 , \16661 , \16663 );
xor \U$16322 ( \16665 , \16657 , \16664 );
and \U$16323 ( \16666 , \1311 , RI9870ab0_99);
and \U$16324 ( \16667 , RI9870d80_105, \1309 );
nor \U$16325 ( \16668 , \16666 , \16667 );
and \U$16326 ( \16669 , \16668 , \1458 );
not \U$16327 ( \16670 , \16668 );
and \U$16328 ( \16671 , \16670 , \1318 );
nor \U$16329 ( \16672 , \16669 , \16671 );
and \U$16330 ( \16673 , \16665 , \16672 );
and \U$16331 ( \16674 , \16657 , \16664 );
nor \U$16332 ( \16675 , \16673 , \16674 );
and \U$16333 ( \16676 , \2464 , RI9870c90_103);
and \U$16334 ( \16677 , RI9871230_115, \2462 );
nor \U$16335 ( \16678 , \16676 , \16677 );
and \U$16336 ( \16679 , \16678 , \2263 );
not \U$16337 ( \16680 , \16678 );
and \U$16338 ( \16681 , \16680 , \2468 );
nor \U$16339 ( \16682 , \16679 , \16681 );
not \U$16340 ( \16683 , \16682 );
and \U$16341 ( \16684 , \3254 , RI9871140_113);
and \U$16342 ( \16685 , RI9871320_117, \3252 );
nor \U$16343 ( \16686 , \16684 , \16685 );
not \U$16344 ( \16687 , \16686 );
not \U$16345 ( \16688 , \2935 );
and \U$16346 ( \16689 , \16687 , \16688 );
and \U$16347 ( \16690 , \16686 , \2935 );
nor \U$16348 ( \16691 , \16689 , \16690 );
not \U$16349 ( \16692 , \16691 );
and \U$16350 ( \16693 , \16683 , \16692 );
and \U$16351 ( \16694 , \16691 , \16682 );
and \U$16352 ( \16695 , \3683 , RI9871410_119);
and \U$16353 ( \16696 , RI98716e0_125, \3681 );
nor \U$16354 ( \16697 , \16695 , \16696 );
not \U$16355 ( \16698 , \16697 );
not \U$16356 ( \16699 , \3918 );
and \U$16357 ( \16700 , \16698 , \16699 );
and \U$16358 ( \16701 , \16697 , \3412 );
nor \U$16359 ( \16702 , \16700 , \16701 );
nor \U$16360 ( \16703 , \16694 , \16702 );
nor \U$16361 ( \16704 , \16693 , \16703 );
xor \U$16362 ( \16705 , \16675 , \16704 );
and \U$16363 ( \16706 , \776 , RI986fca0_69);
and \U$16364 ( \16707 , RI986ff70_75, \774 );
nor \U$16365 ( \16708 , \16706 , \16707 );
and \U$16366 ( \16709 , \16708 , \451 );
not \U$16367 ( \16710 , \16708 );
and \U$16368 ( \16711 , \16710 , \474 );
nor \U$16369 ( \16712 , \16709 , \16711 );
not \U$16370 ( \16713 , \16712 );
and \U$16371 ( \16714 , \1293 , RI986fe80_73);
and \U$16372 ( \16715 , RI9870060_77, \1291 );
nor \U$16373 ( \16716 , \16714 , \16715 );
not \U$16374 ( \16717 , \16716 );
not \U$16375 ( \16718 , \1301 );
and \U$16376 ( \16719 , \16717 , \16718 );
and \U$16377 ( \16720 , \16716 , \1128 );
nor \U$16378 ( \16721 , \16719 , \16720 );
not \U$16379 ( \16722 , \16721 );
and \U$16380 ( \16723 , \16713 , \16722 );
and \U$16381 ( \16724 , \16721 , \16712 );
and \U$16382 ( \16725 , \1329 , RI9870150_79);
and \U$16383 ( \16726 , RI9870f60_109, \1327 );
nor \U$16384 ( \16727 , \16725 , \16726 );
and \U$16385 ( \16728 , \16727 , \1337 );
not \U$16386 ( \16729 , \16727 );
and \U$16387 ( \16730 , \16729 , \1336 );
nor \U$16388 ( \16731 , \16728 , \16730 );
nor \U$16389 ( \16732 , \16724 , \16731 );
nor \U$16390 ( \16733 , \16723 , \16732 );
and \U$16391 ( \16734 , \16705 , \16733 );
and \U$16392 ( \16735 , \16675 , \16704 );
nor \U$16393 ( \16736 , \16734 , \16735 );
and \U$16394 ( \16737 , \15780 , RI986e080_9);
and \U$16395 ( \16738 , RI9873648_192, RI986e260_13);
nor \U$16396 ( \16739 , \16737 , \16738 );
not \U$16397 ( \16740 , \16739 );
not \U$16398 ( \16741 , RI9873558_190);
and \U$16399 ( \16742 , \16740 , \16741 );
and \U$16400 ( \16743 , \16739 , RI9873558_190);
nor \U$16401 ( \16744 , \16742 , \16743 );
not \U$16402 ( \16745 , \16744 );
not \U$16403 ( \16746 , \422 );
and \U$16404 ( \16747 , \16745 , \16746 );
and \U$16405 ( \16748 , \16744 , \422 );
and \U$16406 ( \16749 , \14937 , RI986dcc0_1);
and \U$16407 ( \16750 , RI986e170_11, \14935 );
nor \U$16408 ( \16751 , \16749 , \16750 );
and \U$16409 ( \16752 , \16751 , \14538 );
not \U$16410 ( \16753 , \16751 );
and \U$16411 ( \16754 , \16753 , \14539 );
nor \U$16412 ( \16755 , \16752 , \16754 );
nor \U$16413 ( \16756 , \16748 , \16755 );
nor \U$16414 ( \16757 , \16747 , \16756 );
and \U$16415 ( \16758 , \9505 , RI986e620_21);
and \U$16416 ( \16759 , RI986f7f0_59, \9503 );
nor \U$16417 ( \16760 , \16758 , \16759 );
and \U$16418 ( \16761 , \16760 , \9513 );
not \U$16419 ( \16762 , \16760 );
and \U$16420 ( \16763 , \16762 , \9510 );
nor \U$16421 ( \16764 , \16761 , \16763 );
not \U$16422 ( \16765 , \16764 );
and \U$16423 ( \16766 , \10424 , RI986f700_57);
and \U$16424 ( \16767 , RI986f9d0_63, \10422 );
nor \U$16425 ( \16768 , \16766 , \16767 );
and \U$16426 ( \16769 , \16768 , \10428 );
not \U$16427 ( \16770 , \16768 );
and \U$16428 ( \16771 , \16770 , \9840 );
nor \U$16429 ( \16772 , \16769 , \16771 );
not \U$16430 ( \16773 , \16772 );
and \U$16431 ( \16774 , \16765 , \16773 );
and \U$16432 ( \16775 , \16772 , \16764 );
and \U$16433 ( \16776 , \11696 , RI986f8e0_61);
and \U$16434 ( \16777 , RI986f430_51, \11694 );
nor \U$16435 ( \16778 , \16776 , \16777 );
and \U$16436 ( \16779 , \16778 , \11702 );
not \U$16437 ( \16780 , \16778 );
and \U$16438 ( \16781 , \16780 , \10965 );
nor \U$16439 ( \16782 , \16779 , \16781 );
nor \U$16440 ( \16783 , \16775 , \16782 );
nor \U$16441 ( \16784 , \16774 , \16783 );
xor \U$16442 ( \16785 , \16757 , \16784 );
and \U$16443 ( \16786 , \12293 , RI986f340_49);
and \U$16444 ( \16787 , RI986f520_53, \12291 );
nor \U$16445 ( \16788 , \16786 , \16787 );
and \U$16446 ( \16789 , \16788 , \11686 );
not \U$16447 ( \16790 , \16788 );
and \U$16448 ( \16791 , \16790 , \11687 );
nor \U$16449 ( \16792 , \16789 , \16791 );
not \U$16450 ( \16793 , \16792 );
and \U$16451 ( \16794 , \13045 , RI986f610_55);
and \U$16452 ( \16795 , RI986df90_7, \13043 );
nor \U$16453 ( \16796 , \16794 , \16795 );
and \U$16454 ( \16797 , \16796 , \12619 );
not \U$16455 ( \16798 , \16796 );
and \U$16456 ( \16799 , \16798 , \13047 );
nor \U$16457 ( \16800 , \16797 , \16799 );
not \U$16458 ( \16801 , \16800 );
and \U$16459 ( \16802 , \16793 , \16801 );
and \U$16460 ( \16803 , \16800 , \16792 );
and \U$16461 ( \16804 , \13882 , RI986dea0_5);
and \U$16462 ( \16805 , RI986ddb0_3, \13880 );
nor \U$16463 ( \16806 , \16804 , \16805 );
and \U$16464 ( \16807 , \16806 , \13359 );
not \U$16465 ( \16808 , \16806 );
and \U$16466 ( \16809 , \16808 , \13358 );
nor \U$16467 ( \16810 , \16807 , \16809 );
nor \U$16468 ( \16811 , \16803 , \16810 );
nor \U$16469 ( \16812 , \16802 , \16811 );
and \U$16470 ( \16813 , \16785 , \16812 );
and \U$16471 ( \16814 , \16757 , \16784 );
nor \U$16472 ( \16815 , \16813 , \16814 );
xor \U$16473 ( \16816 , \16736 , \16815 );
not \U$16474 ( \16817 , \4519 );
and \U$16475 ( \16818 , \4710 , RI98715f0_123);
and \U$16476 ( \16819 , RI986ead0_31, \4708 );
nor \U$16477 ( \16820 , \16818 , \16819 );
not \U$16478 ( \16821 , \16820 );
or \U$16479 ( \16822 , \16817 , \16821 );
or \U$16480 ( \16823 , \16820 , \4521 );
nand \U$16481 ( \16824 , \16822 , \16823 );
and \U$16482 ( \16825 , \5318 , RI986e9e0_29);
and \U$16483 ( \16826 , RI986e8f0_27, \5316 );
nor \U$16484 ( \16827 , \16825 , \16826 );
and \U$16485 ( \16828 , \16827 , \5052 );
not \U$16486 ( \16829 , \16827 );
and \U$16487 ( \16830 , \16829 , \5322 );
nor \U$16488 ( \16831 , \16828 , \16830 );
xor \U$16489 ( \16832 , \16824 , \16831 );
and \U$16490 ( \16833 , \4203 , RI98717d0_127);
and \U$16491 ( \16834 , RI9871500_121, \4201 );
nor \U$16492 ( \16835 , \16833 , \16834 );
and \U$16493 ( \16836 , \16835 , \4207 );
not \U$16494 ( \16837 , \16835 );
and \U$16495 ( \16838 , \16837 , \3923 );
nor \U$16496 ( \16839 , \16836 , \16838 );
and \U$16497 ( \16840 , \16832 , \16839 );
and \U$16498 ( \16841 , \16824 , \16831 );
nor \U$16499 ( \16842 , \16840 , \16841 );
and \U$16500 ( \16843 , \7729 , RI986ef80_41);
and \U$16501 ( \16844 , RI986f250_47, \7727 );
nor \U$16502 ( \16845 , \16843 , \16844 );
and \U$16503 ( \16846 , \16845 , \7733 );
not \U$16504 ( \16847 , \16845 );
and \U$16505 ( \16848 , \16847 , \7480 );
nor \U$16506 ( \16849 , \16846 , \16848 );
not \U$16507 ( \16850 , \16849 );
and \U$16508 ( \16851 , \9237 , RI986e440_17);
and \U$16509 ( \16852 , RI986e710_23, \9235 );
nor \U$16510 ( \16853 , \16851 , \16852 );
and \U$16511 ( \16854 , \16853 , \8836 );
not \U$16512 ( \16855 , \16853 );
and \U$16513 ( \16856 , \16855 , \9241 );
nor \U$16514 ( \16857 , \16854 , \16856 );
not \U$16515 ( \16858 , \16857 );
and \U$16516 ( \16859 , \16850 , \16858 );
and \U$16517 ( \16860 , \16857 , \16849 );
and \U$16518 ( \16861 , \8486 , RI986f160_45);
and \U$16519 ( \16862 , RI986e530_19, \8484 );
nor \U$16520 ( \16863 , \16861 , \16862 );
and \U$16521 ( \16864 , \16863 , \8051 );
not \U$16522 ( \16865 , \16863 );
and \U$16523 ( \16866 , \16865 , \8050 );
nor \U$16524 ( \16867 , \16864 , \16866 );
nor \U$16525 ( \16868 , \16860 , \16867 );
nor \U$16526 ( \16869 , \16859 , \16868 );
or \U$16527 ( \16870 , \16842 , \16869 );
not \U$16528 ( \16871 , \16842 );
not \U$16529 ( \16872 , \16869 );
or \U$16530 ( \16873 , \16871 , \16872 );
and \U$16531 ( \16874 , \7079 , RI986ecb0_35);
and \U$16532 ( \16875 , RI986f070_43, \7077 );
nor \U$16533 ( \16876 , \16874 , \16875 );
and \U$16534 ( \16877 , \16876 , \6710 );
not \U$16535 ( \16878 , \16876 );
and \U$16536 ( \16879 , \16878 , \6709 );
nor \U$16537 ( \16880 , \16877 , \16879 );
and \U$16538 ( \16881 , \5881 , RI986e800_25);
and \U$16539 ( \16882 , RI986ee90_39, \5879 );
nor \U$16540 ( \16883 , \16881 , \16882 );
and \U$16541 ( \16884 , \16883 , \5594 );
not \U$16542 ( \16885 , \16883 );
and \U$16543 ( \16886 , \16885 , \5885 );
nor \U$16544 ( \16887 , \16884 , \16886 );
xor \U$16545 ( \16888 , \16880 , \16887 );
and \U$16546 ( \16889 , \6453 , RI986eda0_37);
and \U$16547 ( \16890 , RI986ebc0_33, \6451 );
nor \U$16548 ( \16891 , \16889 , \16890 );
and \U$16549 ( \16892 , \16891 , \6190 );
not \U$16550 ( \16893 , \16891 );
and \U$16551 ( \16894 , \16893 , \6705 );
nor \U$16552 ( \16895 , \16892 , \16894 );
and \U$16553 ( \16896 , \16888 , \16895 );
and \U$16554 ( \16897 , \16880 , \16887 );
or \U$16555 ( \16898 , \16896 , \16897 );
nand \U$16556 ( \16899 , \16873 , \16898 );
nand \U$16557 ( \16900 , \16870 , \16899 );
and \U$16558 ( \16901 , \16816 , \16900 );
and \U$16559 ( \16902 , \16736 , \16815 );
nor \U$16560 ( \16903 , \16901 , \16902 );
not \U$16561 ( \16904 , \16903 );
xor \U$16562 ( \16905 , \16171 , \16179 );
xor \U$16563 ( \16906 , \16905 , \16187 );
not \U$16564 ( \16907 , \16906 );
xor \U$16565 ( \16908 , \16198 , \16205 );
xor \U$16566 ( \16909 , \16908 , \16213 );
nand \U$16567 ( \16910 , \16907 , \16909 );
not \U$16568 ( \16911 , \15777 );
not \U$16569 ( \16912 , \15782 );
and \U$16570 ( \16913 , \16911 , \16912 );
and \U$16571 ( \16914 , \15777 , \15782 );
nor \U$16572 ( \16915 , \16913 , \16914 );
xor \U$16573 ( \16916 , \16910 , \16915 );
xor \U$16574 ( \16917 , \16146 , \16153 );
xor \U$16575 ( \16918 , \16917 , \16161 );
xor \U$16576 ( \16919 , \16318 , \16325 );
xor \U$16577 ( \16920 , \16919 , \16333 );
and \U$16578 ( \16921 , \16918 , \16920 );
xor \U$16579 ( \16922 , \16343 , \16350 );
xor \U$16580 ( \16923 , \16922 , \16358 );
xor \U$16581 ( \16924 , \16318 , \16325 );
xor \U$16582 ( \16925 , \16924 , \16333 );
and \U$16583 ( \16926 , \16923 , \16925 );
and \U$16584 ( \16927 , \16918 , \16923 );
or \U$16585 ( \16928 , \16921 , \16926 , \16927 );
not \U$16586 ( \16929 , \16928 );
and \U$16587 ( \16930 , \16916 , \16929 );
and \U$16588 ( \16931 , \16910 , \16915 );
or \U$16589 ( \16932 , \16930 , \16931 );
not \U$16590 ( \16933 , \16932 );
and \U$16591 ( \16934 , \16904 , \16933 );
and \U$16592 ( \16935 , \16903 , \16932 );
not \U$16593 ( \16936 , \16437 );
xor \U$16594 ( \16937 , \16428 , \16448 );
not \U$16595 ( \16938 , \16937 );
or \U$16596 ( \16939 , \16936 , \16938 );
or \U$16597 ( \16940 , \16937 , \16437 );
nand \U$16598 ( \16941 , \16939 , \16940 );
and \U$16599 ( \16942 , \416 , RI9870420_85);
and \U$16600 ( \16943 , RI9870510_87, \414 );
nor \U$16601 ( \16944 , \16942 , \16943 );
and \U$16602 ( \16945 , \16944 , \422 );
not \U$16603 ( \16946 , \16944 );
and \U$16604 ( \16947 , \16946 , \421 );
nor \U$16605 ( \16948 , \16945 , \16947 );
xor \U$16606 ( \16949 , \16941 , \16948 );
not \U$16607 ( \16950 , \16292 );
xor \U$16608 ( \16951 , \16284 , \16303 );
not \U$16609 ( \16952 , \16951 );
or \U$16610 ( \16953 , \16950 , \16952 );
or \U$16611 ( \16954 , \16951 , \16292 );
nand \U$16612 ( \16955 , \16953 , \16954 );
and \U$16613 ( \16956 , \16949 , \16955 );
and \U$16614 ( \16957 , \16941 , \16948 );
or \U$16615 ( \16958 , \16956 , \16957 );
not \U$16616 ( \16959 , \386 );
and \U$16617 ( \16960 , \395 , RI9870240_81);
and \U$16618 ( \16961 , RI98706f0_91, \393 );
nor \U$16619 ( \16962 , \16960 , \16961 );
not \U$16620 ( \16963 , \16962 );
or \U$16621 ( \16964 , \16959 , \16963 );
or \U$16622 ( \16965 , \16962 , \386 );
nand \U$16623 ( \16966 , \16964 , \16965 );
nand \U$16624 ( \16967 , RI9870420_85, \414 );
and \U$16625 ( \16968 , \16967 , \422 );
not \U$16626 ( \16969 , \16967 );
and \U$16627 ( \16970 , \16969 , \421 );
nor \U$16628 ( \16971 , \16968 , \16970 );
xor \U$16629 ( \16972 , \16966 , \16971 );
not \U$16630 ( \16973 , \345 );
and \U$16631 ( \16974 , \354 , RI9870510_87);
and \U$16632 ( \16975 , RI9870330_83, \352 );
nor \U$16633 ( \16976 , \16974 , \16975 );
not \U$16634 ( \16977 , \16976 );
or \U$16635 ( \16978 , \16973 , \16977 );
or \U$16636 ( \16979 , \16976 , \345 );
nand \U$16637 ( \16980 , \16978 , \16979 );
and \U$16638 ( \16981 , \16972 , \16980 );
and \U$16639 ( \16982 , \16966 , \16971 );
or \U$16640 ( \16983 , \16981 , \16982 );
not \U$16641 ( \16984 , \345 );
and \U$16642 ( \16985 , \354 , RI9870330_83);
and \U$16643 ( \16986 , RI9870240_81, \352 );
nor \U$16644 ( \16987 , \16985 , \16986 );
not \U$16645 ( \16988 , \16987 );
or \U$16646 ( \16989 , \16984 , \16988 );
or \U$16647 ( \16990 , \16987 , \361 );
nand \U$16648 ( \16991 , \16989 , \16990 );
xor \U$16649 ( \16992 , \16983 , \16991 );
and \U$16650 ( \16993 , \438 , RI986fbb0_67);
and \U$16651 ( \16994 , RI986fd90_71, \436 );
nor \U$16652 ( \16995 , \16993 , \16994 );
and \U$16653 ( \16996 , \16995 , \444 );
not \U$16654 ( \16997 , \16995 );
and \U$16655 ( \16998 , \16997 , \443 );
nor \U$16656 ( \16999 , \16996 , \16998 );
not \U$16657 ( \17000 , \456 );
and \U$16658 ( \17001 , \465 , RI98707e0_93);
and \U$16659 ( \17002 , RI986fac0_65, \463 );
nor \U$16660 ( \17003 , \17001 , \17002 );
not \U$16661 ( \17004 , \17003 );
or \U$16662 ( \17005 , \17000 , \17004 );
or \U$16663 ( \17006 , \17003 , \454 );
nand \U$16664 ( \17007 , \17005 , \17006 );
xor \U$16665 ( \17008 , \16999 , \17007 );
not \U$16666 ( \17009 , \367 );
and \U$16667 ( \17010 , \376 , RI9870600_89);
and \U$16668 ( \17011 , RI98708d0_95, \374 );
nor \U$16669 ( \17012 , \17010 , \17011 );
not \U$16670 ( \17013 , \17012 );
or \U$16671 ( \17014 , \17009 , \17013 );
or \U$16672 ( \17015 , \17012 , \365 );
nand \U$16673 ( \17016 , \17014 , \17015 );
and \U$16674 ( \17017 , \17008 , \17016 );
and \U$16675 ( \17018 , \16999 , \17007 );
or \U$16676 ( \17019 , \17017 , \17018 );
and \U$16677 ( \17020 , \16992 , \17019 );
and \U$16678 ( \17021 , \16983 , \16991 );
or \U$16679 ( \17022 , \17020 , \17021 );
xor \U$16680 ( \17023 , \16958 , \17022 );
not \U$16681 ( \17024 , \16255 );
xor \U$16682 ( \17025 , \16263 , \16274 );
not \U$16683 ( \17026 , \17025 );
or \U$16684 ( \17027 , \17024 , \17026 );
or \U$16685 ( \17028 , \17025 , \16255 );
nand \U$16686 ( \17029 , \17027 , \17028 );
xor \U$16687 ( \17030 , \16370 , \16378 );
xor \U$16688 ( \17031 , \17030 , \16386 );
and \U$16689 ( \17032 , \17029 , \17031 );
not \U$16690 ( \17033 , \16227 );
xor \U$16691 ( \17034 , \16235 , \16246 );
not \U$16692 ( \17035 , \17034 );
or \U$16693 ( \17036 , \17033 , \17035 );
or \U$16694 ( \17037 , \17034 , \16227 );
nand \U$16695 ( \17038 , \17036 , \17037 );
xor \U$16696 ( \17039 , \16370 , \16378 );
xor \U$16697 ( \17040 , \17039 , \16386 );
and \U$16698 ( \17041 , \17038 , \17040 );
and \U$16699 ( \17042 , \17029 , \17038 );
or \U$16700 ( \17043 , \17032 , \17041 , \17042 );
and \U$16701 ( \17044 , \17023 , \17043 );
and \U$16702 ( \17045 , \16958 , \17022 );
nor \U$16703 ( \17046 , \17044 , \17045 );
nor \U$16704 ( \17047 , \16935 , \17046 );
nor \U$16705 ( \17048 , \16934 , \17047 );
not \U$16706 ( \17049 , \16115 );
xor \U$16707 ( \17050 , \16099 , \16101 );
not \U$16708 ( \17051 , \17050 );
or \U$16709 ( \17052 , \17049 , \17051 );
or \U$16710 ( \17053 , \17050 , \16115 );
nand \U$16711 ( \17054 , \17052 , \17053 );
xor \U$16712 ( \17055 , \16248 , \16276 );
xor \U$16713 ( \17056 , \17055 , \16305 );
xor \U$16714 ( \17057 , \16450 , \16451 );
xor \U$16715 ( \17058 , \17057 , \16462 );
or \U$16716 ( \17059 , \17056 , \17058 );
not \U$16717 ( \17060 , \17058 );
not \U$16718 ( \17061 , \17056 );
or \U$16719 ( \17062 , \17060 , \17061 );
xor \U$16720 ( \17063 , \16336 , \16361 );
xor \U$16721 ( \17064 , \17063 , \16389 );
nand \U$16722 ( \17065 , \17062 , \17064 );
nand \U$16723 ( \17066 , \17059 , \17065 );
xor \U$16724 ( \17067 , \17054 , \17066 );
xor \U$16725 ( \17068 , \16476 , \16486 );
xor \U$16726 ( \17069 , \17068 , \16497 );
xor \U$16727 ( \17070 , \16514 , \16524 );
xor \U$16728 ( \17071 , \17070 , \16527 );
xor \U$16729 ( \17072 , \17069 , \17071 );
xor \U$16730 ( \17073 , \16404 , \16414 );
xor \U$16731 ( \17074 , \17073 , \16417 );
and \U$16732 ( \17075 , \17072 , \17074 );
and \U$16733 ( \17076 , \17069 , \17071 );
nor \U$16734 ( \17077 , \17075 , \17076 );
and \U$16735 ( \17078 , \17067 , \17077 );
and \U$16736 ( \17079 , \17054 , \17066 );
nor \U$16737 ( \17080 , \17078 , \17079 );
xor \U$16738 ( \17081 , \17048 , \17080 );
xor \U$16739 ( \17082 , \16530 , \16535 );
xor \U$16740 ( \17083 , \17082 , \16538 );
not \U$16741 ( \17084 , \17083 );
xor \U$16742 ( \17085 , \16420 , \16465 );
xor \U$16743 ( \17086 , \17085 , \16500 );
not \U$16744 ( \17087 , \17086 );
and \U$16745 ( \17088 , \17084 , \17087 );
and \U$16746 ( \17089 , \17083 , \17086 );
not \U$16747 ( \17090 , \16125 );
not \U$16748 ( \17091 , \16135 );
or \U$16749 ( \17092 , \17090 , \17091 );
or \U$16750 ( \17093 , \16135 , \16125 );
nand \U$16751 ( \17094 , \17092 , \17093 );
not \U$16752 ( \17095 , \17094 );
not \U$16753 ( \17096 , \16127 );
and \U$16754 ( \17097 , \17095 , \17096 );
and \U$16755 ( \17098 , \17094 , \16127 );
nor \U$16756 ( \17099 , \17097 , \17098 );
nor \U$16757 ( \17100 , \17089 , \17099 );
nor \U$16758 ( \17101 , \17088 , \17100 );
and \U$16759 ( \17102 , \17081 , \17101 );
and \U$16760 ( \17103 , \17048 , \17080 );
nor \U$16761 ( \17104 , \17102 , \17103 );
and \U$16762 ( \17105 , \16649 , \17104 );
and \U$16763 ( \17106 , \16646 , \16648 );
or \U$16764 ( \17107 , \17105 , \17106 );
xor \U$16765 ( \17108 , \16562 , \16564 );
xor \U$16766 ( \17109 , \17108 , \16579 );
xnor \U$16767 ( \17110 , \17107 , \17109 );
not \U$16768 ( \17111 , \17110 );
xor \U$16769 ( \17112 , \16589 , \16593 );
not \U$16770 ( \17113 , \17112 );
and \U$16771 ( \17114 , \17111 , \17113 );
and \U$16772 ( \17115 , \17110 , \17112 );
nor \U$16773 ( \17116 , \17114 , \17115 );
not \U$16774 ( \17117 , \17116 );
xor \U$16775 ( \17118 , \16139 , \16544 );
xor \U$16776 ( \17119 , \17118 , \16559 );
xor \U$16777 ( \17120 , \16646 , \16648 );
xor \U$16778 ( \17121 , \17120 , \17104 );
and \U$16779 ( \17122 , \17119 , \17121 );
xor \U$16780 ( \17123 , \16824 , \16831 );
xor \U$16781 ( \17124 , \17123 , \16839 );
xor \U$16782 ( \17125 , \16880 , \16887 );
xor \U$16783 ( \17126 , \17125 , \16895 );
and \U$16784 ( \17127 , \17124 , \17126 );
not \U$16785 ( \17128 , \16849 );
xor \U$16786 ( \17129 , \16867 , \16857 );
not \U$16787 ( \17130 , \17129 );
or \U$16788 ( \17131 , \17128 , \17130 );
or \U$16789 ( \17132 , \17129 , \16849 );
nand \U$16790 ( \17133 , \17131 , \17132 );
xor \U$16791 ( \17134 , \16880 , \16887 );
xor \U$16792 ( \17135 , \17134 , \16895 );
and \U$16793 ( \17136 , \17133 , \17135 );
and \U$16794 ( \17137 , \17124 , \17133 );
or \U$16795 ( \17138 , \17127 , \17136 , \17137 );
not \U$16796 ( \17139 , \386 );
and \U$16797 ( \17140 , \395 , RI9870330_83);
and \U$16798 ( \17141 , RI9870240_81, \393 );
nor \U$16799 ( \17142 , \17140 , \17141 );
not \U$16800 ( \17143 , \17142 );
or \U$16801 ( \17144 , \17139 , \17143 );
or \U$16802 ( \17145 , \17142 , \487 );
nand \U$16803 ( \17146 , \17144 , \17145 );
not \U$16804 ( \17147 , \454 );
and \U$16805 ( \17148 , \465 , RI98708d0_95);
and \U$16806 ( \17149 , RI98707e0_93, \463 );
nor \U$16807 ( \17150 , \17148 , \17149 );
not \U$16808 ( \17151 , \17150 );
or \U$16809 ( \17152 , \17147 , \17151 );
or \U$16810 ( \17153 , \17150 , \456 );
nand \U$16811 ( \17154 , \17152 , \17153 );
xor \U$16812 ( \17155 , \17146 , \17154 );
not \U$16813 ( \17156 , \365 );
and \U$16814 ( \17157 , \376 , RI98706f0_91);
and \U$16815 ( \17158 , RI9870600_89, \374 );
nor \U$16816 ( \17159 , \17157 , \17158 );
not \U$16817 ( \17160 , \17159 );
or \U$16818 ( \17161 , \17156 , \17160 );
or \U$16819 ( \17162 , \17159 , \367 );
nand \U$16820 ( \17163 , \17161 , \17162 );
and \U$16821 ( \17164 , \17155 , \17163 );
and \U$16822 ( \17165 , \17146 , \17154 );
or \U$16823 ( \17166 , \17164 , \17165 );
xor \U$16824 ( \17167 , \16966 , \16971 );
xor \U$16825 ( \17168 , \17167 , \16980 );
and \U$16826 ( \17169 , \17166 , \17168 );
xor \U$16827 ( \17170 , \16999 , \17007 );
xor \U$16828 ( \17171 , \17170 , \17016 );
xor \U$16829 ( \17172 , \16966 , \16971 );
xor \U$16830 ( \17173 , \17172 , \16980 );
and \U$16831 ( \17174 , \17171 , \17173 );
and \U$16832 ( \17175 , \17166 , \17171 );
or \U$16833 ( \17176 , \17169 , \17174 , \17175 );
xor \U$16834 ( \17177 , \17138 , \17176 );
not \U$16835 ( \17178 , \16682 );
xor \U$16836 ( \17179 , \16691 , \16702 );
not \U$16837 ( \17180 , \17179 );
or \U$16838 ( \17181 , \17178 , \17180 );
or \U$16839 ( \17182 , \17179 , \16682 );
nand \U$16840 ( \17183 , \17181 , \17182 );
not \U$16841 ( \17184 , \16712 );
xor \U$16842 ( \17185 , \16721 , \16731 );
not \U$16843 ( \17186 , \17185 );
or \U$16844 ( \17187 , \17184 , \17186 );
or \U$16845 ( \17188 , \17185 , \16712 );
nand \U$16846 ( \17189 , \17187 , \17188 );
xor \U$16847 ( \17190 , \17183 , \17189 );
xor \U$16848 ( \17191 , \16657 , \16664 );
xor \U$16849 ( \17192 , \17191 , \16672 );
and \U$16850 ( \17193 , \17190 , \17192 );
and \U$16851 ( \17194 , \17183 , \17189 );
or \U$16852 ( \17195 , \17193 , \17194 );
and \U$16853 ( \17196 , \17177 , \17195 );
and \U$16854 ( \17197 , \17138 , \17176 );
or \U$16855 ( \17198 , \17196 , \17197 );
and \U$16856 ( \17199 , \1329 , RI9870060_77);
and \U$16857 ( \17200 , RI9870150_79, \1327 );
nor \U$16858 ( \17201 , \17199 , \17200 );
and \U$16859 ( \17202 , \17201 , \1336 );
not \U$16860 ( \17203 , \17201 );
and \U$16861 ( \17204 , \17203 , \1337 );
nor \U$16862 ( \17205 , \17202 , \17204 );
and \U$16863 ( \17206 , \1311 , RI9870f60_109);
and \U$16864 ( \17207 , RI9870ab0_99, \1309 );
nor \U$16865 ( \17208 , \17206 , \17207 );
and \U$16866 ( \17209 , \17208 , \1458 );
not \U$16867 ( \17210 , \17208 );
and \U$16868 ( \17211 , \17210 , \1318 );
nor \U$16869 ( \17212 , \17209 , \17211 );
xor \U$16870 ( \17213 , \17205 , \17212 );
not \U$16871 ( \17214 , \1462 );
and \U$16872 ( \17215 , \2042 , RI9870d80_105);
and \U$16873 ( \17216 , RI98709c0_97, \2040 );
nor \U$16874 ( \17217 , \17215 , \17216 );
not \U$16875 ( \17218 , \17217 );
or \U$16876 ( \17219 , \17214 , \17218 );
or \U$16877 ( \17220 , \17217 , \2034 );
nand \U$16878 ( \17221 , \17219 , \17220 );
and \U$16879 ( \17222 , \17213 , \17221 );
and \U$16880 ( \17223 , \17205 , \17212 );
or \U$16881 ( \17224 , \17222 , \17223 );
not \U$16882 ( \17225 , \1128 );
and \U$16883 ( \17226 , \1293 , RI986ff70_75);
and \U$16884 ( \17227 , RI986fe80_73, \1291 );
nor \U$16885 ( \17228 , \17226 , \17227 );
not \U$16886 ( \17229 , \17228 );
or \U$16887 ( \17230 , \17225 , \17229 );
or \U$16888 ( \17231 , \17228 , \1128 );
nand \U$16889 ( \17232 , \17230 , \17231 );
and \U$16890 ( \17233 , \776 , RI986fd90_71);
and \U$16891 ( \17234 , RI986fca0_69, \774 );
nor \U$16892 ( \17235 , \17233 , \17234 );
and \U$16893 ( \17236 , \17235 , \474 );
not \U$16894 ( \17237 , \17235 );
and \U$16895 ( \17238 , \17237 , \451 );
nor \U$16896 ( \17239 , \17236 , \17238 );
xor \U$16897 ( \17240 , \17232 , \17239 );
and \U$16898 ( \17241 , \438 , RI986fac0_65);
and \U$16899 ( \17242 , RI986fbb0_67, \436 );
nor \U$16900 ( \17243 , \17241 , \17242 );
and \U$16901 ( \17244 , \17243 , \444 );
not \U$16902 ( \17245 , \17243 );
and \U$16903 ( \17246 , \17245 , \443 );
nor \U$16904 ( \17247 , \17244 , \17246 );
and \U$16905 ( \17248 , \17240 , \17247 );
and \U$16906 ( \17249 , \17232 , \17239 );
or \U$16907 ( \17250 , \17248 , \17249 );
xor \U$16908 ( \17251 , \17224 , \17250 );
not \U$16909 ( \17252 , \2935 );
and \U$16910 ( \17253 , \3254 , RI9871230_115);
and \U$16911 ( \17254 , RI9871140_113, \3252 );
nor \U$16912 ( \17255 , \17253 , \17254 );
not \U$16913 ( \17256 , \17255 );
or \U$16914 ( \17257 , \17252 , \17256 );
or \U$16915 ( \17258 , \17255 , \2935 );
nand \U$16916 ( \17259 , \17257 , \17258 );
and \U$16917 ( \17260 , \2274 , RI9870e70_107);
and \U$16918 ( \17261 , RI9870ba0_101, \2272 );
nor \U$16919 ( \17262 , \17260 , \17261 );
and \U$16920 ( \17263 , \17262 , \2030 );
not \U$16921 ( \17264 , \17262 );
and \U$16922 ( \17265 , \17264 , \2031 );
nor \U$16923 ( \17266 , \17263 , \17265 );
xor \U$16924 ( \17267 , \17259 , \17266 );
and \U$16925 ( \17268 , \2464 , RI9871050_111);
and \U$16926 ( \17269 , RI9870c90_103, \2462 );
nor \U$16927 ( \17270 , \17268 , \17269 );
and \U$16928 ( \17271 , \17270 , \2468 );
not \U$16929 ( \17272 , \17270 );
and \U$16930 ( \17273 , \17272 , \2263 );
nor \U$16931 ( \17274 , \17271 , \17273 );
and \U$16932 ( \17275 , \17267 , \17274 );
and \U$16933 ( \17276 , \17259 , \17266 );
or \U$16934 ( \17277 , \17275 , \17276 );
and \U$16935 ( \17278 , \17251 , \17277 );
and \U$16936 ( \17279 , \17224 , \17250 );
or \U$16937 ( \17280 , \17278 , \17279 );
and \U$16938 ( \17281 , \9237 , RI986e530_19);
and \U$16939 ( \17282 , RI986e440_17, \9235 );
nor \U$16940 ( \17283 , \17281 , \17282 );
and \U$16941 ( \17284 , \17283 , \9241 );
not \U$16942 ( \17285 , \17283 );
and \U$16943 ( \17286 , \17285 , \8836 );
nor \U$16944 ( \17287 , \17284 , \17286 );
and \U$16945 ( \17288 , \9505 , RI986e710_23);
and \U$16946 ( \17289 , RI986e620_21, \9503 );
nor \U$16947 ( \17290 , \17288 , \17289 );
and \U$16948 ( \17291 , \17290 , \9510 );
not \U$16949 ( \17292 , \17290 );
and \U$16950 ( \17293 , \17292 , \9513 );
nor \U$16951 ( \17294 , \17291 , \17293 );
xor \U$16952 ( \17295 , \17287 , \17294 );
and \U$16953 ( \17296 , \10424 , RI986f7f0_59);
and \U$16954 ( \17297 , RI986f700_57, \10422 );
nor \U$16955 ( \17298 , \17296 , \17297 );
and \U$16956 ( \17299 , \17298 , \9840 );
not \U$16957 ( \17300 , \17298 );
and \U$16958 ( \17301 , \17300 , \10428 );
nor \U$16959 ( \17302 , \17299 , \17301 );
and \U$16960 ( \17303 , \17295 , \17302 );
and \U$16961 ( \17304 , \17287 , \17294 );
or \U$16962 ( \17305 , \17303 , \17304 );
and \U$16963 ( \17306 , \13882 , RI986df90_7);
and \U$16964 ( \17307 , RI986dea0_5, \13880 );
nor \U$16965 ( \17308 , \17306 , \17307 );
and \U$16966 ( \17309 , \17308 , \13358 );
not \U$16967 ( \17310 , \17308 );
and \U$16968 ( \17311 , \17310 , \13359 );
nor \U$16969 ( \17312 , \17309 , \17311 );
not \U$16970 ( \17313 , RI9873558_190);
and \U$16971 ( \17314 , \15780 , RI986e170_11);
and \U$16972 ( \17315 , RI9873648_192, RI986e080_9);
nor \U$16973 ( \17316 , \17314 , \17315 );
not \U$16974 ( \17317 , \17316 );
or \U$16975 ( \17318 , \17313 , \17317 );
or \U$16976 ( \17319 , \17316 , RI9873558_190);
nand \U$16977 ( \17320 , \17318 , \17319 );
xor \U$16978 ( \17321 , \17312 , \17320 );
and \U$16979 ( \17322 , \14937 , RI986ddb0_3);
and \U$16980 ( \17323 , RI986dcc0_1, \14935 );
nor \U$16981 ( \17324 , \17322 , \17323 );
and \U$16982 ( \17325 , \17324 , \14539 );
not \U$16983 ( \17326 , \17324 );
and \U$16984 ( \17327 , \17326 , \14538 );
nor \U$16985 ( \17328 , \17325 , \17327 );
and \U$16986 ( \17329 , \17321 , \17328 );
and \U$16987 ( \17330 , \17312 , \17320 );
or \U$16988 ( \17331 , \17329 , \17330 );
xor \U$16989 ( \17332 , \17305 , \17331 );
and \U$16990 ( \17333 , \11696 , RI986f9d0_63);
and \U$16991 ( \17334 , RI986f8e0_61, \11694 );
nor \U$16992 ( \17335 , \17333 , \17334 );
and \U$16993 ( \17336 , \17335 , \10965 );
not \U$16994 ( \17337 , \17335 );
and \U$16995 ( \17338 , \17337 , \11702 );
nor \U$16996 ( \17339 , \17336 , \17338 );
and \U$16997 ( \17340 , \12293 , RI986f430_51);
and \U$16998 ( \17341 , RI986f340_49, \12291 );
nor \U$16999 ( \17342 , \17340 , \17341 );
and \U$17000 ( \17343 , \17342 , \11687 );
not \U$17001 ( \17344 , \17342 );
and \U$17002 ( \17345 , \17344 , \11686 );
nor \U$17003 ( \17346 , \17343 , \17345 );
xor \U$17004 ( \17347 , \17339 , \17346 );
and \U$17005 ( \17348 , \13045 , RI986f520_53);
and \U$17006 ( \17349 , RI986f610_55, \13043 );
nor \U$17007 ( \17350 , \17348 , \17349 );
and \U$17008 ( \17351 , \17350 , \13047 );
not \U$17009 ( \17352 , \17350 );
and \U$17010 ( \17353 , \17352 , \12619 );
nor \U$17011 ( \17354 , \17351 , \17353 );
and \U$17012 ( \17355 , \17347 , \17354 );
and \U$17013 ( \17356 , \17339 , \17346 );
or \U$17014 ( \17357 , \17355 , \17356 );
and \U$17015 ( \17358 , \17332 , \17357 );
and \U$17016 ( \17359 , \17305 , \17331 );
or \U$17017 ( \17360 , \17358 , \17359 );
xor \U$17018 ( \17361 , \17280 , \17360 );
and \U$17019 ( \17362 , \7079 , RI986ebc0_33);
and \U$17020 ( \17363 , RI986ecb0_35, \7077 );
nor \U$17021 ( \17364 , \17362 , \17363 );
and \U$17022 ( \17365 , \17364 , \6710 );
not \U$17023 ( \17366 , \17364 );
and \U$17024 ( \17367 , \17366 , \6709 );
nor \U$17025 ( \17368 , \17365 , \17367 );
and \U$17026 ( \17369 , \7729 , RI986f070_43);
and \U$17027 ( \17370 , RI986ef80_41, \7727 );
nor \U$17028 ( \17371 , \17369 , \17370 );
and \U$17029 ( \17372 , \17371 , \7480 );
not \U$17030 ( \17373 , \17371 );
and \U$17031 ( \17374 , \17373 , \7733 );
nor \U$17032 ( \17375 , \17372 , \17374 );
xor \U$17033 ( \17376 , \17368 , \17375 );
and \U$17034 ( \17377 , \8486 , RI986f250_47);
and \U$17035 ( \17378 , RI986f160_45, \8484 );
nor \U$17036 ( \17379 , \17377 , \17378 );
and \U$17037 ( \17380 , \17379 , \8050 );
not \U$17038 ( \17381 , \17379 );
and \U$17039 ( \17382 , \17381 , \8051 );
nor \U$17040 ( \17383 , \17380 , \17382 );
and \U$17041 ( \17384 , \17376 , \17383 );
and \U$17042 ( \17385 , \17368 , \17375 );
or \U$17043 ( \17386 , \17384 , \17385 );
and \U$17044 ( \17387 , \5318 , RI986ead0_31);
and \U$17045 ( \17388 , RI986e9e0_29, \5316 );
nor \U$17046 ( \17389 , \17387 , \17388 );
and \U$17047 ( \17390 , \17389 , \5052 );
not \U$17048 ( \17391 , \17389 );
and \U$17049 ( \17392 , \17391 , \5322 );
nor \U$17050 ( \17393 , \17390 , \17392 );
and \U$17051 ( \17394 , \5881 , RI986e8f0_27);
and \U$17052 ( \17395 , RI986e800_25, \5879 );
nor \U$17053 ( \17396 , \17394 , \17395 );
and \U$17054 ( \17397 , \17396 , \5594 );
not \U$17055 ( \17398 , \17396 );
and \U$17056 ( \17399 , \17398 , \5885 );
nor \U$17057 ( \17400 , \17397 , \17399 );
xor \U$17058 ( \17401 , \17393 , \17400 );
and \U$17059 ( \17402 , \6453 , RI986ee90_39);
and \U$17060 ( \17403 , RI986eda0_37, \6451 );
nor \U$17061 ( \17404 , \17402 , \17403 );
and \U$17062 ( \17405 , \17404 , \6190 );
not \U$17063 ( \17406 , \17404 );
and \U$17064 ( \17407 , \17406 , \6180 );
nor \U$17065 ( \17408 , \17405 , \17407 );
and \U$17066 ( \17409 , \17401 , \17408 );
and \U$17067 ( \17410 , \17393 , \17400 );
or \U$17068 ( \17411 , \17409 , \17410 );
xor \U$17069 ( \17412 , \17386 , \17411 );
not \U$17070 ( \17413 , \4521 );
and \U$17071 ( \17414 , \4710 , RI9871500_121);
and \U$17072 ( \17415 , RI98715f0_123, \4708 );
nor \U$17073 ( \17416 , \17414 , \17415 );
not \U$17074 ( \17417 , \17416 );
or \U$17075 ( \17418 , \17413 , \17417 );
or \U$17076 ( \17419 , \17416 , \4519 );
nand \U$17077 ( \17420 , \17418 , \17419 );
not \U$17078 ( \17421 , \3412 );
and \U$17079 ( \17422 , \3683 , RI9871320_117);
and \U$17080 ( \17423 , RI9871410_119, \3681 );
nor \U$17081 ( \17424 , \17422 , \17423 );
not \U$17082 ( \17425 , \17424 );
or \U$17083 ( \17426 , \17421 , \17425 );
or \U$17084 ( \17427 , \17424 , \3412 );
nand \U$17085 ( \17428 , \17426 , \17427 );
xor \U$17086 ( \17429 , \17420 , \17428 );
and \U$17087 ( \17430 , \4203 , RI98716e0_125);
and \U$17088 ( \17431 , RI98717d0_127, \4201 );
nor \U$17089 ( \17432 , \17430 , \17431 );
and \U$17090 ( \17433 , \17432 , \4207 );
not \U$17091 ( \17434 , \17432 );
and \U$17092 ( \17435 , \17434 , \3922 );
nor \U$17093 ( \17436 , \17433 , \17435 );
and \U$17094 ( \17437 , \17429 , \17436 );
and \U$17095 ( \17438 , \17420 , \17428 );
or \U$17096 ( \17439 , \17437 , \17438 );
and \U$17097 ( \17440 , \17412 , \17439 );
and \U$17098 ( \17441 , \17386 , \17411 );
or \U$17099 ( \17442 , \17440 , \17441 );
and \U$17100 ( \17443 , \17361 , \17442 );
and \U$17101 ( \17444 , \17280 , \17360 );
or \U$17102 ( \17445 , \17443 , \17444 );
xor \U$17103 ( \17446 , \17198 , \17445 );
not \U$17104 ( \17447 , \421 );
xnor \U$17105 ( \17448 , \16755 , \16744 );
not \U$17106 ( \17449 , \17448 );
or \U$17107 ( \17450 , \17447 , \17449 );
or \U$17108 ( \17451 , \17448 , \421 );
nand \U$17109 ( \17452 , \17450 , \17451 );
not \U$17110 ( \17453 , \16764 );
xor \U$17111 ( \17454 , \16772 , \16782 );
not \U$17112 ( \17455 , \17454 );
or \U$17113 ( \17456 , \17453 , \17455 );
or \U$17114 ( \17457 , \17454 , \16764 );
nand \U$17115 ( \17458 , \17456 , \17457 );
xor \U$17116 ( \17459 , \17452 , \17458 );
not \U$17117 ( \17460 , \16792 );
xor \U$17118 ( \17461 , \16800 , \16810 );
not \U$17119 ( \17462 , \17461 );
or \U$17120 ( \17463 , \17460 , \17462 );
or \U$17121 ( \17464 , \17461 , \16792 );
nand \U$17122 ( \17465 , \17463 , \17464 );
and \U$17123 ( \17466 , \17459 , \17465 );
and \U$17124 ( \17467 , \17452 , \17458 );
or \U$17125 ( \17468 , \17466 , \17467 );
not \U$17126 ( \17469 , \16909 );
not \U$17127 ( \17470 , \16906 );
or \U$17128 ( \17471 , \17469 , \17470 );
or \U$17129 ( \17472 , \16906 , \16909 );
nand \U$17130 ( \17473 , \17471 , \17472 );
xor \U$17131 ( \17474 , \17468 , \17473 );
xor \U$17132 ( \17475 , \16318 , \16325 );
xor \U$17133 ( \17476 , \17475 , \16333 );
xor \U$17134 ( \17477 , \16918 , \16923 );
xor \U$17135 ( \17478 , \17476 , \17477 );
and \U$17136 ( \17479 , \17474 , \17478 );
and \U$17137 ( \17480 , \17468 , \17473 );
or \U$17138 ( \17481 , \17479 , \17480 );
and \U$17139 ( \17482 , \17446 , \17481 );
and \U$17140 ( \17483 , \17198 , \17445 );
nor \U$17141 ( \17484 , \17482 , \17483 );
xor \U$17142 ( \17485 , \16675 , \16704 );
xor \U$17143 ( \17486 , \17485 , \16733 );
not \U$17144 ( \17487 , \17486 );
not \U$17145 ( \17488 , \16898 );
not \U$17146 ( \17489 , \16869 );
or \U$17147 ( \17490 , \17488 , \17489 );
or \U$17148 ( \17491 , \16869 , \16898 );
nand \U$17149 ( \17492 , \17490 , \17491 );
not \U$17150 ( \17493 , \17492 );
not \U$17151 ( \17494 , \16842 );
and \U$17152 ( \17495 , \17493 , \17494 );
and \U$17153 ( \17496 , \17492 , \16842 );
nor \U$17154 ( \17497 , \17495 , \17496 );
not \U$17155 ( \17498 , \17497 );
and \U$17156 ( \17499 , \17487 , \17498 );
and \U$17157 ( \17500 , \17497 , \17486 );
xor \U$17158 ( \17501 , \16757 , \16784 );
xor \U$17159 ( \17502 , \17501 , \16812 );
nor \U$17160 ( \17503 , \17500 , \17502 );
nor \U$17161 ( \17504 , \17499 , \17503 );
not \U$17162 ( \17505 , \17504 );
xor \U$17163 ( \17506 , \16164 , \16190 );
xor \U$17164 ( \17507 , \17506 , \16216 );
not \U$17165 ( \17508 , \17507 );
and \U$17166 ( \17509 , \17505 , \17508 );
and \U$17167 ( \17510 , \17504 , \17507 );
xor \U$17168 ( \17511 , \16983 , \16991 );
xor \U$17169 ( \17512 , \17511 , \17019 );
xor \U$17170 ( \17513 , \16941 , \16948 );
xor \U$17171 ( \17514 , \17513 , \16955 );
and \U$17172 ( \17515 , \17512 , \17514 );
xor \U$17173 ( \17516 , \16370 , \16378 );
xor \U$17174 ( \17517 , \17516 , \16386 );
xor \U$17175 ( \17518 , \17029 , \17038 );
xor \U$17176 ( \17519 , \17517 , \17518 );
xor \U$17177 ( \17520 , \16941 , \16948 );
xor \U$17178 ( \17521 , \17520 , \16955 );
and \U$17179 ( \17522 , \17519 , \17521 );
and \U$17180 ( \17523 , \17512 , \17519 );
or \U$17181 ( \17524 , \17515 , \17522 , \17523 );
not \U$17182 ( \17525 , \17524 );
nor \U$17183 ( \17526 , \17510 , \17525 );
nor \U$17184 ( \17527 , \17509 , \17526 );
xor \U$17185 ( \17528 , \17484 , \17527 );
not \U$17186 ( \17529 , \17056 );
not \U$17187 ( \17530 , \17064 );
or \U$17188 ( \17531 , \17529 , \17530 );
or \U$17189 ( \17532 , \17056 , \17064 );
nand \U$17190 ( \17533 , \17531 , \17532 );
not \U$17191 ( \17534 , \17533 );
not \U$17192 ( \17535 , \17058 );
and \U$17193 ( \17536 , \17534 , \17535 );
and \U$17194 ( \17537 , \17533 , \17058 );
nor \U$17195 ( \17538 , \17536 , \17537 );
not \U$17196 ( \17539 , \17538 );
xor \U$17197 ( \17540 , \16910 , \16915 );
xor \U$17198 ( \17541 , \17540 , \16929 );
not \U$17199 ( \17542 , \17541 );
and \U$17200 ( \17543 , \17539 , \17542 );
and \U$17201 ( \17544 , \17538 , \17541 );
xor \U$17202 ( \17545 , \17069 , \17071 );
xor \U$17203 ( \17546 , \17545 , \17074 );
nor \U$17204 ( \17547 , \17544 , \17546 );
nor \U$17205 ( \17548 , \17543 , \17547 );
and \U$17206 ( \17549 , \17528 , \17548 );
and \U$17207 ( \17550 , \17484 , \17527 );
or \U$17208 ( \17551 , \17549 , \17550 );
not \U$17209 ( \17552 , \16137 );
not \U$17210 ( \17553 , \16117 );
or \U$17211 ( \17554 , \17552 , \17553 );
or \U$17212 ( \17555 , \16117 , \16137 );
nand \U$17213 ( \17556 , \17554 , \17555 );
not \U$17214 ( \17557 , \17556 );
not \U$17215 ( \17558 , \16119 );
and \U$17216 ( \17559 , \17557 , \17558 );
and \U$17217 ( \17560 , \17556 , \16119 );
nor \U$17218 ( \17561 , \17559 , \17560 );
or \U$17219 ( \17562 , \17551 , \17561 );
not \U$17220 ( \17563 , \17561 );
not \U$17221 ( \17564 , \17551 );
or \U$17222 ( \17565 , \17563 , \17564 );
xor \U$17223 ( \17566 , \17054 , \17066 );
xor \U$17224 ( \17567 , \17566 , \17077 );
not \U$17225 ( \17568 , \16308 );
xor \U$17226 ( \17569 , \16219 , \16392 );
not \U$17227 ( \17570 , \17569 );
or \U$17228 ( \17571 , \17568 , \17570 );
or \U$17229 ( \17572 , \17569 , \16308 );
nand \U$17230 ( \17573 , \17571 , \17572 );
xor \U$17231 ( \17574 , \17567 , \17573 );
not \U$17232 ( \17575 , \17083 );
xor \U$17233 ( \17576 , \17086 , \17099 );
not \U$17234 ( \17577 , \17576 );
or \U$17235 ( \17578 , \17575 , \17577 );
or \U$17236 ( \17579 , \17576 , \17083 );
nand \U$17237 ( \17580 , \17578 , \17579 );
and \U$17238 ( \17581 , \17574 , \17580 );
and \U$17239 ( \17582 , \17567 , \17573 );
or \U$17240 ( \17583 , \17581 , \17582 );
nand \U$17241 ( \17584 , \17565 , \17583 );
nand \U$17242 ( \17585 , \17562 , \17584 );
xor \U$17243 ( \17586 , \15638 , \15648 );
xor \U$17244 ( \17587 , \17586 , \15653 );
xor \U$17245 ( \17588 , \16567 , \16574 );
xor \U$17246 ( \17589 , \17587 , \17588 );
xor \U$17247 ( \17590 , \17585 , \17589 );
xor \U$17248 ( \17591 , \17048 , \17080 );
xor \U$17249 ( \17592 , \17591 , \17101 );
xor \U$17250 ( \17593 , \16394 , \16503 );
xor \U$17251 ( \17594 , \17593 , \16541 );
or \U$17252 ( \17595 , \17592 , \17594 );
not \U$17253 ( \17596 , \17594 );
not \U$17254 ( \17597 , \17592 );
or \U$17255 ( \17598 , \17596 , \17597 );
xor \U$17256 ( \17599 , \15959 , \16019 );
xor \U$17257 ( \17600 , \17599 , \16054 );
xor \U$17258 ( \17601 , \16634 , \16641 );
xor \U$17259 ( \17602 , \17600 , \17601 );
nand \U$17260 ( \17603 , \17598 , \17602 );
nand \U$17261 ( \17604 , \17595 , \17603 );
and \U$17262 ( \17605 , \17590 , \17604 );
and \U$17263 ( \17606 , \17585 , \17589 );
or \U$17264 ( \17607 , \17605 , \17606 );
xor \U$17265 ( \17608 , \17122 , \17607 );
not \U$17266 ( \17609 , \17608 );
or \U$17267 ( \17610 , \17117 , \17609 );
or \U$17268 ( \17611 , \17608 , \17116 );
nand \U$17269 ( \17612 , \17610 , \17611 );
xor \U$17270 ( \17613 , \17119 , \17121 );
not \U$17271 ( \17614 , \17613 );
xor \U$17272 ( \17615 , \17585 , \17589 );
xor \U$17273 ( \17616 , \17615 , \17604 );
not \U$17274 ( \17617 , \17616 );
or \U$17275 ( \17618 , \17614 , \17617 );
or \U$17276 ( \17619 , \17616 , \17613 );
not \U$17277 ( \17620 , \17551 );
not \U$17278 ( \17621 , \17583 );
or \U$17279 ( \17622 , \17620 , \17621 );
or \U$17280 ( \17623 , \17583 , \17551 );
nand \U$17281 ( \17624 , \17622 , \17623 );
not \U$17282 ( \17625 , \17624 );
not \U$17283 ( \17626 , \17561 );
and \U$17284 ( \17627 , \17625 , \17626 );
and \U$17285 ( \17628 , \17624 , \17561 );
nor \U$17286 ( \17629 , \17627 , \17628 );
xnor \U$17287 ( \17630 , \17594 , \17592 );
not \U$17288 ( \17631 , \17630 );
not \U$17289 ( \17632 , \17602 );
and \U$17290 ( \17633 , \17631 , \17632 );
and \U$17291 ( \17634 , \17630 , \17602 );
nor \U$17292 ( \17635 , \17633 , \17634 );
or \U$17293 ( \17636 , \17629 , \17635 );
not \U$17294 ( \17637 , \17635 );
not \U$17295 ( \17638 , \17629 );
or \U$17296 ( \17639 , \17637 , \17638 );
xor \U$17297 ( \17640 , \16958 , \17022 );
xor \U$17298 ( \17641 , \17640 , \17043 );
xor \U$17299 ( \17642 , \16736 , \16815 );
xor \U$17300 ( \17643 , \17642 , \16900 );
xor \U$17301 ( \17644 , \17641 , \17643 );
not \U$17302 ( \17645 , \17541 );
xor \U$17303 ( \17646 , \17538 , \17546 );
not \U$17304 ( \17647 , \17646 );
or \U$17305 ( \17648 , \17645 , \17647 );
or \U$17306 ( \17649 , \17646 , \17541 );
nand \U$17307 ( \17650 , \17648 , \17649 );
and \U$17308 ( \17651 , \17644 , \17650 );
and \U$17309 ( \17652 , \17641 , \17643 );
or \U$17310 ( \17653 , \17651 , \17652 );
not \U$17311 ( \17654 , \16932 );
xor \U$17312 ( \17655 , \16903 , \17046 );
not \U$17313 ( \17656 , \17655 );
or \U$17314 ( \17657 , \17654 , \17656 );
or \U$17315 ( \17658 , \17655 , \16932 );
nand \U$17316 ( \17659 , \17657 , \17658 );
xor \U$17317 ( \17660 , \17653 , \17659 );
xor \U$17318 ( \17661 , \17138 , \17176 );
xor \U$17319 ( \17662 , \17661 , \17195 );
xor \U$17320 ( \17663 , \17280 , \17360 );
xor \U$17321 ( \17664 , \17663 , \17442 );
xor \U$17322 ( \17665 , \17662 , \17664 );
xor \U$17323 ( \17666 , \17468 , \17473 );
xor \U$17324 ( \17667 , \17666 , \17478 );
and \U$17325 ( \17668 , \17665 , \17667 );
and \U$17326 ( \17669 , \17662 , \17664 );
or \U$17327 ( \17670 , \17668 , \17669 );
xor \U$17328 ( \17671 , \17205 , \17212 );
xor \U$17329 ( \17672 , \17671 , \17221 );
xor \U$17330 ( \17673 , \17146 , \17154 );
xor \U$17331 ( \17674 , \17673 , \17163 );
xor \U$17332 ( \17675 , \17672 , \17674 );
xor \U$17333 ( \17676 , \17232 , \17239 );
xor \U$17334 ( \17677 , \17676 , \17247 );
and \U$17335 ( \17678 , \17675 , \17677 );
and \U$17336 ( \17679 , \17672 , \17674 );
or \U$17337 ( \17680 , \17678 , \17679 );
nand \U$17338 ( \17681 , RI9870420_85, \352 );
not \U$17339 ( \17682 , \17681 );
not \U$17340 ( \17683 , \345 );
or \U$17341 ( \17684 , \17682 , \17683 );
or \U$17342 ( \17685 , \345 , \17681 );
nand \U$17343 ( \17686 , \17684 , \17685 );
not \U$17344 ( \17687 , \487 );
and \U$17345 ( \17688 , \395 , RI9870510_87);
and \U$17346 ( \17689 , RI9870330_83, \393 );
nor \U$17347 ( \17690 , \17688 , \17689 );
not \U$17348 ( \17691 , \17690 );
or \U$17349 ( \17692 , \17687 , \17691 );
or \U$17350 ( \17693 , \17690 , \386 );
nand \U$17351 ( \17694 , \17692 , \17693 );
and \U$17352 ( \17695 , \17686 , \17694 );
not \U$17353 ( \17696 , \345 );
and \U$17354 ( \17697 , \354 , RI9870420_85);
and \U$17355 ( \17698 , RI9870510_87, \352 );
nor \U$17356 ( \17699 , \17697 , \17698 );
not \U$17357 ( \17700 , \17699 );
or \U$17358 ( \17701 , \17696 , \17700 );
or \U$17359 ( \17702 , \17699 , \345 );
nand \U$17360 ( \17703 , \17701 , \17702 );
xor \U$17361 ( \17704 , \17695 , \17703 );
and \U$17362 ( \17705 , \438 , RI98707e0_93);
and \U$17363 ( \17706 , RI986fac0_65, \436 );
nor \U$17364 ( \17707 , \17705 , \17706 );
and \U$17365 ( \17708 , \17707 , \444 );
not \U$17366 ( \17709 , \17707 );
and \U$17367 ( \17710 , \17709 , \443 );
nor \U$17368 ( \17711 , \17708 , \17710 );
not \U$17369 ( \17712 , \454 );
and \U$17370 ( \17713 , \465 , RI9870600_89);
and \U$17371 ( \17714 , RI98708d0_95, \463 );
nor \U$17372 ( \17715 , \17713 , \17714 );
not \U$17373 ( \17716 , \17715 );
or \U$17374 ( \17717 , \17712 , \17716 );
or \U$17375 ( \17718 , \17715 , \456 );
nand \U$17376 ( \17719 , \17717 , \17718 );
xor \U$17377 ( \17720 , \17711 , \17719 );
not \U$17378 ( \17721 , \367 );
and \U$17379 ( \17722 , \376 , RI9870240_81);
and \U$17380 ( \17723 , RI98706f0_91, \374 );
nor \U$17381 ( \17724 , \17722 , \17723 );
not \U$17382 ( \17725 , \17724 );
or \U$17383 ( \17726 , \17721 , \17725 );
or \U$17384 ( \17727 , \17724 , \367 );
nand \U$17385 ( \17728 , \17726 , \17727 );
and \U$17386 ( \17729 , \17720 , \17728 );
and \U$17387 ( \17730 , \17711 , \17719 );
or \U$17388 ( \17731 , \17729 , \17730 );
and \U$17389 ( \17732 , \17704 , \17731 );
and \U$17390 ( \17733 , \17695 , \17703 );
or \U$17391 ( \17734 , \17732 , \17733 );
xor \U$17392 ( \17735 , \17680 , \17734 );
xor \U$17393 ( \17736 , \17259 , \17266 );
xor \U$17394 ( \17737 , \17736 , \17274 );
xor \U$17395 ( \17738 , \17393 , \17400 );
xor \U$17396 ( \17739 , \17738 , \17408 );
and \U$17397 ( \17740 , \17737 , \17739 );
xor \U$17398 ( \17741 , \17420 , \17428 );
xor \U$17399 ( \17742 , \17741 , \17436 );
xor \U$17400 ( \17743 , \17393 , \17400 );
xor \U$17401 ( \17744 , \17743 , \17408 );
and \U$17402 ( \17745 , \17742 , \17744 );
and \U$17403 ( \17746 , \17737 , \17742 );
or \U$17404 ( \17747 , \17740 , \17745 , \17746 );
and \U$17405 ( \17748 , \17735 , \17747 );
and \U$17406 ( \17749 , \17680 , \17734 );
or \U$17407 ( \17750 , \17748 , \17749 );
and \U$17408 ( \17751 , \2464 , RI9870ba0_101);
and \U$17409 ( \17752 , RI9871050_111, \2462 );
nor \U$17410 ( \17753 , \17751 , \17752 );
and \U$17411 ( \17754 , \17753 , \2468 );
not \U$17412 ( \17755 , \17753 );
and \U$17413 ( \17756 , \17755 , \2263 );
nor \U$17414 ( \17757 , \17754 , \17756 );
not \U$17415 ( \17758 , \3406 );
and \U$17416 ( \17759 , \3254 , RI9870c90_103);
and \U$17417 ( \17760 , RI9871230_115, \3252 );
nor \U$17418 ( \17761 , \17759 , \17760 );
not \U$17419 ( \17762 , \17761 );
or \U$17420 ( \17763 , \17758 , \17762 );
or \U$17421 ( \17764 , \17761 , \3406 );
nand \U$17422 ( \17765 , \17763 , \17764 );
xor \U$17423 ( \17766 , \17757 , \17765 );
not \U$17424 ( \17767 , \3412 );
and \U$17425 ( \17768 , \3683 , RI9871140_113);
and \U$17426 ( \17769 , RI9871320_117, \3681 );
nor \U$17427 ( \17770 , \17768 , \17769 );
not \U$17428 ( \17771 , \17770 );
or \U$17429 ( \17772 , \17767 , \17771 );
or \U$17430 ( \17773 , \17770 , \3412 );
nand \U$17431 ( \17774 , \17772 , \17773 );
and \U$17432 ( \17775 , \17766 , \17774 );
and \U$17433 ( \17776 , \17757 , \17765 );
or \U$17434 ( \17777 , \17775 , \17776 );
and \U$17435 ( \17778 , \776 , RI986fbb0_67);
and \U$17436 ( \17779 , RI986fd90_71, \774 );
nor \U$17437 ( \17780 , \17778 , \17779 );
and \U$17438 ( \17781 , \17780 , \474 );
not \U$17439 ( \17782 , \17780 );
and \U$17440 ( \17783 , \17782 , \451 );
nor \U$17441 ( \17784 , \17781 , \17783 );
not \U$17442 ( \17785 , \1301 );
and \U$17443 ( \17786 , \1293 , RI986fca0_69);
and \U$17444 ( \17787 , RI986ff70_75, \1291 );
nor \U$17445 ( \17788 , \17786 , \17787 );
not \U$17446 ( \17789 , \17788 );
or \U$17447 ( \17790 , \17785 , \17789 );
or \U$17448 ( \17791 , \17788 , \1128 );
nand \U$17449 ( \17792 , \17790 , \17791 );
xor \U$17450 ( \17793 , \17784 , \17792 );
and \U$17451 ( \17794 , \1329 , RI986fe80_73);
and \U$17452 ( \17795 , RI9870060_77, \1327 );
nor \U$17453 ( \17796 , \17794 , \17795 );
and \U$17454 ( \17797 , \17796 , \1336 );
not \U$17455 ( \17798 , \17796 );
and \U$17456 ( \17799 , \17798 , \1337 );
nor \U$17457 ( \17800 , \17797 , \17799 );
and \U$17458 ( \17801 , \17793 , \17800 );
and \U$17459 ( \17802 , \17784 , \17792 );
or \U$17460 ( \17803 , \17801 , \17802 );
xor \U$17461 ( \17804 , \17777 , \17803 );
and \U$17462 ( \17805 , \1311 , RI9870150_79);
and \U$17463 ( \17806 , RI9870f60_109, \1309 );
nor \U$17464 ( \17807 , \17805 , \17806 );
and \U$17465 ( \17808 , \17807 , \1458 );
not \U$17466 ( \17809 , \17807 );
and \U$17467 ( \17810 , \17809 , \1318 );
nor \U$17468 ( \17811 , \17808 , \17810 );
not \U$17469 ( \17812 , \1462 );
and \U$17470 ( \17813 , \2042 , RI9870ab0_99);
and \U$17471 ( \17814 , RI9870d80_105, \2040 );
nor \U$17472 ( \17815 , \17813 , \17814 );
not \U$17473 ( \17816 , \17815 );
or \U$17474 ( \17817 , \17812 , \17816 );
or \U$17475 ( \17818 , \17815 , \1462 );
nand \U$17476 ( \17819 , \17817 , \17818 );
xor \U$17477 ( \17820 , \17811 , \17819 );
and \U$17478 ( \17821 , \2274 , RI98709c0_97);
and \U$17479 ( \17822 , RI9870e70_107, \2272 );
nor \U$17480 ( \17823 , \17821 , \17822 );
and \U$17481 ( \17824 , \17823 , \2030 );
not \U$17482 ( \17825 , \17823 );
and \U$17483 ( \17826 , \17825 , \2031 );
nor \U$17484 ( \17827 , \17824 , \17826 );
and \U$17485 ( \17828 , \17820 , \17827 );
and \U$17486 ( \17829 , \17811 , \17819 );
or \U$17487 ( \17830 , \17828 , \17829 );
and \U$17488 ( \17831 , \17804 , \17830 );
and \U$17489 ( \17832 , \17777 , \17803 );
or \U$17490 ( \17833 , \17831 , \17832 );
and \U$17491 ( \17834 , \12293 , RI986f8e0_61);
and \U$17492 ( \17835 , RI986f430_51, \12291 );
nor \U$17493 ( \17836 , \17834 , \17835 );
and \U$17494 ( \17837 , \17836 , \11687 );
not \U$17495 ( \17838 , \17836 );
and \U$17496 ( \17839 , \17838 , \11686 );
nor \U$17497 ( \17840 , \17837 , \17839 );
and \U$17498 ( \17841 , \13045 , RI986f340_49);
and \U$17499 ( \17842 , RI986f520_53, \13043 );
nor \U$17500 ( \17843 , \17841 , \17842 );
and \U$17501 ( \17844 , \17843 , \13047 );
not \U$17502 ( \17845 , \17843 );
and \U$17503 ( \17846 , \17845 , \12619 );
nor \U$17504 ( \17847 , \17844 , \17846 );
xor \U$17505 ( \17848 , \17840 , \17847 );
and \U$17506 ( \17849 , \13882 , RI986f610_55);
and \U$17507 ( \17850 , RI986df90_7, \13880 );
nor \U$17508 ( \17851 , \17849 , \17850 );
and \U$17509 ( \17852 , \17851 , \13358 );
not \U$17510 ( \17853 , \17851 );
and \U$17511 ( \17854 , \17853 , \13359 );
nor \U$17512 ( \17855 , \17852 , \17854 );
and \U$17513 ( \17856 , \17848 , \17855 );
and \U$17514 ( \17857 , \17840 , \17847 );
or \U$17515 ( \17858 , \17856 , \17857 );
not \U$17516 ( \17859 , RI9873558_190);
and \U$17517 ( \17860 , \15780 , RI986dcc0_1);
and \U$17518 ( \17861 , RI9873648_192, RI986e170_11);
nor \U$17519 ( \17862 , \17860 , \17861 );
not \U$17520 ( \17863 , \17862 );
or \U$17521 ( \17864 , \17859 , \17863 );
or \U$17522 ( \17865 , \17862 , RI9873558_190);
nand \U$17523 ( \17866 , \17864 , \17865 );
xor \U$17524 ( \17867 , \17866 , \361 );
and \U$17525 ( \17868 , \14937 , RI986dea0_5);
and \U$17526 ( \17869 , RI986ddb0_3, \14935 );
nor \U$17527 ( \17870 , \17868 , \17869 );
and \U$17528 ( \17871 , \17870 , \14539 );
not \U$17529 ( \17872 , \17870 );
and \U$17530 ( \17873 , \17872 , \14538 );
nor \U$17531 ( \17874 , \17871 , \17873 );
and \U$17532 ( \17875 , \17867 , \17874 );
and \U$17533 ( \17876 , \17866 , \361 );
or \U$17534 ( \17877 , \17875 , \17876 );
xor \U$17535 ( \17878 , \17858 , \17877 );
and \U$17536 ( \17879 , \9505 , RI986e440_17);
and \U$17537 ( \17880 , RI986e710_23, \9503 );
nor \U$17538 ( \17881 , \17879 , \17880 );
and \U$17539 ( \17882 , \17881 , \9510 );
not \U$17540 ( \17883 , \17881 );
and \U$17541 ( \17884 , \17883 , \9513 );
nor \U$17542 ( \17885 , \17882 , \17884 );
and \U$17543 ( \17886 , \10424 , RI986e620_21);
and \U$17544 ( \17887 , RI986f7f0_59, \10422 );
nor \U$17545 ( \17888 , \17886 , \17887 );
and \U$17546 ( \17889 , \17888 , \9840 );
not \U$17547 ( \17890 , \17888 );
and \U$17548 ( \17891 , \17890 , \10428 );
nor \U$17549 ( \17892 , \17889 , \17891 );
xor \U$17550 ( \17893 , \17885 , \17892 );
and \U$17551 ( \17894 , \11696 , RI986f700_57);
and \U$17552 ( \17895 , RI986f9d0_63, \11694 );
nor \U$17553 ( \17896 , \17894 , \17895 );
and \U$17554 ( \17897 , \17896 , \10965 );
not \U$17555 ( \17898 , \17896 );
and \U$17556 ( \17899 , \17898 , \11702 );
nor \U$17557 ( \17900 , \17897 , \17899 );
and \U$17558 ( \17901 , \17893 , \17900 );
and \U$17559 ( \17902 , \17885 , \17892 );
or \U$17560 ( \17903 , \17901 , \17902 );
and \U$17561 ( \17904 , \17878 , \17903 );
and \U$17562 ( \17905 , \17858 , \17877 );
or \U$17563 ( \17906 , \17904 , \17905 );
xor \U$17564 ( \17907 , \17833 , \17906 );
and \U$17565 ( \17908 , \7729 , RI986ecb0_35);
and \U$17566 ( \17909 , RI986f070_43, \7727 );
nor \U$17567 ( \17910 , \17908 , \17909 );
and \U$17568 ( \17911 , \17910 , \7480 );
not \U$17569 ( \17912 , \17910 );
and \U$17570 ( \17913 , \17912 , \7733 );
nor \U$17571 ( \17914 , \17911 , \17913 );
and \U$17572 ( \17915 , \8486 , RI986ef80_41);
and \U$17573 ( \17916 , RI986f250_47, \8484 );
nor \U$17574 ( \17917 , \17915 , \17916 );
and \U$17575 ( \17918 , \17917 , \8050 );
not \U$17576 ( \17919 , \17917 );
and \U$17577 ( \17920 , \17919 , \8051 );
nor \U$17578 ( \17921 , \17918 , \17920 );
xor \U$17579 ( \17922 , \17914 , \17921 );
and \U$17580 ( \17923 , \9237 , RI986f160_45);
and \U$17581 ( \17924 , RI986e530_19, \9235 );
nor \U$17582 ( \17925 , \17923 , \17924 );
and \U$17583 ( \17926 , \17925 , \9241 );
not \U$17584 ( \17927 , \17925 );
and \U$17585 ( \17928 , \17927 , \8836 );
nor \U$17586 ( \17929 , \17926 , \17928 );
and \U$17587 ( \17930 , \17922 , \17929 );
and \U$17588 ( \17931 , \17914 , \17921 );
or \U$17589 ( \17932 , \17930 , \17931 );
and \U$17590 ( \17933 , \5881 , RI986e9e0_29);
and \U$17591 ( \17934 , RI986e8f0_27, \5879 );
nor \U$17592 ( \17935 , \17933 , \17934 );
and \U$17593 ( \17936 , \17935 , \5594 );
not \U$17594 ( \17937 , \17935 );
and \U$17595 ( \17938 , \17937 , \5885 );
nor \U$17596 ( \17939 , \17936 , \17938 );
and \U$17597 ( \17940 , \6453 , RI986e800_25);
and \U$17598 ( \17941 , RI986ee90_39, \6451 );
nor \U$17599 ( \17942 , \17940 , \17941 );
and \U$17600 ( \17943 , \17942 , \6190 );
not \U$17601 ( \17944 , \17942 );
and \U$17602 ( \17945 , \17944 , \6705 );
nor \U$17603 ( \17946 , \17943 , \17945 );
xor \U$17604 ( \17947 , \17939 , \17946 );
and \U$17605 ( \17948 , \7079 , RI986eda0_37);
and \U$17606 ( \17949 , RI986ebc0_33, \7077 );
nor \U$17607 ( \17950 , \17948 , \17949 );
and \U$17608 ( \17951 , \17950 , \6710 );
not \U$17609 ( \17952 , \17950 );
and \U$17610 ( \17953 , \17952 , \6709 );
nor \U$17611 ( \17954 , \17951 , \17953 );
and \U$17612 ( \17955 , \17947 , \17954 );
and \U$17613 ( \17956 , \17939 , \17946 );
or \U$17614 ( \17957 , \17955 , \17956 );
xor \U$17615 ( \17958 , \17932 , \17957 );
and \U$17616 ( \17959 , \4203 , RI9871410_119);
and \U$17617 ( \17960 , RI98716e0_125, \4201 );
nor \U$17618 ( \17961 , \17959 , \17960 );
and \U$17619 ( \17962 , \17961 , \4207 );
not \U$17620 ( \17963 , \17961 );
and \U$17621 ( \17964 , \17963 , \3922 );
nor \U$17622 ( \17965 , \17962 , \17964 );
not \U$17623 ( \17966 , \4521 );
and \U$17624 ( \17967 , \4710 , RI98717d0_127);
and \U$17625 ( \17968 , RI9871500_121, \4708 );
nor \U$17626 ( \17969 , \17967 , \17968 );
not \U$17627 ( \17970 , \17969 );
or \U$17628 ( \17971 , \17966 , \17970 );
or \U$17629 ( \17972 , \17969 , \4521 );
nand \U$17630 ( \17973 , \17971 , \17972 );
xor \U$17631 ( \17974 , \17965 , \17973 );
and \U$17632 ( \17975 , \5318 , RI98715f0_123);
and \U$17633 ( \17976 , RI986ead0_31, \5316 );
nor \U$17634 ( \17977 , \17975 , \17976 );
and \U$17635 ( \17978 , \17977 , \5052 );
not \U$17636 ( \17979 , \17977 );
and \U$17637 ( \17980 , \17979 , \5322 );
nor \U$17638 ( \17981 , \17978 , \17980 );
and \U$17639 ( \17982 , \17974 , \17981 );
and \U$17640 ( \17983 , \17965 , \17973 );
or \U$17641 ( \17984 , \17982 , \17983 );
and \U$17642 ( \17985 , \17958 , \17984 );
and \U$17643 ( \17986 , \17932 , \17957 );
or \U$17644 ( \17987 , \17985 , \17986 );
and \U$17645 ( \17988 , \17907 , \17987 );
and \U$17646 ( \17989 , \17833 , \17906 );
or \U$17647 ( \17990 , \17988 , \17989 );
xor \U$17648 ( \17991 , \17750 , \17990 );
xor \U$17649 ( \17992 , \17368 , \17375 );
xor \U$17650 ( \17993 , \17992 , \17383 );
xor \U$17651 ( \17994 , \17287 , \17294 );
xor \U$17652 ( \17995 , \17994 , \17302 );
and \U$17653 ( \17996 , \17993 , \17995 );
xor \U$17654 ( \17997 , \17339 , \17346 );
xor \U$17655 ( \17998 , \17997 , \17354 );
xor \U$17656 ( \17999 , \17287 , \17294 );
xor \U$17657 ( \18000 , \17999 , \17302 );
and \U$17658 ( \18001 , \17998 , \18000 );
and \U$17659 ( \18002 , \17993 , \17998 );
or \U$17660 ( \18003 , \17996 , \18001 , \18002 );
xor \U$17661 ( \18004 , \17452 , \17458 );
xor \U$17662 ( \18005 , \18004 , \17465 );
and \U$17663 ( \18006 , \18003 , \18005 );
xor \U$17664 ( \18007 , \16880 , \16887 );
xor \U$17665 ( \18008 , \18007 , \16895 );
xor \U$17666 ( \18009 , \17124 , \17133 );
xor \U$17667 ( \18010 , \18008 , \18009 );
xor \U$17668 ( \18011 , \17452 , \17458 );
xor \U$17669 ( \18012 , \18011 , \17465 );
and \U$17670 ( \18013 , \18010 , \18012 );
and \U$17671 ( \18014 , \18003 , \18010 );
or \U$17672 ( \18015 , \18006 , \18013 , \18014 );
and \U$17673 ( \18016 , \17991 , \18015 );
and \U$17674 ( \18017 , \17750 , \17990 );
or \U$17675 ( \18018 , \18016 , \18017 );
xor \U$17676 ( \18019 , \17670 , \18018 );
not \U$17677 ( \18020 , \17497 );
xor \U$17678 ( \18021 , \17502 , \17486 );
not \U$17679 ( \18022 , \18021 );
or \U$17680 ( \18023 , \18020 , \18022 );
or \U$17681 ( \18024 , \18021 , \17497 );
nand \U$17682 ( \18025 , \18023 , \18024 );
xor \U$17683 ( \18026 , \16966 , \16971 );
xor \U$17684 ( \18027 , \18026 , \16980 );
xor \U$17685 ( \18028 , \17166 , \17171 );
xor \U$17686 ( \18029 , \18027 , \18028 );
xor \U$17687 ( \18030 , \17224 , \17250 );
xor \U$17688 ( \18031 , \18030 , \17277 );
xor \U$17689 ( \18032 , \18029 , \18031 );
xor \U$17690 ( \18033 , \17183 , \17189 );
xor \U$17691 ( \18034 , \18033 , \17192 );
and \U$17692 ( \18035 , \18032 , \18034 );
and \U$17693 ( \18036 , \18029 , \18031 );
or \U$17694 ( \18037 , \18035 , \18036 );
xor \U$17695 ( \18038 , \18025 , \18037 );
xor \U$17696 ( \18039 , \16941 , \16948 );
xor \U$17697 ( \18040 , \18039 , \16955 );
xor \U$17698 ( \18041 , \17512 , \17519 );
xor \U$17699 ( \18042 , \18040 , \18041 );
and \U$17700 ( \18043 , \18038 , \18042 );
and \U$17701 ( \18044 , \18025 , \18037 );
or \U$17702 ( \18045 , \18043 , \18044 );
and \U$17703 ( \18046 , \18019 , \18045 );
and \U$17704 ( \18047 , \17670 , \18018 );
or \U$17705 ( \18048 , \18046 , \18047 );
and \U$17706 ( \18049 , \17660 , \18048 );
and \U$17707 ( \18050 , \17653 , \17659 );
or \U$17708 ( \18051 , \18049 , \18050 );
nand \U$17709 ( \18052 , \17639 , \18051 );
nand \U$17710 ( \18053 , \17636 , \18052 );
nand \U$17711 ( \18054 , \17619 , \18053 );
nand \U$17712 ( \18055 , \17618 , \18054 );
and \U$17713 ( \18056 , \17612 , \18055 );
xor \U$17714 ( \18057 , \17612 , \18055 );
xor \U$17715 ( \18058 , \17932 , \17957 );
xor \U$17716 ( \18059 , \18058 , \17984 );
xor \U$17717 ( \18060 , \17858 , \17877 );
xor \U$17718 ( \18061 , \18060 , \17903 );
xor \U$17719 ( \18062 , \18059 , \18061 );
xor \U$17720 ( \18063 , \17777 , \17803 );
xor \U$17721 ( \18064 , \18063 , \17830 );
and \U$17722 ( \18065 , \18062 , \18064 );
and \U$17723 ( \18066 , \18059 , \18061 );
or \U$17724 ( \18067 , \18065 , \18066 );
xor \U$17725 ( \18068 , \17386 , \17411 );
xor \U$17726 ( \18069 , \18068 , \17439 );
xor \U$17727 ( \18070 , \18067 , \18069 );
xor \U$17728 ( \18071 , \17695 , \17703 );
xor \U$17729 ( \18072 , \18071 , \17731 );
xor \U$17730 ( \18073 , \17672 , \17674 );
xor \U$17731 ( \18074 , \18073 , \17677 );
and \U$17732 ( \18075 , \18072 , \18074 );
xor \U$17733 ( \18076 , \17393 , \17400 );
xor \U$17734 ( \18077 , \18076 , \17408 );
xor \U$17735 ( \18078 , \17737 , \17742 );
xor \U$17736 ( \18079 , \18077 , \18078 );
xor \U$17737 ( \18080 , \17672 , \17674 );
xor \U$17738 ( \18081 , \18080 , \17677 );
and \U$17739 ( \18082 , \18079 , \18081 );
and \U$17740 ( \18083 , \18072 , \18079 );
or \U$17741 ( \18084 , \18075 , \18082 , \18083 );
and \U$17742 ( \18085 , \18070 , \18084 );
and \U$17743 ( \18086 , \18067 , \18069 );
or \U$17744 ( \18087 , \18085 , \18086 );
xor \U$17745 ( \18088 , \17811 , \17819 );
xor \U$17746 ( \18089 , \18088 , \17827 );
xor \U$17747 ( \18090 , \17784 , \17792 );
xor \U$17748 ( \18091 , \18090 , \17800 );
and \U$17749 ( \18092 , \18089 , \18091 );
xor \U$17750 ( \18093 , \17757 , \17765 );
xor \U$17751 ( \18094 , \18093 , \17774 );
xor \U$17752 ( \18095 , \17784 , \17792 );
xor \U$17753 ( \18096 , \18095 , \17800 );
and \U$17754 ( \18097 , \18094 , \18096 );
and \U$17755 ( \18098 , \18089 , \18094 );
or \U$17756 ( \18099 , \18092 , \18097 , \18098 );
not \U$17757 ( \18100 , \487 );
and \U$17758 ( \18101 , \395 , RI9870420_85);
and \U$17759 ( \18102 , RI9870510_87, \393 );
nor \U$17760 ( \18103 , \18101 , \18102 );
not \U$17761 ( \18104 , \18103 );
or \U$17762 ( \18105 , \18100 , \18104 );
or \U$17763 ( \18106 , \18103 , \386 );
nand \U$17764 ( \18107 , \18105 , \18106 );
not \U$17765 ( \18108 , \456 );
and \U$17766 ( \18109 , \465 , RI98706f0_91);
and \U$17767 ( \18110 , RI9870600_89, \463 );
nor \U$17768 ( \18111 , \18109 , \18110 );
not \U$17769 ( \18112 , \18111 );
or \U$17770 ( \18113 , \18108 , \18112 );
or \U$17771 ( \18114 , \18111 , \454 );
nand \U$17772 ( \18115 , \18113 , \18114 );
xor \U$17773 ( \18116 , \18107 , \18115 );
not \U$17774 ( \18117 , \367 );
and \U$17775 ( \18118 , \376 , RI9870330_83);
and \U$17776 ( \18119 , RI9870240_81, \374 );
nor \U$17777 ( \18120 , \18118 , \18119 );
not \U$17778 ( \18121 , \18120 );
or \U$17779 ( \18122 , \18117 , \18121 );
or \U$17780 ( \18123 , \18120 , \365 );
nand \U$17781 ( \18124 , \18122 , \18123 );
and \U$17782 ( \18125 , \18116 , \18124 );
and \U$17783 ( \18126 , \18107 , \18115 );
or \U$17784 ( \18127 , \18125 , \18126 );
xor \U$17785 ( \18128 , \17686 , \17694 );
xor \U$17786 ( \18129 , \18127 , \18128 );
xor \U$17787 ( \18130 , \17711 , \17719 );
xor \U$17788 ( \18131 , \18130 , \17728 );
and \U$17789 ( \18132 , \18129 , \18131 );
and \U$17790 ( \18133 , \18127 , \18128 );
or \U$17791 ( \18134 , \18132 , \18133 );
xor \U$17792 ( \18135 , \18099 , \18134 );
xor \U$17793 ( \18136 , \17939 , \17946 );
xor \U$17794 ( \18137 , \18136 , \17954 );
xor \U$17795 ( \18138 , \17965 , \17973 );
xor \U$17796 ( \18139 , \18138 , \17981 );
and \U$17797 ( \18140 , \18137 , \18139 );
xor \U$17798 ( \18141 , \17914 , \17921 );
xor \U$17799 ( \18142 , \18141 , \17929 );
xor \U$17800 ( \18143 , \17965 , \17973 );
xor \U$17801 ( \18144 , \18143 , \17981 );
and \U$17802 ( \18145 , \18142 , \18144 );
and \U$17803 ( \18146 , \18137 , \18142 );
or \U$17804 ( \18147 , \18140 , \18145 , \18146 );
and \U$17805 ( \18148 , \18135 , \18147 );
and \U$17806 ( \18149 , \18099 , \18134 );
or \U$17807 ( \18150 , \18148 , \18149 );
and \U$17808 ( \18151 , \8486 , RI986f070_43);
and \U$17809 ( \18152 , RI986ef80_41, \8484 );
nor \U$17810 ( \18153 , \18151 , \18152 );
and \U$17811 ( \18154 , \18153 , \8050 );
not \U$17812 ( \18155 , \18153 );
and \U$17813 ( \18156 , \18155 , \8051 );
nor \U$17814 ( \18157 , \18154 , \18156 );
and \U$17815 ( \18158 , \7079 , RI986ee90_39);
and \U$17816 ( \18159 , RI986eda0_37, \7077 );
nor \U$17817 ( \18160 , \18158 , \18159 );
and \U$17818 ( \18161 , \18160 , \6710 );
not \U$17819 ( \18162 , \18160 );
and \U$17820 ( \18163 , \18162 , \6709 );
nor \U$17821 ( \18164 , \18161 , \18163 );
xor \U$17822 ( \18165 , \18157 , \18164 );
and \U$17823 ( \18166 , \7729 , RI986ebc0_33);
and \U$17824 ( \18167 , RI986ecb0_35, \7727 );
nor \U$17825 ( \18168 , \18166 , \18167 );
and \U$17826 ( \18169 , \18168 , \7480 );
not \U$17827 ( \18170 , \18168 );
and \U$17828 ( \18171 , \18170 , \7733 );
nor \U$17829 ( \18172 , \18169 , \18171 );
and \U$17830 ( \18173 , \18165 , \18172 );
and \U$17831 ( \18174 , \18157 , \18164 );
or \U$17832 ( \18175 , \18173 , \18174 );
and \U$17833 ( \18176 , \4203 , RI9871320_117);
and \U$17834 ( \18177 , RI9871410_119, \4201 );
nor \U$17835 ( \18178 , \18176 , \18177 );
and \U$17836 ( \18179 , \18178 , \4207 );
not \U$17837 ( \18180 , \18178 );
and \U$17838 ( \18181 , \18180 , \3922 );
nor \U$17839 ( \18182 , \18179 , \18181 );
not \U$17840 ( \18183 , \3918 );
and \U$17841 ( \18184 , \3683 , RI9871230_115);
and \U$17842 ( \18185 , RI9871140_113, \3681 );
nor \U$17843 ( \18186 , \18184 , \18185 );
not \U$17844 ( \18187 , \18186 );
or \U$17845 ( \18188 , \18183 , \18187 );
or \U$17846 ( \18189 , \18186 , \3412 );
nand \U$17847 ( \18190 , \18188 , \18189 );
xor \U$17848 ( \18191 , \18182 , \18190 );
not \U$17849 ( \18192 , \4519 );
and \U$17850 ( \18193 , \4710 , RI98716e0_125);
and \U$17851 ( \18194 , RI98717d0_127, \4708 );
nor \U$17852 ( \18195 , \18193 , \18194 );
not \U$17853 ( \18196 , \18195 );
or \U$17854 ( \18197 , \18192 , \18196 );
or \U$17855 ( \18198 , \18195 , \4519 );
nand \U$17856 ( \18199 , \18197 , \18198 );
and \U$17857 ( \18200 , \18191 , \18199 );
and \U$17858 ( \18201 , \18182 , \18190 );
or \U$17859 ( \18202 , \18200 , \18201 );
xor \U$17860 ( \18203 , \18175 , \18202 );
and \U$17861 ( \18204 , \6453 , RI986e8f0_27);
and \U$17862 ( \18205 , RI986e800_25, \6451 );
nor \U$17863 ( \18206 , \18204 , \18205 );
and \U$17864 ( \18207 , \18206 , \6190 );
not \U$17865 ( \18208 , \18206 );
and \U$17866 ( \18209 , \18208 , \6180 );
nor \U$17867 ( \18210 , \18207 , \18209 );
and \U$17868 ( \18211 , \5318 , RI9871500_121);
and \U$17869 ( \18212 , RI98715f0_123, \5316 );
nor \U$17870 ( \18213 , \18211 , \18212 );
and \U$17871 ( \18214 , \18213 , \5052 );
not \U$17872 ( \18215 , \18213 );
and \U$17873 ( \18216 , \18215 , \5322 );
nor \U$17874 ( \18217 , \18214 , \18216 );
xor \U$17875 ( \18218 , \18210 , \18217 );
and \U$17876 ( \18219 , \5881 , RI986ead0_31);
and \U$17877 ( \18220 , RI986e9e0_29, \5879 );
nor \U$17878 ( \18221 , \18219 , \18220 );
and \U$17879 ( \18222 , \18221 , \5594 );
not \U$17880 ( \18223 , \18221 );
and \U$17881 ( \18224 , \18223 , \5885 );
nor \U$17882 ( \18225 , \18222 , \18224 );
and \U$17883 ( \18226 , \18218 , \18225 );
and \U$17884 ( \18227 , \18210 , \18217 );
or \U$17885 ( \18228 , \18226 , \18227 );
and \U$17886 ( \18229 , \18203 , \18228 );
and \U$17887 ( \18230 , \18175 , \18202 );
or \U$17888 ( \18231 , \18229 , \18230 );
and \U$17889 ( \18232 , \10424 , RI986e710_23);
and \U$17890 ( \18233 , RI986e620_21, \10422 );
nor \U$17891 ( \18234 , \18232 , \18233 );
and \U$17892 ( \18235 , \18234 , \9840 );
not \U$17893 ( \18236 , \18234 );
and \U$17894 ( \18237 , \18236 , \10428 );
nor \U$17895 ( \18238 , \18235 , \18237 );
and \U$17896 ( \18239 , \9237 , RI986f250_47);
and \U$17897 ( \18240 , RI986f160_45, \9235 );
nor \U$17898 ( \18241 , \18239 , \18240 );
and \U$17899 ( \18242 , \18241 , \9241 );
not \U$17900 ( \18243 , \18241 );
and \U$17901 ( \18244 , \18243 , \8836 );
nor \U$17902 ( \18245 , \18242 , \18244 );
xor \U$17903 ( \18246 , \18238 , \18245 );
and \U$17904 ( \18247 , \9505 , RI986e530_19);
and \U$17905 ( \18248 , RI986e440_17, \9503 );
nor \U$17906 ( \18249 , \18247 , \18248 );
and \U$17907 ( \18250 , \18249 , \9510 );
not \U$17908 ( \18251 , \18249 );
and \U$17909 ( \18252 , \18251 , \9513 );
nor \U$17910 ( \18253 , \18250 , \18252 );
and \U$17911 ( \18254 , \18246 , \18253 );
and \U$17912 ( \18255 , \18238 , \18245 );
or \U$17913 ( \18256 , \18254 , \18255 );
and \U$17914 ( \18257 , \14937 , RI986df90_7);
and \U$17915 ( \18258 , RI986dea0_5, \14935 );
nor \U$17916 ( \18259 , \18257 , \18258 );
and \U$17917 ( \18260 , \18259 , \14539 );
not \U$17918 ( \18261 , \18259 );
and \U$17919 ( \18262 , \18261 , \14538 );
nor \U$17920 ( \18263 , \18260 , \18262 );
not \U$17921 ( \18264 , RI9873558_190);
and \U$17922 ( \18265 , \15780 , RI986ddb0_3);
and \U$17923 ( \18266 , RI9873648_192, RI986dcc0_1);
nor \U$17924 ( \18267 , \18265 , \18266 );
not \U$17925 ( \18268 , \18267 );
or \U$17926 ( \18269 , \18264 , \18268 );
or \U$17927 ( \18270 , \18267 , RI9873558_190);
nand \U$17928 ( \18271 , \18269 , \18270 );
xor \U$17929 ( \18272 , \18263 , \18271 );
and \U$17930 ( \18273 , \13882 , RI986f520_53);
and \U$17931 ( \18274 , RI986f610_55, \13880 );
nor \U$17932 ( \18275 , \18273 , \18274 );
and \U$17933 ( \18276 , \18275 , \13358 );
not \U$17934 ( \18277 , \18275 );
and \U$17935 ( \18278 , \18277 , \13359 );
nor \U$17936 ( \18279 , \18276 , \18278 );
and \U$17937 ( \18280 , \18272 , \18279 );
and \U$17938 ( \18281 , \18263 , \18271 );
or \U$17939 ( \18282 , \18280 , \18281 );
xor \U$17940 ( \18283 , \18256 , \18282 );
and \U$17941 ( \18284 , \13045 , RI986f430_51);
and \U$17942 ( \18285 , RI986f340_49, \13043 );
nor \U$17943 ( \18286 , \18284 , \18285 );
and \U$17944 ( \18287 , \18286 , \13047 );
not \U$17945 ( \18288 , \18286 );
and \U$17946 ( \18289 , \18288 , \12619 );
nor \U$17947 ( \18290 , \18287 , \18289 );
and \U$17948 ( \18291 , \11696 , RI986f7f0_59);
and \U$17949 ( \18292 , RI986f700_57, \11694 );
nor \U$17950 ( \18293 , \18291 , \18292 );
and \U$17951 ( \18294 , \18293 , \10965 );
not \U$17952 ( \18295 , \18293 );
and \U$17953 ( \18296 , \18295 , \11702 );
nor \U$17954 ( \18297 , \18294 , \18296 );
xor \U$17955 ( \18298 , \18290 , \18297 );
and \U$17956 ( \18299 , \12293 , RI986f9d0_63);
and \U$17957 ( \18300 , RI986f8e0_61, \12291 );
nor \U$17958 ( \18301 , \18299 , \18300 );
and \U$17959 ( \18302 , \18301 , \11687 );
not \U$17960 ( \18303 , \18301 );
and \U$17961 ( \18304 , \18303 , \11686 );
nor \U$17962 ( \18305 , \18302 , \18304 );
and \U$17963 ( \18306 , \18298 , \18305 );
and \U$17964 ( \18307 , \18290 , \18297 );
or \U$17965 ( \18308 , \18306 , \18307 );
and \U$17966 ( \18309 , \18283 , \18308 );
and \U$17967 ( \18310 , \18256 , \18282 );
or \U$17968 ( \18311 , \18309 , \18310 );
xor \U$17969 ( \18312 , \18231 , \18311 );
not \U$17970 ( \18313 , \3406 );
and \U$17971 ( \18314 , \3254 , RI9871050_111);
and \U$17972 ( \18315 , RI9870c90_103, \3252 );
nor \U$17973 ( \18316 , \18314 , \18315 );
not \U$17974 ( \18317 , \18316 );
or \U$17975 ( \18318 , \18313 , \18317 );
or \U$17976 ( \18319 , \18316 , \2935 );
nand \U$17977 ( \18320 , \18318 , \18319 );
and \U$17978 ( \18321 , \2274 , RI9870d80_105);
and \U$17979 ( \18322 , RI98709c0_97, \2272 );
nor \U$17980 ( \18323 , \18321 , \18322 );
and \U$17981 ( \18324 , \18323 , \2030 );
not \U$17982 ( \18325 , \18323 );
and \U$17983 ( \18326 , \18325 , \2031 );
nor \U$17984 ( \18327 , \18324 , \18326 );
xor \U$17985 ( \18328 , \18320 , \18327 );
and \U$17986 ( \18329 , \2464 , RI9870e70_107);
and \U$17987 ( \18330 , RI9870ba0_101, \2462 );
nor \U$17988 ( \18331 , \18329 , \18330 );
and \U$17989 ( \18332 , \18331 , \2468 );
not \U$17990 ( \18333 , \18331 );
and \U$17991 ( \18334 , \18333 , \2263 );
nor \U$17992 ( \18335 , \18332 , \18334 );
and \U$17993 ( \18336 , \18328 , \18335 );
and \U$17994 ( \18337 , \18320 , \18327 );
or \U$17995 ( \18338 , \18336 , \18337 );
not \U$17996 ( \18339 , \1128 );
and \U$17997 ( \18340 , \1293 , RI986fd90_71);
and \U$17998 ( \18341 , RI986fca0_69, \1291 );
nor \U$17999 ( \18342 , \18340 , \18341 );
not \U$18000 ( \18343 , \18342 );
or \U$18001 ( \18344 , \18339 , \18343 );
or \U$18002 ( \18345 , \18342 , \1301 );
nand \U$18003 ( \18346 , \18344 , \18345 );
and \U$18004 ( \18347 , \776 , RI986fac0_65);
and \U$18005 ( \18348 , RI986fbb0_67, \774 );
nor \U$18006 ( \18349 , \18347 , \18348 );
and \U$18007 ( \18350 , \18349 , \474 );
not \U$18008 ( \18351 , \18349 );
and \U$18009 ( \18352 , \18351 , \451 );
nor \U$18010 ( \18353 , \18350 , \18352 );
xor \U$18011 ( \18354 , \18346 , \18353 );
and \U$18012 ( \18355 , \438 , RI98708d0_95);
and \U$18013 ( \18356 , RI98707e0_93, \436 );
nor \U$18014 ( \18357 , \18355 , \18356 );
and \U$18015 ( \18358 , \18357 , \444 );
not \U$18016 ( \18359 , \18357 );
and \U$18017 ( \18360 , \18359 , \443 );
nor \U$18018 ( \18361 , \18358 , \18360 );
and \U$18019 ( \18362 , \18354 , \18361 );
and \U$18020 ( \18363 , \18346 , \18353 );
or \U$18021 ( \18364 , \18362 , \18363 );
xor \U$18022 ( \18365 , \18338 , \18364 );
and \U$18023 ( \18366 , \1311 , RI9870060_77);
and \U$18024 ( \18367 , RI9870150_79, \1309 );
nor \U$18025 ( \18368 , \18366 , \18367 );
and \U$18026 ( \18369 , \18368 , \1458 );
not \U$18027 ( \18370 , \18368 );
and \U$18028 ( \18371 , \18370 , \1318 );
nor \U$18029 ( \18372 , \18369 , \18371 );
and \U$18030 ( \18373 , \1329 , RI986ff70_75);
and \U$18031 ( \18374 , RI986fe80_73, \1327 );
nor \U$18032 ( \18375 , \18373 , \18374 );
and \U$18033 ( \18376 , \18375 , \1336 );
not \U$18034 ( \18377 , \18375 );
and \U$18035 ( \18378 , \18377 , \1337 );
nor \U$18036 ( \18379 , \18376 , \18378 );
xor \U$18037 ( \18380 , \18372 , \18379 );
not \U$18038 ( \18381 , \1462 );
and \U$18039 ( \18382 , \2042 , RI9870f60_109);
and \U$18040 ( \18383 , RI9870ab0_99, \2040 );
nor \U$18041 ( \18384 , \18382 , \18383 );
not \U$18042 ( \18385 , \18384 );
or \U$18043 ( \18386 , \18381 , \18385 );
or \U$18044 ( \18387 , \18384 , \1462 );
nand \U$18045 ( \18388 , \18386 , \18387 );
and \U$18046 ( \18389 , \18380 , \18388 );
and \U$18047 ( \18390 , \18372 , \18379 );
or \U$18048 ( \18391 , \18389 , \18390 );
and \U$18049 ( \18392 , \18365 , \18391 );
and \U$18050 ( \18393 , \18338 , \18364 );
or \U$18051 ( \18394 , \18392 , \18393 );
and \U$18052 ( \18395 , \18312 , \18394 );
and \U$18053 ( \18396 , \18231 , \18311 );
or \U$18054 ( \18397 , \18395 , \18396 );
xor \U$18055 ( \18398 , \18150 , \18397 );
xor \U$18056 ( \18399 , \17866 , \361 );
xor \U$18057 ( \18400 , \18399 , \17874 );
xor \U$18058 ( \18401 , \17885 , \17892 );
xor \U$18059 ( \18402 , \18401 , \17900 );
xor \U$18060 ( \18403 , \18400 , \18402 );
xor \U$18061 ( \18404 , \17840 , \17847 );
xor \U$18062 ( \18405 , \18404 , \17855 );
and \U$18063 ( \18406 , \18403 , \18405 );
and \U$18064 ( \18407 , \18400 , \18402 );
or \U$18065 ( \18408 , \18406 , \18407 );
xor \U$18066 ( \18409 , \17312 , \17320 );
xor \U$18067 ( \18410 , \18409 , \17328 );
xor \U$18068 ( \18411 , \18408 , \18410 );
xor \U$18069 ( \18412 , \17287 , \17294 );
xor \U$18070 ( \18413 , \18412 , \17302 );
xor \U$18071 ( \18414 , \17993 , \17998 );
xor \U$18072 ( \18415 , \18413 , \18414 );
and \U$18073 ( \18416 , \18411 , \18415 );
and \U$18074 ( \18417 , \18408 , \18410 );
or \U$18075 ( \18418 , \18416 , \18417 );
and \U$18076 ( \18419 , \18398 , \18418 );
and \U$18077 ( \18420 , \18150 , \18397 );
or \U$18078 ( \18421 , \18419 , \18420 );
xor \U$18079 ( \18422 , \18087 , \18421 );
xor \U$18080 ( \18423 , \17305 , \17331 );
xor \U$18081 ( \18424 , \18423 , \17357 );
xor \U$18082 ( \18425 , \18029 , \18031 );
xor \U$18083 ( \18426 , \18425 , \18034 );
and \U$18084 ( \18427 , \18424 , \18426 );
xor \U$18085 ( \18428 , \17452 , \17458 );
xor \U$18086 ( \18429 , \18428 , \17465 );
xor \U$18087 ( \18430 , \18003 , \18010 );
xor \U$18088 ( \18431 , \18429 , \18430 );
xor \U$18089 ( \18432 , \18029 , \18031 );
xor \U$18090 ( \18433 , \18432 , \18034 );
and \U$18091 ( \18434 , \18431 , \18433 );
and \U$18092 ( \18435 , \18424 , \18431 );
or \U$18093 ( \18436 , \18427 , \18434 , \18435 );
xor \U$18094 ( \18437 , \18422 , \18436 );
not \U$18095 ( \18438 , \2935 );
and \U$18096 ( \18439 , \3254 , RI9870ba0_101);
and \U$18097 ( \18440 , RI9871050_111, \3252 );
nor \U$18098 ( \18441 , \18439 , \18440 );
not \U$18099 ( \18442 , \18441 );
or \U$18100 ( \18443 , \18438 , \18442 );
or \U$18101 ( \18444 , \18441 , \2935 );
nand \U$18102 ( \18445 , \18443 , \18444 );
and \U$18103 ( \18446 , \2464 , RI98709c0_97);
and \U$18104 ( \18447 , RI9870e70_107, \2462 );
nor \U$18105 ( \18448 , \18446 , \18447 );
and \U$18106 ( \18449 , \18448 , \2468 );
not \U$18107 ( \18450 , \18448 );
and \U$18108 ( \18451 , \18450 , \2263 );
nor \U$18109 ( \18452 , \18449 , \18451 );
xor \U$18110 ( \18453 , \18445 , \18452 );
not \U$18111 ( \18454 , \3412 );
and \U$18112 ( \18455 , \3683 , RI9870c90_103);
and \U$18113 ( \18456 , RI9871230_115, \3681 );
nor \U$18114 ( \18457 , \18455 , \18456 );
not \U$18115 ( \18458 , \18457 );
or \U$18116 ( \18459 , \18454 , \18458 );
or \U$18117 ( \18460 , \18457 , \3918 );
nand \U$18118 ( \18461 , \18459 , \18460 );
and \U$18119 ( \18462 , \18453 , \18461 );
and \U$18120 ( \18463 , \18445 , \18452 );
or \U$18121 ( \18464 , \18462 , \18463 );
and \U$18122 ( \18465 , \1311 , RI986fe80_73);
and \U$18123 ( \18466 , RI9870060_77, \1309 );
nor \U$18124 ( \18467 , \18465 , \18466 );
and \U$18125 ( \18468 , \18467 , \1458 );
not \U$18126 ( \18469 , \18467 );
and \U$18127 ( \18470 , \18469 , \1318 );
nor \U$18128 ( \18471 , \18468 , \18470 );
not \U$18129 ( \18472 , \1462 );
and \U$18130 ( \18473 , \2042 , RI9870150_79);
and \U$18131 ( \18474 , RI9870f60_109, \2040 );
nor \U$18132 ( \18475 , \18473 , \18474 );
not \U$18133 ( \18476 , \18475 );
or \U$18134 ( \18477 , \18472 , \18476 );
or \U$18135 ( \18478 , \18475 , \2034 );
nand \U$18136 ( \18479 , \18477 , \18478 );
xor \U$18137 ( \18480 , \18471 , \18479 );
and \U$18138 ( \18481 , \2274 , RI9870ab0_99);
and \U$18139 ( \18482 , RI9870d80_105, \2272 );
nor \U$18140 ( \18483 , \18481 , \18482 );
and \U$18141 ( \18484 , \18483 , \2030 );
not \U$18142 ( \18485 , \18483 );
and \U$18143 ( \18486 , \18485 , \2031 );
nor \U$18144 ( \18487 , \18484 , \18486 );
and \U$18145 ( \18488 , \18480 , \18487 );
and \U$18146 ( \18489 , \18471 , \18479 );
or \U$18147 ( \18490 , \18488 , \18489 );
xor \U$18148 ( \18491 , \18464 , \18490 );
and \U$18149 ( \18492 , \776 , RI98707e0_93);
and \U$18150 ( \18493 , RI986fac0_65, \774 );
nor \U$18151 ( \18494 , \18492 , \18493 );
and \U$18152 ( \18495 , \18494 , \474 );
not \U$18153 ( \18496 , \18494 );
and \U$18154 ( \18497 , \18496 , \451 );
nor \U$18155 ( \18498 , \18495 , \18497 );
not \U$18156 ( \18499 , \1301 );
and \U$18157 ( \18500 , \1293 , RI986fbb0_67);
and \U$18158 ( \18501 , RI986fd90_71, \1291 );
nor \U$18159 ( \18502 , \18500 , \18501 );
not \U$18160 ( \18503 , \18502 );
or \U$18161 ( \18504 , \18499 , \18503 );
or \U$18162 ( \18505 , \18502 , \1301 );
nand \U$18163 ( \18506 , \18504 , \18505 );
xor \U$18164 ( \18507 , \18498 , \18506 );
and \U$18165 ( \18508 , \1329 , RI986fca0_69);
and \U$18166 ( \18509 , RI986ff70_75, \1327 );
nor \U$18167 ( \18510 , \18508 , \18509 );
and \U$18168 ( \18511 , \18510 , \1336 );
not \U$18169 ( \18512 , \18510 );
and \U$18170 ( \18513 , \18512 , \1337 );
nor \U$18171 ( \18514 , \18511 , \18513 );
and \U$18172 ( \18515 , \18507 , \18514 );
and \U$18173 ( \18516 , \18498 , \18506 );
or \U$18174 ( \18517 , \18515 , \18516 );
xor \U$18175 ( \18518 , \18491 , \18517 );
xor \U$18176 ( \18519 , \18320 , \18327 );
xor \U$18177 ( \18520 , \18519 , \18335 );
xor \U$18178 ( \18521 , \18372 , \18379 );
xor \U$18179 ( \18522 , \18521 , \18388 );
xor \U$18180 ( \18523 , \18520 , \18522 );
xor \U$18181 ( \18524 , \18182 , \18190 );
xor \U$18182 ( \18525 , \18524 , \18199 );
xor \U$18183 ( \18526 , \18523 , \18525 );
and \U$18184 ( \18527 , \18518 , \18526 );
xor \U$18185 ( \18528 , \18107 , \18115 );
xor \U$18186 ( \18529 , \18528 , \18124 );
and \U$18187 ( \18530 , \438 , RI9870600_89);
and \U$18188 ( \18531 , RI98708d0_95, \436 );
nor \U$18189 ( \18532 , \18530 , \18531 );
and \U$18190 ( \18533 , \18532 , \444 );
not \U$18191 ( \18534 , \18532 );
and \U$18192 ( \18535 , \18534 , \443 );
nor \U$18193 ( \18536 , \18533 , \18535 );
not \U$18194 ( \18537 , \454 );
and \U$18195 ( \18538 , \465 , RI9870240_81);
and \U$18196 ( \18539 , RI98706f0_91, \463 );
nor \U$18197 ( \18540 , \18538 , \18539 );
not \U$18198 ( \18541 , \18540 );
or \U$18199 ( \18542 , \18537 , \18541 );
or \U$18200 ( \18543 , \18540 , \454 );
nand \U$18201 ( \18544 , \18542 , \18543 );
xor \U$18202 ( \18545 , \18536 , \18544 );
not \U$18203 ( \18546 , \367 );
and \U$18204 ( \18547 , \376 , RI9870510_87);
and \U$18205 ( \18548 , RI9870330_83, \374 );
nor \U$18206 ( \18549 , \18547 , \18548 );
not \U$18207 ( \18550 , \18549 );
or \U$18208 ( \18551 , \18546 , \18550 );
or \U$18209 ( \18552 , \18549 , \367 );
nand \U$18210 ( \18553 , \18551 , \18552 );
and \U$18211 ( \18554 , \18545 , \18553 );
and \U$18212 ( \18555 , \18536 , \18544 );
or \U$18213 ( \18556 , \18554 , \18555 );
xor \U$18214 ( \18557 , \18346 , \18353 );
xor \U$18215 ( \18558 , \18557 , \18361 );
xor \U$18216 ( \18559 , \18556 , \18558 );
xor \U$18217 ( \18560 , \18529 , \18559 );
xor \U$18218 ( \18561 , \18520 , \18522 );
xor \U$18219 ( \18562 , \18561 , \18525 );
and \U$18220 ( \18563 , \18560 , \18562 );
and \U$18221 ( \18564 , \18518 , \18560 );
or \U$18222 ( \18565 , \18527 , \18563 , \18564 );
xor \U$18223 ( \18566 , \18256 , \18282 );
xor \U$18224 ( \18567 , \18566 , \18308 );
xor \U$18225 ( \18568 , \18565 , \18567 );
xor \U$18226 ( \18569 , \18175 , \18202 );
xor \U$18227 ( \18570 , \18569 , \18228 );
xor \U$18228 ( \18571 , \18338 , \18364 );
xor \U$18229 ( \18572 , \18571 , \18391 );
xor \U$18230 ( \18573 , \18127 , \18128 );
xor \U$18231 ( \18574 , \18573 , \18131 );
xor \U$18232 ( \18575 , \18572 , \18574 );
xor \U$18233 ( \18576 , \18570 , \18575 );
and \U$18234 ( \18577 , \18568 , \18576 );
and \U$18235 ( \18578 , \18565 , \18567 );
or \U$18236 ( \18579 , \18577 , \18578 );
xor \U$18237 ( \18580 , \18290 , \18297 );
xor \U$18238 ( \18581 , \18580 , \18305 );
xor \U$18239 ( \18582 , \18263 , \18271 );
xor \U$18240 ( \18583 , \18582 , \18279 );
xor \U$18241 ( \18584 , \18581 , \18583 );
xor \U$18242 ( \18585 , \18238 , \18245 );
xor \U$18243 ( \18586 , \18585 , \18253 );
xor \U$18244 ( \18587 , \18210 , \18217 );
xor \U$18245 ( \18588 , \18587 , \18225 );
xor \U$18246 ( \18589 , \18157 , \18164 );
xor \U$18247 ( \18590 , \18589 , \18172 );
xor \U$18248 ( \18591 , \18588 , \18590 );
xor \U$18249 ( \18592 , \18586 , \18591 );
and \U$18250 ( \18593 , \18584 , \18592 );
and \U$18251 ( \18594 , \18581 , \18583 );
or \U$18252 ( \18595 , \18593 , \18594 );
and \U$18253 ( \18596 , \6453 , RI986ead0_31);
and \U$18254 ( \18597 , RI986e9e0_29, \6451 );
nor \U$18255 ( \18598 , \18596 , \18597 );
and \U$18256 ( \18599 , \18598 , \6190 );
not \U$18257 ( \18600 , \18598 );
and \U$18258 ( \18601 , \18600 , \6180 );
nor \U$18259 ( \18602 , \18599 , \18601 );
and \U$18260 ( \18603 , \5318 , RI98716e0_125);
and \U$18261 ( \18604 , RI98717d0_127, \5316 );
nor \U$18262 ( \18605 , \18603 , \18604 );
and \U$18263 ( \18606 , \18605 , \5052 );
not \U$18264 ( \18607 , \18605 );
and \U$18265 ( \18608 , \18607 , \5322 );
nor \U$18266 ( \18609 , \18606 , \18608 );
xor \U$18267 ( \18610 , \18602 , \18609 );
and \U$18268 ( \18611 , \5881 , RI9871500_121);
and \U$18269 ( \18612 , RI98715f0_123, \5879 );
nor \U$18270 ( \18613 , \18611 , \18612 );
and \U$18271 ( \18614 , \18613 , \5594 );
not \U$18272 ( \18615 , \18613 );
and \U$18273 ( \18616 , \18615 , \5885 );
nor \U$18274 ( \18617 , \18614 , \18616 );
and \U$18275 ( \18618 , \18610 , \18617 );
and \U$18276 ( \18619 , \18602 , \18609 );
or \U$18277 ( \18620 , \18618 , \18619 );
not \U$18278 ( \18621 , \3412 );
and \U$18279 ( \18622 , \3683 , RI9871050_111);
and \U$18280 ( \18623 , RI9870c90_103, \3681 );
nor \U$18281 ( \18624 , \18622 , \18623 );
not \U$18282 ( \18625 , \18624 );
or \U$18283 ( \18626 , \18621 , \18625 );
or \U$18284 ( \18627 , \18624 , \3412 );
nand \U$18285 ( \18628 , \18626 , \18627 );
and \U$18286 ( \18629 , \4203 , RI9871230_115);
and \U$18287 ( \18630 , RI9871140_113, \4201 );
nor \U$18288 ( \18631 , \18629 , \18630 );
and \U$18289 ( \18632 , \18631 , \4207 );
not \U$18290 ( \18633 , \18631 );
and \U$18291 ( \18634 , \18633 , \3922 );
nor \U$18292 ( \18635 , \18632 , \18634 );
xor \U$18293 ( \18636 , \18628 , \18635 );
not \U$18294 ( \18637 , \4521 );
and \U$18295 ( \18638 , \4710 , RI9871320_117);
and \U$18296 ( \18639 , RI9871410_119, \4708 );
nor \U$18297 ( \18640 , \18638 , \18639 );
not \U$18298 ( \18641 , \18640 );
or \U$18299 ( \18642 , \18637 , \18641 );
or \U$18300 ( \18643 , \18640 , \4519 );
nand \U$18301 ( \18644 , \18642 , \18643 );
and \U$18302 ( \18645 , \18636 , \18644 );
and \U$18303 ( \18646 , \18628 , \18635 );
or \U$18304 ( \18647 , \18645 , \18646 );
xor \U$18305 ( \18648 , \18620 , \18647 );
and \U$18306 ( \18649 , \7079 , RI986e8f0_27);
and \U$18307 ( \18650 , RI986e800_25, \7077 );
nor \U$18308 ( \18651 , \18649 , \18650 );
and \U$18309 ( \18652 , \18651 , \6710 );
not \U$18310 ( \18653 , \18651 );
and \U$18311 ( \18654 , \18653 , \6709 );
nor \U$18312 ( \18655 , \18652 , \18654 );
and \U$18313 ( \18656 , \7729 , RI986ee90_39);
and \U$18314 ( \18657 , RI986eda0_37, \7727 );
nor \U$18315 ( \18658 , \18656 , \18657 );
and \U$18316 ( \18659 , \18658 , \7480 );
not \U$18317 ( \18660 , \18658 );
and \U$18318 ( \18661 , \18660 , \7733 );
nor \U$18319 ( \18662 , \18659 , \18661 );
xor \U$18320 ( \18663 , \18655 , \18662 );
and \U$18321 ( \18664 , \8486 , RI986ebc0_33);
and \U$18322 ( \18665 , RI986ecb0_35, \8484 );
nor \U$18323 ( \18666 , \18664 , \18665 );
and \U$18324 ( \18667 , \18666 , \8050 );
not \U$18325 ( \18668 , \18666 );
and \U$18326 ( \18669 , \18668 , \8051 );
nor \U$18327 ( \18670 , \18667 , \18669 );
and \U$18328 ( \18671 , \18663 , \18670 );
and \U$18329 ( \18672 , \18655 , \18662 );
or \U$18330 ( \18673 , \18671 , \18672 );
and \U$18331 ( \18674 , \18648 , \18673 );
and \U$18332 ( \18675 , \18620 , \18647 );
or \U$18333 ( \18676 , \18674 , \18675 );
and \U$18334 ( \18677 , \13045 , RI986f9d0_63);
and \U$18335 ( \18678 , RI986f8e0_61, \13043 );
nor \U$18336 ( \18679 , \18677 , \18678 );
and \U$18337 ( \18680 , \18679 , \13047 );
not \U$18338 ( \18681 , \18679 );
and \U$18339 ( \18682 , \18681 , \12619 );
nor \U$18340 ( \18683 , \18680 , \18682 );
and \U$18341 ( \18684 , \11696 , RI986e710_23);
and \U$18342 ( \18685 , RI986e620_21, \11694 );
nor \U$18343 ( \18686 , \18684 , \18685 );
and \U$18344 ( \18687 , \18686 , \10965 );
not \U$18345 ( \18688 , \18686 );
and \U$18346 ( \18689 , \18688 , \11702 );
nor \U$18347 ( \18690 , \18687 , \18689 );
xor \U$18348 ( \18691 , \18683 , \18690 );
and \U$18349 ( \18692 , \12293 , RI986f7f0_59);
and \U$18350 ( \18693 , RI986f700_57, \12291 );
nor \U$18351 ( \18694 , \18692 , \18693 );
and \U$18352 ( \18695 , \18694 , \11687 );
not \U$18353 ( \18696 , \18694 );
and \U$18354 ( \18697 , \18696 , \11686 );
nor \U$18355 ( \18698 , \18695 , \18697 );
and \U$18356 ( \18699 , \18691 , \18698 );
and \U$18357 ( \18700 , \18683 , \18690 );
or \U$18358 ( \18701 , \18699 , \18700 );
and \U$18359 ( \18702 , \13882 , RI986f430_51);
and \U$18360 ( \18703 , RI986f340_49, \13880 );
nor \U$18361 ( \18704 , \18702 , \18703 );
and \U$18362 ( \18705 , \18704 , \13358 );
not \U$18363 ( \18706 , \18704 );
and \U$18364 ( \18707 , \18706 , \13359 );
nor \U$18365 ( \18708 , \18705 , \18707 );
not \U$18366 ( \18709 , RI9873558_190);
and \U$18367 ( \18710 , \15780 , RI986df90_7);
and \U$18368 ( \18711 , RI9873648_192, RI986dea0_5);
nor \U$18369 ( \18712 , \18710 , \18711 );
not \U$18370 ( \18713 , \18712 );
or \U$18371 ( \18714 , \18709 , \18713 );
or \U$18372 ( \18715 , \18712 , RI9873558_190);
nand \U$18373 ( \18716 , \18714 , \18715 );
xor \U$18374 ( \18717 , \18708 , \18716 );
and \U$18375 ( \18718 , \14937 , RI986f520_53);
and \U$18376 ( \18719 , RI986f610_55, \14935 );
nor \U$18377 ( \18720 , \18718 , \18719 );
and \U$18378 ( \18721 , \18720 , \14539 );
not \U$18379 ( \18722 , \18720 );
and \U$18380 ( \18723 , \18722 , \14538 );
nor \U$18381 ( \18724 , \18721 , \18723 );
and \U$18382 ( \18725 , \18717 , \18724 );
and \U$18383 ( \18726 , \18708 , \18716 );
or \U$18384 ( \18727 , \18725 , \18726 );
xor \U$18385 ( \18728 , \18701 , \18727 );
and \U$18386 ( \18729 , \9505 , RI986f250_47);
and \U$18387 ( \18730 , RI986f160_45, \9503 );
nor \U$18388 ( \18731 , \18729 , \18730 );
and \U$18389 ( \18732 , \18731 , \9510 );
not \U$18390 ( \18733 , \18731 );
and \U$18391 ( \18734 , \18733 , \9513 );
nor \U$18392 ( \18735 , \18732 , \18734 );
and \U$18393 ( \18736 , \9237 , RI986f070_43);
and \U$18394 ( \18737 , RI986ef80_41, \9235 );
nor \U$18395 ( \18738 , \18736 , \18737 );
and \U$18396 ( \18739 , \18738 , \9241 );
not \U$18397 ( \18740 , \18738 );
and \U$18398 ( \18741 , \18740 , \8836 );
nor \U$18399 ( \18742 , \18739 , \18741 );
xor \U$18400 ( \18743 , \18735 , \18742 );
and \U$18401 ( \18744 , \10424 , RI986e530_19);
and \U$18402 ( \18745 , RI986e440_17, \10422 );
nor \U$18403 ( \18746 , \18744 , \18745 );
and \U$18404 ( \18747 , \18746 , \9840 );
not \U$18405 ( \18748 , \18746 );
and \U$18406 ( \18749 , \18748 , \10428 );
nor \U$18407 ( \18750 , \18747 , \18749 );
and \U$18408 ( \18751 , \18743 , \18750 );
and \U$18409 ( \18752 , \18735 , \18742 );
or \U$18410 ( \18753 , \18751 , \18752 );
and \U$18411 ( \18754 , \18728 , \18753 );
and \U$18412 ( \18755 , \18701 , \18727 );
or \U$18413 ( \18756 , \18754 , \18755 );
xor \U$18414 ( \18757 , \18676 , \18756 );
and \U$18415 ( \18758 , \1311 , RI986ff70_75);
and \U$18416 ( \18759 , RI986fe80_73, \1309 );
nor \U$18417 ( \18760 , \18758 , \18759 );
and \U$18418 ( \18761 , \18760 , \1319 );
not \U$18419 ( \18762 , \18760 );
and \U$18420 ( \18763 , \18762 , \1315 );
nor \U$18421 ( \18764 , \18761 , \18763 );
and \U$18422 ( \18765 , \1329 , RI986fd90_71);
and \U$18423 ( \18766 , RI986fca0_69, \1327 );
nor \U$18424 ( \18767 , \18765 , \18766 );
and \U$18425 ( \18768 , \18767 , \1336 );
not \U$18426 ( \18769 , \18767 );
and \U$18427 ( \18770 , \18769 , \1337 );
nor \U$18428 ( \18771 , \18768 , \18770 );
xor \U$18429 ( \18772 , \18764 , \18771 );
not \U$18430 ( \18773 , \2034 );
and \U$18431 ( \18774 , \2042 , RI9870060_77);
and \U$18432 ( \18775 , RI9870150_79, \2040 );
nor \U$18433 ( \18776 , \18774 , \18775 );
not \U$18434 ( \18777 , \18776 );
or \U$18435 ( \18778 , \18773 , \18777 );
or \U$18436 ( \18779 , \18776 , \2034 );
nand \U$18437 ( \18780 , \18778 , \18779 );
and \U$18438 ( \18781 , \18772 , \18780 );
and \U$18439 ( \18782 , \18764 , \18771 );
or \U$18440 ( \18783 , \18781 , \18782 );
not \U$18441 ( \18784 , \1301 );
and \U$18442 ( \18785 , \1293 , RI986fac0_65);
and \U$18443 ( \18786 , RI986fbb0_67, \1291 );
nor \U$18444 ( \18787 , \18785 , \18786 );
not \U$18445 ( \18788 , \18787 );
or \U$18446 ( \18789 , \18784 , \18788 );
or \U$18447 ( \18790 , \18787 , \1301 );
nand \U$18448 ( \18791 , \18789 , \18790 );
and \U$18449 ( \18792 , \776 , RI98708d0_95);
and \U$18450 ( \18793 , RI98707e0_93, \774 );
nor \U$18451 ( \18794 , \18792 , \18793 );
and \U$18452 ( \18795 , \18794 , \474 );
not \U$18453 ( \18796 , \18794 );
and \U$18454 ( \18797 , \18796 , \451 );
nor \U$18455 ( \18798 , \18795 , \18797 );
xor \U$18456 ( \18799 , \18791 , \18798 );
and \U$18457 ( \18800 , \438 , RI98706f0_91);
and \U$18458 ( \18801 , RI9870600_89, \436 );
nor \U$18459 ( \18802 , \18800 , \18801 );
and \U$18460 ( \18803 , \18802 , \444 );
not \U$18461 ( \18804 , \18802 );
and \U$18462 ( \18805 , \18804 , \443 );
nor \U$18463 ( \18806 , \18803 , \18805 );
and \U$18464 ( \18807 , \18799 , \18806 );
and \U$18465 ( \18808 , \18791 , \18798 );
or \U$18466 ( \18809 , \18807 , \18808 );
xor \U$18467 ( \18810 , \18783 , \18809 );
not \U$18468 ( \18811 , \3406 );
and \U$18469 ( \18812 , \3254 , RI9870e70_107);
and \U$18470 ( \18813 , RI9870ba0_101, \3252 );
nor \U$18471 ( \18814 , \18812 , \18813 );
not \U$18472 ( \18815 , \18814 );
or \U$18473 ( \18816 , \18811 , \18815 );
or \U$18474 ( \18817 , \18814 , \3406 );
nand \U$18475 ( \18818 , \18816 , \18817 );
and \U$18476 ( \18819 , \2274 , RI9870f60_109);
and \U$18477 ( \18820 , RI9870ab0_99, \2272 );
nor \U$18478 ( \18821 , \18819 , \18820 );
and \U$18479 ( \18822 , \18821 , \2030 );
not \U$18480 ( \18823 , \18821 );
and \U$18481 ( \18824 , \18823 , \2031 );
nor \U$18482 ( \18825 , \18822 , \18824 );
xor \U$18483 ( \18826 , \18818 , \18825 );
and \U$18484 ( \18827 , \2464 , RI9870d80_105);
and \U$18485 ( \18828 , RI98709c0_97, \2462 );
nor \U$18486 ( \18829 , \18827 , \18828 );
and \U$18487 ( \18830 , \18829 , \2468 );
not \U$18488 ( \18831 , \18829 );
and \U$18489 ( \18832 , \18831 , \2263 );
nor \U$18490 ( \18833 , \18830 , \18832 );
and \U$18491 ( \18834 , \18826 , \18833 );
and \U$18492 ( \18835 , \18818 , \18825 );
or \U$18493 ( \18836 , \18834 , \18835 );
and \U$18494 ( \18837 , \18810 , \18836 );
and \U$18495 ( \18838 , \18783 , \18809 );
or \U$18496 ( \18839 , \18837 , \18838 );
and \U$18497 ( \18840 , \18757 , \18839 );
and \U$18498 ( \18841 , \18676 , \18756 );
or \U$18499 ( \18842 , \18840 , \18841 );
xor \U$18500 ( \18843 , \18595 , \18842 );
and \U$18501 ( \18844 , \5881 , RI98715f0_123);
and \U$18502 ( \18845 , RI986ead0_31, \5879 );
nor \U$18503 ( \18846 , \18844 , \18845 );
and \U$18504 ( \18847 , \18846 , \5885 );
not \U$18505 ( \18848 , \18846 );
and \U$18506 ( \18849 , \18848 , \5594 );
nor \U$18507 ( \18850 , \18847 , \18849 );
not \U$18508 ( \18851 , \18850 );
and \U$18509 ( \18852 , \6453 , RI986e9e0_29);
and \U$18510 ( \18853 , RI986e8f0_27, \6451 );
nor \U$18511 ( \18854 , \18852 , \18853 );
and \U$18512 ( \18855 , \18854 , \6180 );
not \U$18513 ( \18856 , \18854 );
and \U$18514 ( \18857 , \18856 , \6190 );
nor \U$18515 ( \18858 , \18855 , \18857 );
and \U$18516 ( \18859 , \7079 , RI986e800_25);
and \U$18517 ( \18860 , RI986ee90_39, \7077 );
nor \U$18518 ( \18861 , \18859 , \18860 );
and \U$18519 ( \18862 , \18861 , \6709 );
not \U$18520 ( \18863 , \18861 );
and \U$18521 ( \18864 , \18863 , \6710 );
nor \U$18522 ( \18865 , \18862 , \18864 );
xor \U$18523 ( \18866 , \18858 , \18865 );
not \U$18524 ( \18867 , \18866 );
or \U$18525 ( \18868 , \18851 , \18867 );
or \U$18526 ( \18869 , \18866 , \18850 );
nand \U$18527 ( \18870 , \18868 , \18869 );
and \U$18528 ( \18871 , \9505 , RI986f160_45);
and \U$18529 ( \18872 , RI986e530_19, \9503 );
nor \U$18530 ( \18873 , \18871 , \18872 );
and \U$18531 ( \18874 , \18873 , \9510 );
not \U$18532 ( \18875 , \18873 );
and \U$18533 ( \18876 , \18875 , \9513 );
nor \U$18534 ( \18877 , \18874 , \18876 );
and \U$18535 ( \18878 , \10424 , RI986e440_17);
and \U$18536 ( \18879 , RI986e710_23, \10422 );
nor \U$18537 ( \18880 , \18878 , \18879 );
and \U$18538 ( \18881 , \18880 , \9840 );
not \U$18539 ( \18882 , \18880 );
and \U$18540 ( \18883 , \18882 , \10428 );
nor \U$18541 ( \18884 , \18881 , \18883 );
xor \U$18542 ( \18885 , \18877 , \18884 );
and \U$18543 ( \18886 , \11696 , RI986e620_21);
and \U$18544 ( \18887 , RI986f7f0_59, \11694 );
nor \U$18545 ( \18888 , \18886 , \18887 );
and \U$18546 ( \18889 , \18888 , \10965 );
not \U$18547 ( \18890 , \18888 );
and \U$18548 ( \18891 , \18890 , \11702 );
nor \U$18549 ( \18892 , \18889 , \18891 );
xor \U$18550 ( \18893 , \18885 , \18892 );
and \U$18551 ( \18894 , \18870 , \18893 );
and \U$18552 ( \18895 , \7729 , RI986eda0_37);
and \U$18553 ( \18896 , RI986ebc0_33, \7727 );
nor \U$18554 ( \18897 , \18895 , \18896 );
and \U$18555 ( \18898 , \18897 , \7733 );
not \U$18556 ( \18899 , \18897 );
and \U$18557 ( \18900 , \18899 , \7480 );
nor \U$18558 ( \18901 , \18898 , \18900 );
not \U$18559 ( \18902 , \18901 );
and \U$18560 ( \18903 , \8486 , RI986ecb0_35);
and \U$18561 ( \18904 , RI986f070_43, \8484 );
nor \U$18562 ( \18905 , \18903 , \18904 );
and \U$18563 ( \18906 , \18905 , \8051 );
not \U$18564 ( \18907 , \18905 );
and \U$18565 ( \18908 , \18907 , \8050 );
nor \U$18566 ( \18909 , \18906 , \18908 );
and \U$18567 ( \18910 , \9237 , RI986ef80_41);
and \U$18568 ( \18911 , RI986f250_47, \9235 );
nor \U$18569 ( \18912 , \18910 , \18911 );
and \U$18570 ( \18913 , \18912 , \8836 );
not \U$18571 ( \18914 , \18912 );
and \U$18572 ( \18915 , \18914 , \9241 );
nor \U$18573 ( \18916 , \18913 , \18915 );
xor \U$18574 ( \18917 , \18909 , \18916 );
not \U$18575 ( \18918 , \18917 );
or \U$18576 ( \18919 , \18902 , \18918 );
or \U$18577 ( \18920 , \18917 , \18901 );
nand \U$18578 ( \18921 , \18919 , \18920 );
xor \U$18579 ( \18922 , \18877 , \18884 );
xor \U$18580 ( \18923 , \18922 , \18892 );
and \U$18581 ( \18924 , \18921 , \18923 );
and \U$18582 ( \18925 , \18870 , \18921 );
or \U$18583 ( \18926 , \18894 , \18924 , \18925 );
xor \U$18584 ( \18927 , \18498 , \18506 );
xor \U$18585 ( \18928 , \18927 , \18514 );
nand \U$18586 ( \18929 , RI9870420_85, \393 );
not \U$18587 ( \18930 , \18929 );
not \U$18588 ( \18931 , \487 );
or \U$18589 ( \18932 , \18930 , \18931 );
or \U$18590 ( \18933 , \386 , \18929 );
nand \U$18591 ( \18934 , \18932 , \18933 );
xor \U$18592 ( \18935 , \18928 , \18934 );
xor \U$18593 ( \18936 , \18536 , \18544 );
xor \U$18594 ( \18937 , \18936 , \18553 );
and \U$18595 ( \18938 , \18935 , \18937 );
and \U$18596 ( \18939 , \18928 , \18934 );
or \U$18597 ( \18940 , \18938 , \18939 );
xor \U$18598 ( \18941 , \18926 , \18940 );
xor \U$18599 ( \18942 , \18471 , \18479 );
xor \U$18600 ( \18943 , \18942 , \18487 );
xor \U$18601 ( \18944 , \18445 , \18452 );
xor \U$18602 ( \18945 , \18944 , \18461 );
and \U$18603 ( \18946 , \18943 , \18945 );
and \U$18604 ( \18947 , \4203 , RI9871140_113);
and \U$18605 ( \18948 , RI9871320_117, \4201 );
nor \U$18606 ( \18949 , \18947 , \18948 );
and \U$18607 ( \18950 , \18949 , \3922 );
not \U$18608 ( \18951 , \18949 );
and \U$18609 ( \18952 , \18951 , \4207 );
nor \U$18610 ( \18953 , \18950 , \18952 );
not \U$18611 ( \18954 , \18953 );
and \U$18612 ( \18955 , \4710 , RI9871410_119);
and \U$18613 ( \18956 , RI98716e0_125, \4708 );
nor \U$18614 ( \18957 , \18955 , \18956 );
not \U$18615 ( \18958 , \18957 );
not \U$18616 ( \18959 , \4521 );
and \U$18617 ( \18960 , \18958 , \18959 );
and \U$18618 ( \18961 , \18957 , \4521 );
nor \U$18619 ( \18962 , \18960 , \18961 );
and \U$18620 ( \18963 , \5318 , RI98717d0_127);
and \U$18621 ( \18964 , RI9871500_121, \5316 );
nor \U$18622 ( \18965 , \18963 , \18964 );
and \U$18623 ( \18966 , \18965 , \5322 );
not \U$18624 ( \18967 , \18965 );
and \U$18625 ( \18968 , \18967 , \5052 );
nor \U$18626 ( \18969 , \18966 , \18968 );
xor \U$18627 ( \18970 , \18962 , \18969 );
not \U$18628 ( \18971 , \18970 );
or \U$18629 ( \18972 , \18954 , \18971 );
or \U$18630 ( \18973 , \18970 , \18953 );
nand \U$18631 ( \18974 , \18972 , \18973 );
xor \U$18632 ( \18975 , \18445 , \18452 );
xor \U$18633 ( \18976 , \18975 , \18461 );
and \U$18634 ( \18977 , \18974 , \18976 );
and \U$18635 ( \18978 , \18943 , \18974 );
or \U$18636 ( \18979 , \18946 , \18977 , \18978 );
and \U$18637 ( \18980 , \18941 , \18979 );
and \U$18638 ( \18981 , \18926 , \18940 );
or \U$18639 ( \18982 , \18980 , \18981 );
and \U$18640 ( \18983 , \18843 , \18982 );
and \U$18641 ( \18984 , \18595 , \18842 );
or \U$18642 ( \18985 , \18983 , \18984 );
xor \U$18643 ( \18986 , \18579 , \18985 );
not \U$18644 ( \18987 , \18953 );
not \U$18645 ( \18988 , \18962 );
and \U$18646 ( \18989 , \18987 , \18988 );
and \U$18647 ( \18990 , \18962 , \18953 );
nor \U$18648 ( \18991 , \18990 , \18969 );
nor \U$18649 ( \18992 , \18989 , \18991 );
not \U$18650 ( \18993 , \18850 );
not \U$18651 ( \18994 , \18858 );
and \U$18652 ( \18995 , \18993 , \18994 );
and \U$18653 ( \18996 , \18858 , \18850 );
nor \U$18654 ( \18997 , \18996 , \18865 );
nor \U$18655 ( \18998 , \18995 , \18997 );
xor \U$18656 ( \18999 , \18992 , \18998 );
not \U$18657 ( \19000 , \18901 );
not \U$18658 ( \19001 , \18909 );
and \U$18659 ( \19002 , \19000 , \19001 );
and \U$18660 ( \19003 , \18909 , \18901 );
nor \U$18661 ( \19004 , \19003 , \18916 );
nor \U$18662 ( \19005 , \19002 , \19004 );
and \U$18663 ( \19006 , \18999 , \19005 );
and \U$18664 ( \19007 , \18992 , \18998 );
nor \U$18665 ( \19008 , \19006 , \19007 );
xor \U$18666 ( \19009 , \18877 , \18884 );
and \U$18667 ( \19010 , \19009 , \18892 );
and \U$18668 ( \19011 , \18877 , \18884 );
or \U$18669 ( \19012 , \19010 , \19011 );
not \U$18670 ( \19013 , RI9873558_190);
and \U$18671 ( \19014 , \15780 , RI986dea0_5);
and \U$18672 ( \19015 , RI9873648_192, RI986ddb0_3);
nor \U$18673 ( \19016 , \19014 , \19015 );
not \U$18674 ( \19017 , \19016 );
or \U$18675 ( \19018 , \19013 , \19017 );
or \U$18676 ( \19019 , \19016 , RI9873558_190);
nand \U$18677 ( \19020 , \19018 , \19019 );
xor \U$18678 ( \19021 , \19020 , \487 );
and \U$18679 ( \19022 , \14937 , RI986f610_55);
and \U$18680 ( \19023 , RI986df90_7, \14935 );
nor \U$18681 ( \19024 , \19022 , \19023 );
and \U$18682 ( \19025 , \19024 , \14539 );
not \U$18683 ( \19026 , \19024 );
and \U$18684 ( \19027 , \19026 , \14538 );
nor \U$18685 ( \19028 , \19025 , \19027 );
and \U$18686 ( \19029 , \19021 , \19028 );
and \U$18687 ( \19030 , \19020 , \487 );
or \U$18688 ( \19031 , \19029 , \19030 );
xor \U$18689 ( \19032 , \19012 , \19031 );
and \U$18690 ( \19033 , \13045 , RI986f8e0_61);
and \U$18691 ( \19034 , RI986f430_51, \13043 );
nor \U$18692 ( \19035 , \19033 , \19034 );
and \U$18693 ( \19036 , \19035 , \13047 );
not \U$18694 ( \19037 , \19035 );
and \U$18695 ( \19038 , \19037 , \12619 );
nor \U$18696 ( \19039 , \19036 , \19038 );
and \U$18697 ( \19040 , \12293 , RI986f700_57);
and \U$18698 ( \19041 , RI986f9d0_63, \12291 );
nor \U$18699 ( \19042 , \19040 , \19041 );
and \U$18700 ( \19043 , \19042 , \11687 );
not \U$18701 ( \19044 , \19042 );
and \U$18702 ( \19045 , \19044 , \11686 );
nor \U$18703 ( \19046 , \19043 , \19045 );
xor \U$18704 ( \19047 , \19039 , \19046 );
and \U$18705 ( \19048 , \13882 , RI986f340_49);
and \U$18706 ( \19049 , RI986f520_53, \13880 );
nor \U$18707 ( \19050 , \19048 , \19049 );
and \U$18708 ( \19051 , \19050 , \13358 );
not \U$18709 ( \19052 , \19050 );
and \U$18710 ( \19053 , \19052 , \13359 );
nor \U$18711 ( \19054 , \19051 , \19053 );
and \U$18712 ( \19055 , \19047 , \19054 );
and \U$18713 ( \19056 , \19039 , \19046 );
or \U$18714 ( \19057 , \19055 , \19056 );
and \U$18715 ( \19058 , \19032 , \19057 );
and \U$18716 ( \19059 , \19012 , \19031 );
or \U$18717 ( \19060 , \19058 , \19059 );
xor \U$18718 ( \19061 , \19008 , \19060 );
xor \U$18719 ( \19062 , \18464 , \18490 );
and \U$18720 ( \19063 , \19062 , \18517 );
and \U$18721 ( \19064 , \18464 , \18490 );
or \U$18722 ( \19065 , \19063 , \19064 );
xor \U$18723 ( \19066 , \19061 , \19065 );
xor \U$18724 ( \19067 , \18520 , \18522 );
and \U$18725 ( \19068 , \19067 , \18525 );
and \U$18726 ( \19069 , \18520 , \18522 );
or \U$18727 ( \19070 , \19068 , \19069 );
xor \U$18728 ( \19071 , \18107 , \18115 );
xor \U$18729 ( \19072 , \19071 , \18124 );
and \U$18730 ( \19073 , \18556 , \19072 );
xor \U$18731 ( \19074 , \18107 , \18115 );
xor \U$18732 ( \19075 , \19074 , \18124 );
and \U$18733 ( \19076 , \18558 , \19075 );
and \U$18734 ( \19077 , \18556 , \18558 );
or \U$18735 ( \19078 , \19073 , \19076 , \19077 );
xor \U$18736 ( \19079 , \19070 , \19078 );
xor \U$18737 ( \19080 , \18238 , \18245 );
xor \U$18738 ( \19081 , \19080 , \18253 );
and \U$18739 ( \19082 , \18588 , \19081 );
xor \U$18740 ( \19083 , \18238 , \18245 );
xor \U$18741 ( \19084 , \19083 , \18253 );
and \U$18742 ( \19085 , \18590 , \19084 );
and \U$18743 ( \19086 , \18588 , \18590 );
or \U$18744 ( \19087 , \19082 , \19085 , \19086 );
xor \U$18745 ( \19088 , \19079 , \19087 );
and \U$18746 ( \19089 , \19066 , \19088 );
xor \U$18747 ( \19090 , \18400 , \18402 );
xor \U$18748 ( \19091 , \19090 , \18405 );
xor \U$18749 ( \19092 , \17784 , \17792 );
xor \U$18750 ( \19093 , \19092 , \17800 );
xor \U$18751 ( \19094 , \18089 , \18094 );
xor \U$18752 ( \19095 , \19093 , \19094 );
xor \U$18753 ( \19096 , \17965 , \17973 );
xor \U$18754 ( \19097 , \19096 , \17981 );
xor \U$18755 ( \19098 , \18137 , \18142 );
xor \U$18756 ( \19099 , \19097 , \19098 );
xor \U$18757 ( \19100 , \19095 , \19099 );
xor \U$18758 ( \19101 , \19091 , \19100 );
xor \U$18759 ( \19102 , \19070 , \19078 );
xor \U$18760 ( \19103 , \19102 , \19087 );
and \U$18761 ( \19104 , \19101 , \19103 );
and \U$18762 ( \19105 , \19066 , \19101 );
or \U$18763 ( \19106 , \19089 , \19104 , \19105 );
and \U$18764 ( \19107 , \18986 , \19106 );
and \U$18765 ( \19108 , \18579 , \18985 );
or \U$18766 ( \19109 , \19107 , \19108 );
xor \U$18767 ( \19110 , \18067 , \18069 );
xor \U$18768 ( \19111 , \19110 , \18084 );
xor \U$18769 ( \19112 , \19109 , \19111 );
xor \U$18770 ( \19113 , \19070 , \19078 );
and \U$18771 ( \19114 , \19113 , \19087 );
and \U$18772 ( \19115 , \19070 , \19078 );
or \U$18773 ( \19116 , \19114 , \19115 );
xor \U$18774 ( \19117 , \19008 , \19060 );
and \U$18775 ( \19118 , \19117 , \19065 );
and \U$18776 ( \19119 , \19008 , \19060 );
or \U$18777 ( \19120 , \19118 , \19119 );
xor \U$18778 ( \19121 , \19116 , \19120 );
xor \U$18779 ( \19122 , \18400 , \18402 );
xor \U$18780 ( \19123 , \19122 , \18405 );
and \U$18781 ( \19124 , \19095 , \19123 );
xor \U$18782 ( \19125 , \18400 , \18402 );
xor \U$18783 ( \19126 , \19125 , \18405 );
and \U$18784 ( \19127 , \19099 , \19126 );
and \U$18785 ( \19128 , \19095 , \19099 );
or \U$18786 ( \19129 , \19124 , \19127 , \19128 );
xor \U$18787 ( \19130 , \19121 , \19129 );
xor \U$18788 ( \19131 , \18408 , \18410 );
xor \U$18789 ( \19132 , \19131 , \18415 );
xor \U$18790 ( \19133 , \18231 , \18311 );
xor \U$18791 ( \19134 , \19133 , \18394 );
xor \U$18792 ( \19135 , \19132 , \19134 );
xor \U$18793 ( \19136 , \18099 , \18134 );
xor \U$18794 ( \19137 , \19136 , \18147 );
xor \U$18795 ( \19138 , \19135 , \19137 );
and \U$18796 ( \19139 , \19130 , \19138 );
xor \U$18797 ( \19140 , \18059 , \18061 );
xor \U$18798 ( \19141 , \19140 , \18064 );
xor \U$18799 ( \19142 , \18175 , \18202 );
xor \U$18800 ( \19143 , \19142 , \18228 );
and \U$18801 ( \19144 , \18572 , \19143 );
xor \U$18802 ( \19145 , \18175 , \18202 );
xor \U$18803 ( \19146 , \19145 , \18228 );
and \U$18804 ( \19147 , \18574 , \19146 );
and \U$18805 ( \19148 , \18572 , \18574 );
or \U$18806 ( \19149 , \19144 , \19147 , \19148 );
xor \U$18807 ( \19150 , \17672 , \17674 );
xor \U$18808 ( \19151 , \19150 , \17677 );
xor \U$18809 ( \19152 , \18072 , \18079 );
xor \U$18810 ( \19153 , \19151 , \19152 );
xor \U$18811 ( \19154 , \19149 , \19153 );
xor \U$18812 ( \19155 , \19141 , \19154 );
xor \U$18813 ( \19156 , \19132 , \19134 );
xor \U$18814 ( \19157 , \19156 , \19137 );
and \U$18815 ( \19158 , \19155 , \19157 );
and \U$18816 ( \19159 , \19130 , \19155 );
or \U$18817 ( \19160 , \19139 , \19158 , \19159 );
and \U$18818 ( \19161 , \19112 , \19160 );
and \U$18819 ( \19162 , \19109 , \19111 );
or \U$18820 ( \19163 , \19161 , \19162 );
xor \U$18821 ( \19164 , \18437 , \19163 );
xor \U$18822 ( \19165 , \17680 , \17734 );
xor \U$18823 ( \19166 , \19165 , \17747 );
xor \U$18824 ( \19167 , \17833 , \17906 );
xor \U$18825 ( \19168 , \19167 , \17987 );
xor \U$18826 ( \19169 , \18029 , \18031 );
xor \U$18827 ( \19170 , \19169 , \18034 );
xor \U$18828 ( \19171 , \18424 , \18431 );
xor \U$18829 ( \19172 , \19170 , \19171 );
xor \U$18830 ( \19173 , \19168 , \19172 );
xor \U$18831 ( \19174 , \19166 , \19173 );
xor \U$18832 ( \19175 , \18150 , \18397 );
xor \U$18833 ( \19176 , \19175 , \18418 );
xor \U$18834 ( \19177 , \19174 , \19176 );
xor \U$18835 ( \19178 , \18059 , \18061 );
xor \U$18836 ( \19179 , \19178 , \18064 );
and \U$18837 ( \19180 , \19149 , \19179 );
xor \U$18838 ( \19181 , \18059 , \18061 );
xor \U$18839 ( \19182 , \19181 , \18064 );
and \U$18840 ( \19183 , \19153 , \19182 );
and \U$18841 ( \19184 , \19149 , \19153 );
or \U$18842 ( \19185 , \19180 , \19183 , \19184 );
xor \U$18843 ( \19186 , \19116 , \19120 );
and \U$18844 ( \19187 , \19186 , \19129 );
and \U$18845 ( \19188 , \19116 , \19120 );
or \U$18846 ( \19189 , \19187 , \19188 );
xor \U$18847 ( \19190 , \19185 , \19189 );
xor \U$18848 ( \19191 , \19132 , \19134 );
and \U$18849 ( \19192 , \19191 , \19137 );
and \U$18850 ( \19193 , \19132 , \19134 );
or \U$18851 ( \19194 , \19192 , \19193 );
xor \U$18852 ( \19195 , \19190 , \19194 );
and \U$18853 ( \19196 , \19177 , \19195 );
and \U$18854 ( \19197 , \19174 , \19176 );
or \U$18855 ( \19198 , \19196 , \19197 );
and \U$18856 ( \19199 , \19164 , \19198 );
and \U$18857 ( \19200 , \18437 , \19163 );
nor \U$18858 ( \19201 , \19199 , \19200 );
not \U$18859 ( \19202 , \19201 );
xor \U$18860 ( \19203 , \17641 , \17643 );
xor \U$18861 ( \19204 , \19203 , \17650 );
xor \U$18862 ( \19205 , \17198 , \17445 );
xor \U$18863 ( \19206 , \19205 , \17481 );
xor \U$18864 ( \19207 , \19204 , \19206 );
xor \U$18865 ( \19208 , \17670 , \18018 );
xor \U$18866 ( \19209 , \19208 , \18045 );
xor \U$18867 ( \19210 , \19207 , \19209 );
xor \U$18868 ( \19211 , \19185 , \19189 );
and \U$18869 ( \19212 , \19211 , \19194 );
and \U$18870 ( \19213 , \19185 , \19189 );
or \U$18871 ( \19214 , \19212 , \19213 );
xor \U$18872 ( \19215 , \17680 , \17734 );
xor \U$18873 ( \19216 , \19215 , \17747 );
and \U$18874 ( \19217 , \19168 , \19216 );
xor \U$18875 ( \19218 , \17680 , \17734 );
xor \U$18876 ( \19219 , \19218 , \17747 );
and \U$18877 ( \19220 , \19172 , \19219 );
and \U$18878 ( \19221 , \19168 , \19172 );
or \U$18879 ( \19222 , \19217 , \19220 , \19221 );
xor \U$18880 ( \19223 , \19214 , \19222 );
xor \U$18881 ( \19224 , \17662 , \17664 );
xor \U$18882 ( \19225 , \19224 , \17667 );
xor \U$18883 ( \19226 , \17750 , \17990 );
xor \U$18884 ( \19227 , \19226 , \18015 );
xor \U$18885 ( \19228 , \18025 , \18037 );
xor \U$18886 ( \19229 , \19228 , \18042 );
xor \U$18887 ( \19230 , \19227 , \19229 );
xor \U$18888 ( \19231 , \19225 , \19230 );
and \U$18889 ( \19232 , \19223 , \19231 );
and \U$18890 ( \19233 , \19214 , \19222 );
or \U$18891 ( \19234 , \19232 , \19233 );
xor \U$18892 ( \19235 , \18087 , \18421 );
and \U$18893 ( \19236 , \19235 , \18436 );
and \U$18894 ( \19237 , \18087 , \18421 );
or \U$18895 ( \19238 , \19236 , \19237 );
not \U$18896 ( \19239 , \17507 );
xor \U$18897 ( \19240 , \17504 , \17525 );
not \U$18898 ( \19241 , \19240 );
or \U$18899 ( \19242 , \19239 , \19241 );
or \U$18900 ( \19243 , \19240 , \17507 );
nand \U$18901 ( \19244 , \19242 , \19243 );
xor \U$18902 ( \19245 , \19238 , \19244 );
xor \U$18903 ( \19246 , \17662 , \17664 );
xor \U$18904 ( \19247 , \19246 , \17667 );
and \U$18905 ( \19248 , \19227 , \19247 );
xor \U$18906 ( \19249 , \17662 , \17664 );
xor \U$18907 ( \19250 , \19249 , \17667 );
and \U$18908 ( \19251 , \19229 , \19250 );
and \U$18909 ( \19252 , \19227 , \19229 );
or \U$18910 ( \19253 , \19248 , \19251 , \19252 );
xor \U$18911 ( \19254 , \19245 , \19253 );
xor \U$18912 ( \19255 , \19234 , \19254 );
xor \U$18913 ( \19256 , \19210 , \19255 );
not \U$18914 ( \19257 , \19256 );
or \U$18915 ( \19258 , \19202 , \19257 );
or \U$18916 ( \19259 , \19256 , \19201 );
nand \U$18917 ( \19260 , \19258 , \19259 );
xor \U$18918 ( \19261 , \19214 , \19222 );
xor \U$18919 ( \19262 , \19261 , \19231 );
not \U$18920 ( \19263 , \19262 );
xor \U$18921 ( \19264 , \18437 , \19163 );
xor \U$18922 ( \19265 , \19264 , \19198 );
not \U$18923 ( \19266 , \19265 );
or \U$18924 ( \19267 , \19263 , \19266 );
or \U$18925 ( \19268 , \19265 , \19262 );
xor \U$18926 ( \19269 , \18595 , \18842 );
xor \U$18927 ( \19270 , \19269 , \18982 );
xor \U$18928 ( \19271 , \18565 , \18567 );
xor \U$18929 ( \19272 , \19271 , \18576 );
and \U$18930 ( \19273 , \19270 , \19272 );
xor \U$18931 ( \19274 , \19070 , \19078 );
xor \U$18932 ( \19275 , \19274 , \19087 );
xor \U$18933 ( \19276 , \19066 , \19101 );
xor \U$18934 ( \19277 , \19275 , \19276 );
xor \U$18935 ( \19278 , \18565 , \18567 );
xor \U$18936 ( \19279 , \19278 , \18576 );
and \U$18937 ( \19280 , \19277 , \19279 );
and \U$18938 ( \19281 , \19270 , \19277 );
or \U$18939 ( \19282 , \19273 , \19280 , \19281 );
xor \U$18940 ( \19283 , \19012 , \19031 );
xor \U$18941 ( \19284 , \19283 , \19057 );
xor \U$18942 ( \19285 , \18581 , \18583 );
xor \U$18943 ( \19286 , \19285 , \18592 );
and \U$18944 ( \19287 , \19284 , \19286 );
xor \U$18945 ( \19288 , \18520 , \18522 );
xor \U$18946 ( \19289 , \19288 , \18525 );
xor \U$18947 ( \19290 , \18518 , \18560 );
xor \U$18948 ( \19291 , \19289 , \19290 );
xor \U$18949 ( \19292 , \18581 , \18583 );
xor \U$18950 ( \19293 , \19292 , \18592 );
and \U$18951 ( \19294 , \19291 , \19293 );
and \U$18952 ( \19295 , \19284 , \19291 );
or \U$18953 ( \19296 , \19287 , \19294 , \19295 );
and \U$18954 ( \19297 , \1293 , RI98707e0_93);
and \U$18955 ( \19298 , RI986fac0_65, \1291 );
nor \U$18956 ( \19299 , \19297 , \19298 );
not \U$18957 ( \19300 , \19299 );
not \U$18958 ( \19301 , \1128 );
and \U$18959 ( \19302 , \19300 , \19301 );
and \U$18960 ( \19303 , \19299 , \1301 );
nor \U$18961 ( \19304 , \19302 , \19303 );
and \U$18962 ( \19305 , \776 , RI9870600_89);
and \U$18963 ( \19306 , RI98708d0_95, \774 );
nor \U$18964 ( \19307 , \19305 , \19306 );
and \U$18965 ( \19308 , \19307 , \451 );
not \U$18966 ( \19309 , \19307 );
and \U$18967 ( \19310 , \19309 , \474 );
nor \U$18968 ( \19311 , \19308 , \19310 );
xor \U$18969 ( \19312 , \19304 , \19311 );
and \U$18970 ( \19313 , \1329 , RI986fbb0_67);
and \U$18971 ( \19314 , RI986fd90_71, \1327 );
nor \U$18972 ( \19315 , \19313 , \19314 );
and \U$18973 ( \19316 , \19315 , \1337 );
not \U$18974 ( \19317 , \19315 );
and \U$18975 ( \19318 , \19317 , \1336 );
nor \U$18976 ( \19319 , \19316 , \19318 );
and \U$18977 ( \19320 , \19312 , \19319 );
and \U$18978 ( \19321 , \19304 , \19311 );
or \U$18979 ( \19322 , \19320 , \19321 );
and \U$18980 ( \19323 , \2464 , RI9870ab0_99);
and \U$18981 ( \19324 , RI9870d80_105, \2462 );
nor \U$18982 ( \19325 , \19323 , \19324 );
and \U$18983 ( \19326 , \19325 , \2263 );
not \U$18984 ( \19327 , \19325 );
and \U$18985 ( \19328 , \19327 , \2468 );
nor \U$18986 ( \19329 , \19326 , \19328 );
not \U$18987 ( \19330 , \19329 );
and \U$18988 ( \19331 , \3254 , RI98709c0_97);
and \U$18989 ( \19332 , RI9870e70_107, \3252 );
nor \U$18990 ( \19333 , \19331 , \19332 );
not \U$18991 ( \19334 , \19333 );
not \U$18992 ( \19335 , \2935 );
and \U$18993 ( \19336 , \19334 , \19335 );
and \U$18994 ( \19337 , \19333 , \3406 );
nor \U$18995 ( \19338 , \19336 , \19337 );
not \U$18996 ( \19339 , \19338 );
and \U$18997 ( \19340 , \19330 , \19339 );
and \U$18998 ( \19341 , \19338 , \19329 );
and \U$18999 ( \19342 , \3683 , RI9870ba0_101);
and \U$19000 ( \19343 , RI9871050_111, \3681 );
nor \U$19001 ( \19344 , \19342 , \19343 );
not \U$19002 ( \19345 , \19344 );
not \U$19003 ( \19346 , \3918 );
and \U$19004 ( \19347 , \19345 , \19346 );
and \U$19005 ( \19348 , \19344 , \3918 );
nor \U$19006 ( \19349 , \19347 , \19348 );
nor \U$19007 ( \19350 , \19341 , \19349 );
nor \U$19008 ( \19351 , \19340 , \19350 );
or \U$19009 ( \19352 , \19322 , \19351 );
not \U$19010 ( \19353 , \19322 );
not \U$19011 ( \19354 , \19351 );
or \U$19012 ( \19355 , \19353 , \19354 );
and \U$19013 ( \19356 , \1311 , RI986fca0_69);
and \U$19014 ( \19357 , RI986ff70_75, \1309 );
nor \U$19015 ( \19358 , \19356 , \19357 );
and \U$19016 ( \19359 , \19358 , \1315 );
not \U$19017 ( \19360 , \19358 );
and \U$19018 ( \19361 , \19360 , \1458 );
nor \U$19019 ( \19362 , \19359 , \19361 );
and \U$19020 ( \19363 , \2042 , RI986fe80_73);
and \U$19021 ( \19364 , RI9870060_77, \2040 );
nor \U$19022 ( \19365 , \19363 , \19364 );
not \U$19023 ( \19366 , \19365 );
not \U$19024 ( \19367 , \1462 );
and \U$19025 ( \19368 , \19366 , \19367 );
and \U$19026 ( \19369 , \19365 , \1462 );
nor \U$19027 ( \19370 , \19368 , \19369 );
or \U$19028 ( \19371 , \19362 , \19370 );
not \U$19029 ( \19372 , \19370 );
not \U$19030 ( \19373 , \19362 );
or \U$19031 ( \19374 , \19372 , \19373 );
and \U$19032 ( \19375 , \2274 , RI9870150_79);
and \U$19033 ( \19376 , RI9870f60_109, \2272 );
nor \U$19034 ( \19377 , \19375 , \19376 );
and \U$19035 ( \19378 , \19377 , \2030 );
not \U$19036 ( \19379 , \19377 );
and \U$19037 ( \19380 , \19379 , \2031 );
nor \U$19038 ( \19381 , \19378 , \19380 );
nand \U$19039 ( \19382 , \19374 , \19381 );
nand \U$19040 ( \19383 , \19371 , \19382 );
nand \U$19041 ( \19384 , \19355 , \19383 );
nand \U$19042 ( \19385 , \19352 , \19384 );
not \U$19043 ( \19386 , RI9873558_190);
and \U$19044 ( \19387 , \15780 , RI986f610_55);
and \U$19045 ( \19388 , RI9873648_192, RI986df90_7);
nor \U$19046 ( \19389 , \19387 , \19388 );
not \U$19047 ( \19390 , \19389 );
or \U$19048 ( \19391 , \19386 , \19390 );
or \U$19049 ( \19392 , \19389 , RI9873558_190);
nand \U$19050 ( \19393 , \19391 , \19392 );
xor \U$19051 ( \19394 , \19393 , \367 );
and \U$19052 ( \19395 , \14937 , RI986f340_49);
and \U$19053 ( \19396 , RI986f520_53, \14935 );
nor \U$19054 ( \19397 , \19395 , \19396 );
and \U$19055 ( \19398 , \19397 , \14539 );
not \U$19056 ( \19399 , \19397 );
and \U$19057 ( \19400 , \19399 , \14538 );
nor \U$19058 ( \19401 , \19398 , \19400 );
and \U$19059 ( \19402 , \19394 , \19401 );
and \U$19060 ( \19403 , \19393 , \367 );
or \U$19061 ( \19404 , \19402 , \19403 );
not \U$19062 ( \19405 , \19404 );
and \U$19063 ( \19406 , \12293 , RI986e620_21);
and \U$19064 ( \19407 , RI986f7f0_59, \12291 );
nor \U$19065 ( \19408 , \19406 , \19407 );
and \U$19066 ( \19409 , \19408 , \11687 );
not \U$19067 ( \19410 , \19408 );
and \U$19068 ( \19411 , \19410 , \11686 );
nor \U$19069 ( \19412 , \19409 , \19411 );
and \U$19070 ( \19413 , \13045 , RI986f700_57);
and \U$19071 ( \19414 , RI986f9d0_63, \13043 );
nor \U$19072 ( \19415 , \19413 , \19414 );
and \U$19073 ( \19416 , \19415 , \13047 );
not \U$19074 ( \19417 , \19415 );
and \U$19075 ( \19418 , \19417 , \12619 );
nor \U$19076 ( \19419 , \19416 , \19418 );
xor \U$19077 ( \19420 , \19412 , \19419 );
and \U$19078 ( \19421 , \13882 , RI986f8e0_61);
and \U$19079 ( \19422 , RI986f430_51, \13880 );
nor \U$19080 ( \19423 , \19421 , \19422 );
and \U$19081 ( \19424 , \19423 , \13358 );
not \U$19082 ( \19425 , \19423 );
and \U$19083 ( \19426 , \19425 , \13359 );
nor \U$19084 ( \19427 , \19424 , \19426 );
and \U$19085 ( \19428 , \19420 , \19427 );
and \U$19086 ( \19429 , \19412 , \19419 );
or \U$19087 ( \19430 , \19428 , \19429 );
not \U$19088 ( \19431 , \19430 );
or \U$19089 ( \19432 , \19405 , \19431 );
or \U$19090 ( \19433 , \19430 , \19404 );
and \U$19091 ( \19434 , \11696 , RI986e440_17);
and \U$19092 ( \19435 , RI986e710_23, \11694 );
nor \U$19093 ( \19436 , \19434 , \19435 );
and \U$19094 ( \19437 , \19436 , \10965 );
not \U$19095 ( \19438 , \19436 );
and \U$19096 ( \19439 , \19438 , \11702 );
nor \U$19097 ( \19440 , \19437 , \19439 );
and \U$19098 ( \19441 , \9505 , RI986ef80_41);
and \U$19099 ( \19442 , RI986f250_47, \9503 );
nor \U$19100 ( \19443 , \19441 , \19442 );
and \U$19101 ( \19444 , \19443 , \9510 );
not \U$19102 ( \19445 , \19443 );
and \U$19103 ( \19446 , \19445 , \9513 );
nor \U$19104 ( \19447 , \19444 , \19446 );
xor \U$19105 ( \19448 , \19440 , \19447 );
and \U$19106 ( \19449 , \10424 , RI986f160_45);
and \U$19107 ( \19450 , RI986e530_19, \10422 );
nor \U$19108 ( \19451 , \19449 , \19450 );
and \U$19109 ( \19452 , \19451 , \9840 );
not \U$19110 ( \19453 , \19451 );
and \U$19111 ( \19454 , \19453 , \10428 );
nor \U$19112 ( \19455 , \19452 , \19454 );
and \U$19113 ( \19456 , \19448 , \19455 );
and \U$19114 ( \19457 , \19440 , \19447 );
or \U$19115 ( \19458 , \19456 , \19457 );
nand \U$19116 ( \19459 , \19433 , \19458 );
nand \U$19117 ( \19460 , \19432 , \19459 );
xor \U$19118 ( \19461 , \19385 , \19460 );
not \U$19119 ( \19462 , \4521 );
and \U$19120 ( \19463 , \4710 , RI9871140_113);
and \U$19121 ( \19464 , RI9871320_117, \4708 );
nor \U$19122 ( \19465 , \19463 , \19464 );
not \U$19123 ( \19466 , \19465 );
or \U$19124 ( \19467 , \19462 , \19466 );
or \U$19125 ( \19468 , \19465 , \4521 );
nand \U$19126 ( \19469 , \19467 , \19468 );
and \U$19127 ( \19470 , \5318 , RI9871410_119);
and \U$19128 ( \19471 , RI98716e0_125, \5316 );
nor \U$19129 ( \19472 , \19470 , \19471 );
and \U$19130 ( \19473 , \19472 , \5052 );
not \U$19131 ( \19474 , \19472 );
and \U$19132 ( \19475 , \19474 , \5322 );
nor \U$19133 ( \19476 , \19473 , \19475 );
xor \U$19134 ( \19477 , \19469 , \19476 );
and \U$19135 ( \19478 , \4203 , RI9870c90_103);
and \U$19136 ( \19479 , RI9871230_115, \4201 );
nor \U$19137 ( \19480 , \19478 , \19479 );
and \U$19138 ( \19481 , \19480 , \4207 );
not \U$19139 ( \19482 , \19480 );
and \U$19140 ( \19483 , \19482 , \3922 );
nor \U$19141 ( \19484 , \19481 , \19483 );
and \U$19142 ( \19485 , \19477 , \19484 );
and \U$19143 ( \19486 , \19469 , \19476 );
nor \U$19144 ( \19487 , \19485 , \19486 );
and \U$19145 ( \19488 , \8486 , RI986eda0_37);
and \U$19146 ( \19489 , RI986ebc0_33, \8484 );
nor \U$19147 ( \19490 , \19488 , \19489 );
and \U$19148 ( \19491 , \19490 , \8050 );
not \U$19149 ( \19492 , \19490 );
and \U$19150 ( \19493 , \19492 , \8051 );
nor \U$19151 ( \19494 , \19491 , \19493 );
and \U$19152 ( \19495 , \9237 , RI986ecb0_35);
and \U$19153 ( \19496 , RI986f070_43, \9235 );
nor \U$19154 ( \19497 , \19495 , \19496 );
and \U$19155 ( \19498 , \19497 , \9241 );
not \U$19156 ( \19499 , \19497 );
and \U$19157 ( \19500 , \19499 , \8836 );
nor \U$19158 ( \19501 , \19498 , \19500 );
xor \U$19159 ( \19502 , \19494 , \19501 );
and \U$19160 ( \19503 , \7729 , RI986e800_25);
and \U$19161 ( \19504 , RI986ee90_39, \7727 );
nor \U$19162 ( \19505 , \19503 , \19504 );
and \U$19163 ( \19506 , \19505 , \7480 );
not \U$19164 ( \19507 , \19505 );
and \U$19165 ( \19508 , \19507 , \7733 );
nor \U$19166 ( \19509 , \19506 , \19508 );
and \U$19167 ( \19510 , \19502 , \19509 );
and \U$19168 ( \19511 , \19494 , \19501 );
nor \U$19169 ( \19512 , \19510 , \19511 );
xor \U$19170 ( \19513 , \19487 , \19512 );
and \U$19171 ( \19514 , \6453 , RI98715f0_123);
and \U$19172 ( \19515 , RI986ead0_31, \6451 );
nor \U$19173 ( \19516 , \19514 , \19515 );
and \U$19174 ( \19517 , \19516 , \6190 );
not \U$19175 ( \19518 , \19516 );
and \U$19176 ( \19519 , \19518 , \6180 );
nor \U$19177 ( \19520 , \19517 , \19519 );
and \U$19178 ( \19521 , \7079 , RI986e9e0_29);
and \U$19179 ( \19522 , RI986e8f0_27, \7077 );
nor \U$19180 ( \19523 , \19521 , \19522 );
and \U$19181 ( \19524 , \19523 , \6710 );
not \U$19182 ( \19525 , \19523 );
and \U$19183 ( \19526 , \19525 , \6709 );
nor \U$19184 ( \19527 , \19524 , \19526 );
xor \U$19185 ( \19528 , \19520 , \19527 );
and \U$19186 ( \19529 , \5881 , RI98717d0_127);
and \U$19187 ( \19530 , RI9871500_121, \5879 );
nor \U$19188 ( \19531 , \19529 , \19530 );
and \U$19189 ( \19532 , \19531 , \5594 );
not \U$19190 ( \19533 , \19531 );
and \U$19191 ( \19534 , \19533 , \5885 );
nor \U$19192 ( \19535 , \19532 , \19534 );
and \U$19193 ( \19536 , \19528 , \19535 );
and \U$19194 ( \19537 , \19520 , \19527 );
nor \U$19195 ( \19538 , \19536 , \19537 );
and \U$19196 ( \19539 , \19513 , \19538 );
and \U$19197 ( \19540 , \19487 , \19512 );
nor \U$19198 ( \19541 , \19539 , \19540 );
and \U$19199 ( \19542 , \19461 , \19541 );
and \U$19200 ( \19543 , \19385 , \19460 );
or \U$19201 ( \19544 , \19542 , \19543 );
xor \U$19202 ( \19545 , \19039 , \19046 );
xor \U$19203 ( \19546 , \19545 , \19054 );
xor \U$19204 ( \19547 , \19020 , \487 );
xor \U$19205 ( \19548 , \19547 , \19028 );
and \U$19206 ( \19549 , \19546 , \19548 );
xor \U$19207 ( \19550 , \18683 , \18690 );
xor \U$19208 ( \19551 , \19550 , \18698 );
xor \U$19209 ( \19552 , \18708 , \18716 );
xor \U$19210 ( \19553 , \19552 , \18724 );
xor \U$19211 ( \19554 , \19551 , \19553 );
xor \U$19212 ( \19555 , \18735 , \18742 );
xor \U$19213 ( \19556 , \19555 , \18750 );
and \U$19214 ( \19557 , \19554 , \19556 );
and \U$19215 ( \19558 , \19551 , \19553 );
or \U$19216 ( \19559 , \19557 , \19558 );
xor \U$19217 ( \19560 , \19020 , \487 );
xor \U$19218 ( \19561 , \19560 , \19028 );
and \U$19219 ( \19562 , \19559 , \19561 );
and \U$19220 ( \19563 , \19546 , \19559 );
or \U$19221 ( \19564 , \19549 , \19562 , \19563 );
xor \U$19222 ( \19565 , \19544 , \19564 );
xor \U$19223 ( \19566 , \18628 , \18635 );
xor \U$19224 ( \19567 , \19566 , \18644 );
xor \U$19225 ( \19568 , \18602 , \18609 );
xor \U$19226 ( \19569 , \19568 , \18617 );
and \U$19227 ( \19570 , \19567 , \19569 );
xor \U$19228 ( \19571 , \18655 , \18662 );
xor \U$19229 ( \19572 , \19571 , \18670 );
xor \U$19230 ( \19573 , \18602 , \18609 );
xor \U$19231 ( \19574 , \19573 , \18617 );
and \U$19232 ( \19575 , \19572 , \19574 );
and \U$19233 ( \19576 , \19567 , \19572 );
or \U$19234 ( \19577 , \19570 , \19575 , \19576 );
not \U$19235 ( \19578 , \367 );
and \U$19236 ( \19579 , \376 , RI9870420_85);
and \U$19237 ( \19580 , RI9870510_87, \374 );
nor \U$19238 ( \19581 , \19579 , \19580 );
not \U$19239 ( \19582 , \19581 );
or \U$19240 ( \19583 , \19578 , \19582 );
or \U$19241 ( \19584 , \19581 , \367 );
nand \U$19242 ( \19585 , \19583 , \19584 );
not \U$19243 ( \19586 , \456 );
and \U$19244 ( \19587 , \465 , RI9870330_83);
and \U$19245 ( \19588 , RI9870240_81, \463 );
nor \U$19246 ( \19589 , \19587 , \19588 );
not \U$19247 ( \19590 , \19589 );
or \U$19248 ( \19591 , \19586 , \19590 );
or \U$19249 ( \19592 , \19589 , \454 );
nand \U$19250 ( \19593 , \19591 , \19592 );
xor \U$19251 ( \19594 , \19585 , \19593 );
and \U$19252 ( \19595 , \438 , RI9870240_81);
and \U$19253 ( \19596 , RI98706f0_91, \436 );
nor \U$19254 ( \19597 , \19595 , \19596 );
and \U$19255 ( \19598 , \19597 , \444 );
not \U$19256 ( \19599 , \19597 );
and \U$19257 ( \19600 , \19599 , \443 );
nor \U$19258 ( \19601 , \19598 , \19600 );
nand \U$19259 ( \19602 , RI9870420_85, \374 );
not \U$19260 ( \19603 , \19602 );
not \U$19261 ( \19604 , \367 );
or \U$19262 ( \19605 , \19603 , \19604 );
or \U$19263 ( \19606 , \365 , \19602 );
nand \U$19264 ( \19607 , \19605 , \19606 );
xor \U$19265 ( \19608 , \19601 , \19607 );
not \U$19266 ( \19609 , \456 );
and \U$19267 ( \19610 , \465 , RI9870510_87);
and \U$19268 ( \19611 , RI9870330_83, \463 );
nor \U$19269 ( \19612 , \19610 , \19611 );
not \U$19270 ( \19613 , \19612 );
or \U$19271 ( \19614 , \19609 , \19613 );
or \U$19272 ( \19615 , \19612 , \454 );
nand \U$19273 ( \19616 , \19614 , \19615 );
and \U$19274 ( \19617 , \19608 , \19616 );
and \U$19275 ( \19618 , \19601 , \19607 );
or \U$19276 ( \19619 , \19617 , \19618 );
and \U$19277 ( \19620 , \19594 , \19619 );
and \U$19278 ( \19621 , \19585 , \19593 );
or \U$19279 ( \19622 , \19620 , \19621 );
xor \U$19280 ( \19623 , \19577 , \19622 );
xor \U$19281 ( \19624 , \18764 , \18771 );
xor \U$19282 ( \19625 , \19624 , \18780 );
xor \U$19283 ( \19626 , \18791 , \18798 );
xor \U$19284 ( \19627 , \19626 , \18806 );
and \U$19285 ( \19628 , \19625 , \19627 );
xor \U$19286 ( \19629 , \18818 , \18825 );
xor \U$19287 ( \19630 , \19629 , \18833 );
xor \U$19288 ( \19631 , \18791 , \18798 );
xor \U$19289 ( \19632 , \19631 , \18806 );
and \U$19290 ( \19633 , \19630 , \19632 );
and \U$19291 ( \19634 , \19625 , \19630 );
or \U$19292 ( \19635 , \19628 , \19633 , \19634 );
and \U$19293 ( \19636 , \19623 , \19635 );
and \U$19294 ( \19637 , \19577 , \19622 );
or \U$19295 ( \19638 , \19636 , \19637 );
and \U$19296 ( \19639 , \19565 , \19638 );
and \U$19297 ( \19640 , \19544 , \19564 );
or \U$19298 ( \19641 , \19639 , \19640 );
xor \U$19299 ( \19642 , \19296 , \19641 );
xor \U$19300 ( \19643 , \18620 , \18647 );
xor \U$19301 ( \19644 , \19643 , \18673 );
xor \U$19302 ( \19645 , \18783 , \18809 );
xor \U$19303 ( \19646 , \19645 , \18836 );
and \U$19304 ( \19647 , \19644 , \19646 );
xor \U$19305 ( \19648 , \18701 , \18727 );
xor \U$19306 ( \19649 , \19648 , \18753 );
xor \U$19307 ( \19650 , \18783 , \18809 );
xor \U$19308 ( \19651 , \19650 , \18836 );
and \U$19309 ( \19652 , \19649 , \19651 );
and \U$19310 ( \19653 , \19644 , \19649 );
or \U$19311 ( \19654 , \19647 , \19652 , \19653 );
not \U$19312 ( \19655 , \19654 );
xor \U$19313 ( \19656 , \18992 , \18998 );
xor \U$19314 ( \19657 , \19656 , \19005 );
or \U$19315 ( \19658 , \19655 , \19657 );
not \U$19316 ( \19659 , \19657 );
not \U$19317 ( \19660 , \19655 );
or \U$19318 ( \19661 , \19659 , \19660 );
xor \U$19319 ( \19662 , \18445 , \18452 );
xor \U$19320 ( \19663 , \19662 , \18461 );
xor \U$19321 ( \19664 , \18943 , \18974 );
xor \U$19322 ( \19665 , \19663 , \19664 );
xor \U$19323 ( \19666 , \18928 , \18934 );
xor \U$19324 ( \19667 , \19666 , \18937 );
and \U$19325 ( \19668 , \19665 , \19667 );
xor \U$19326 ( \19669 , \18877 , \18884 );
xor \U$19327 ( \19670 , \19669 , \18892 );
xor \U$19328 ( \19671 , \18870 , \18921 );
xor \U$19329 ( \19672 , \19670 , \19671 );
xor \U$19330 ( \19673 , \18928 , \18934 );
xor \U$19331 ( \19674 , \19673 , \18937 );
and \U$19332 ( \19675 , \19672 , \19674 );
and \U$19333 ( \19676 , \19665 , \19672 );
or \U$19334 ( \19677 , \19668 , \19675 , \19676 );
nand \U$19335 ( \19678 , \19661 , \19677 );
nand \U$19336 ( \19679 , \19658 , \19678 );
and \U$19337 ( \19680 , \19642 , \19679 );
and \U$19338 ( \19681 , \19296 , \19641 );
or \U$19339 ( \19682 , \19680 , \19681 );
xor \U$19340 ( \19683 , \19282 , \19682 );
xor \U$19341 ( \19684 , \19132 , \19134 );
xor \U$19342 ( \19685 , \19684 , \19137 );
xor \U$19343 ( \19686 , \19130 , \19155 );
xor \U$19344 ( \19687 , \19685 , \19686 );
and \U$19345 ( \19688 , \19683 , \19687 );
and \U$19346 ( \19689 , \19282 , \19682 );
or \U$19347 ( \19690 , \19688 , \19689 );
xor \U$19348 ( \19691 , \19174 , \19176 );
xor \U$19349 ( \19692 , \19691 , \19195 );
and \U$19350 ( \19693 , \19690 , \19692 );
xor \U$19351 ( \19694 , \19109 , \19111 );
xor \U$19352 ( \19695 , \19694 , \19160 );
xor \U$19353 ( \19696 , \19174 , \19176 );
xor \U$19354 ( \19697 , \19696 , \19195 );
and \U$19355 ( \19698 , \19695 , \19697 );
and \U$19356 ( \19699 , \19690 , \19695 );
or \U$19357 ( \19700 , \19693 , \19698 , \19699 );
nand \U$19358 ( \19701 , \19268 , \19700 );
nand \U$19359 ( \19702 , \19267 , \19701 );
and \U$19360 ( \19703 , \19260 , \19702 );
xor \U$19361 ( \19704 , \19702 , \19260 );
xnor \U$19362 ( \19705 , \19265 , \19700 );
not \U$19363 ( \19706 , \19705 );
not \U$19364 ( \19707 , \19262 );
and \U$19365 ( \19708 , \19706 , \19707 );
and \U$19366 ( \19709 , \19705 , \19262 );
nor \U$19367 ( \19710 , \19708 , \19709 );
xor \U$19368 ( \19711 , \19282 , \19682 );
xor \U$19369 ( \19712 , \19711 , \19687 );
xor \U$19370 ( \19713 , \18579 , \18985 );
xor \U$19371 ( \19714 , \19713 , \19106 );
xor \U$19372 ( \19715 , \19712 , \19714 );
xor \U$19373 ( \19716 , \19520 , \19527 );
xor \U$19374 ( \19717 , \19716 , \19535 );
not \U$19375 ( \19718 , \19329 );
xor \U$19376 ( \19719 , \19338 , \19349 );
not \U$19377 ( \19720 , \19719 );
or \U$19378 ( \19721 , \19718 , \19720 );
or \U$19379 ( \19722 , \19719 , \19329 );
nand \U$19380 ( \19723 , \19721 , \19722 );
xor \U$19381 ( \19724 , \19717 , \19723 );
xor \U$19382 ( \19725 , \19469 , \19476 );
xor \U$19383 ( \19726 , \19725 , \19484 );
and \U$19384 ( \19727 , \19724 , \19726 );
and \U$19385 ( \19728 , \19717 , \19723 );
or \U$19386 ( \19729 , \19727 , \19728 );
xor \U$19387 ( \19730 , \19304 , \19311 );
xor \U$19388 ( \19731 , \19730 , \19319 );
not \U$19389 ( \19732 , \19370 );
not \U$19390 ( \19733 , \19381 );
or \U$19391 ( \19734 , \19732 , \19733 );
or \U$19392 ( \19735 , \19370 , \19381 );
nand \U$19393 ( \19736 , \19734 , \19735 );
not \U$19394 ( \19737 , \19736 );
not \U$19395 ( \19738 , \19362 );
and \U$19396 ( \19739 , \19737 , \19738 );
and \U$19397 ( \19740 , \19736 , \19362 );
nor \U$19398 ( \19741 , \19739 , \19740 );
or \U$19399 ( \19742 , \19731 , \19741 );
not \U$19400 ( \19743 , \19741 );
not \U$19401 ( \19744 , \19731 );
or \U$19402 ( \19745 , \19743 , \19744 );
xor \U$19403 ( \19746 , \19601 , \19607 );
xor \U$19404 ( \19747 , \19746 , \19616 );
nand \U$19405 ( \19748 , \19745 , \19747 );
nand \U$19406 ( \19749 , \19742 , \19748 );
xor \U$19407 ( \19750 , \19729 , \19749 );
xor \U$19408 ( \19751 , \19412 , \19419 );
xor \U$19409 ( \19752 , \19751 , \19427 );
xor \U$19410 ( \19753 , \19494 , \19501 );
xor \U$19411 ( \19754 , \19753 , \19509 );
xor \U$19412 ( \19755 , \19752 , \19754 );
xor \U$19413 ( \19756 , \19440 , \19447 );
xor \U$19414 ( \19757 , \19756 , \19455 );
and \U$19415 ( \19758 , \19755 , \19757 );
and \U$19416 ( \19759 , \19752 , \19754 );
or \U$19417 ( \19760 , \19758 , \19759 );
and \U$19418 ( \19761 , \19750 , \19760 );
and \U$19419 ( \19762 , \19729 , \19749 );
or \U$19420 ( \19763 , \19761 , \19762 );
and \U$19421 ( \19764 , \2042 , RI986ff70_75);
and \U$19422 ( \19765 , RI986fe80_73, \2040 );
nor \U$19423 ( \19766 , \19764 , \19765 );
not \U$19424 ( \19767 , \19766 );
not \U$19425 ( \19768 , \1462 );
and \U$19426 ( \19769 , \19767 , \19768 );
and \U$19427 ( \19770 , \19766 , \1462 );
nor \U$19428 ( \19771 , \19769 , \19770 );
and \U$19429 ( \19772 , \1329 , RI986fac0_65);
and \U$19430 ( \19773 , RI986fbb0_67, \1327 );
nor \U$19431 ( \19774 , \19772 , \19773 );
and \U$19432 ( \19775 , \19774 , \1337 );
not \U$19433 ( \19776 , \19774 );
and \U$19434 ( \19777 , \19776 , \1336 );
nor \U$19435 ( \19778 , \19775 , \19777 );
xor \U$19436 ( \19779 , \19771 , \19778 );
and \U$19437 ( \19780 , \1311 , RI986fd90_71);
and \U$19438 ( \19781 , RI986fca0_69, \1309 );
nor \U$19439 ( \19782 , \19780 , \19781 );
and \U$19440 ( \19783 , \19782 , \1315 );
not \U$19441 ( \19784 , \19782 );
and \U$19442 ( \19785 , \19784 , \1319 );
nor \U$19443 ( \19786 , \19783 , \19785 );
and \U$19444 ( \19787 , \19779 , \19786 );
and \U$19445 ( \19788 , \19771 , \19778 );
or \U$19446 ( \19789 , \19787 , \19788 );
and \U$19447 ( \19790 , \3254 , RI9870d80_105);
and \U$19448 ( \19791 , RI98709c0_97, \3252 );
nor \U$19449 ( \19792 , \19790 , \19791 );
not \U$19450 ( \19793 , \19792 );
not \U$19451 ( \19794 , \2935 );
and \U$19452 ( \19795 , \19793 , \19794 );
and \U$19453 ( \19796 , \19792 , \3406 );
nor \U$19454 ( \19797 , \19795 , \19796 );
and \U$19455 ( \19798 , \2274 , RI9870060_77);
and \U$19456 ( \19799 , RI9870150_79, \2272 );
nor \U$19457 ( \19800 , \19798 , \19799 );
and \U$19458 ( \19801 , \19800 , \2031 );
not \U$19459 ( \19802 , \19800 );
and \U$19460 ( \19803 , \19802 , \2030 );
nor \U$19461 ( \19804 , \19801 , \19803 );
xor \U$19462 ( \19805 , \19797 , \19804 );
and \U$19463 ( \19806 , \2464 , RI9870f60_109);
and \U$19464 ( \19807 , RI9870ab0_99, \2462 );
nor \U$19465 ( \19808 , \19806 , \19807 );
and \U$19466 ( \19809 , \19808 , \2263 );
not \U$19467 ( \19810 , \19808 );
and \U$19468 ( \19811 , \19810 , \2468 );
nor \U$19469 ( \19812 , \19809 , \19811 );
and \U$19470 ( \19813 , \19805 , \19812 );
and \U$19471 ( \19814 , \19797 , \19804 );
or \U$19472 ( \19815 , \19813 , \19814 );
or \U$19473 ( \19816 , \19789 , \19815 );
not \U$19474 ( \19817 , \19789 );
not \U$19475 ( \19818 , \19815 );
or \U$19476 ( \19819 , \19817 , \19818 );
not \U$19477 ( \19820 , \1128 );
and \U$19478 ( \19821 , \1293 , RI98708d0_95);
and \U$19479 ( \19822 , RI98707e0_93, \1291 );
nor \U$19480 ( \19823 , \19821 , \19822 );
not \U$19481 ( \19824 , \19823 );
or \U$19482 ( \19825 , \19820 , \19824 );
or \U$19483 ( \19826 , \19823 , \1301 );
nand \U$19484 ( \19827 , \19825 , \19826 );
and \U$19485 ( \19828 , \776 , RI98706f0_91);
and \U$19486 ( \19829 , RI9870600_89, \774 );
nor \U$19487 ( \19830 , \19828 , \19829 );
and \U$19488 ( \19831 , \19830 , \474 );
not \U$19489 ( \19832 , \19830 );
and \U$19490 ( \19833 , \19832 , \451 );
nor \U$19491 ( \19834 , \19831 , \19833 );
xor \U$19492 ( \19835 , \19827 , \19834 );
and \U$19493 ( \19836 , \438 , RI9870330_83);
and \U$19494 ( \19837 , RI9870240_81, \436 );
nor \U$19495 ( \19838 , \19836 , \19837 );
and \U$19496 ( \19839 , \19838 , \444 );
not \U$19497 ( \19840 , \19838 );
and \U$19498 ( \19841 , \19840 , \443 );
nor \U$19499 ( \19842 , \19839 , \19841 );
and \U$19500 ( \19843 , \19835 , \19842 );
and \U$19501 ( \19844 , \19827 , \19834 );
or \U$19502 ( \19845 , \19843 , \19844 );
nand \U$19503 ( \19846 , \19819 , \19845 );
nand \U$19504 ( \19847 , \19816 , \19846 );
and \U$19505 ( \19848 , \14937 , RI986f430_51);
and \U$19506 ( \19849 , RI986f340_49, \14935 );
nor \U$19507 ( \19850 , \19848 , \19849 );
and \U$19508 ( \19851 , \19850 , \14538 );
not \U$19509 ( \19852 , \19850 );
and \U$19510 ( \19853 , \19852 , \14539 );
nor \U$19511 ( \19854 , \19851 , \19853 );
and \U$19512 ( \19855 , \15780 , RI986f520_53);
and \U$19513 ( \19856 , RI9873648_192, RI986f610_55);
nor \U$19514 ( \19857 , \19855 , \19856 );
not \U$19515 ( \19858 , \19857 );
not \U$19516 ( \19859 , RI9873558_190);
and \U$19517 ( \19860 , \19858 , \19859 );
and \U$19518 ( \19861 , \19857 , RI9873558_190);
nor \U$19519 ( \19862 , \19860 , \19861 );
xor \U$19520 ( \19863 , \19854 , \19862 );
and \U$19521 ( \19864 , \13882 , RI986f9d0_63);
and \U$19522 ( \19865 , RI986f8e0_61, \13880 );
nor \U$19523 ( \19866 , \19864 , \19865 );
and \U$19524 ( \19867 , \19866 , \13359 );
not \U$19525 ( \19868 , \19866 );
and \U$19526 ( \19869 , \19868 , \13358 );
nor \U$19527 ( \19870 , \19867 , \19869 );
and \U$19528 ( \19871 , \19863 , \19870 );
and \U$19529 ( \19872 , \19854 , \19862 );
or \U$19530 ( \19873 , \19871 , \19872 );
and \U$19531 ( \19874 , \9505 , RI986f070_43);
and \U$19532 ( \19875 , RI986ef80_41, \9503 );
nor \U$19533 ( \19876 , \19874 , \19875 );
and \U$19534 ( \19877 , \19876 , \9513 );
not \U$19535 ( \19878 , \19876 );
and \U$19536 ( \19879 , \19878 , \9510 );
nor \U$19537 ( \19880 , \19877 , \19879 );
and \U$19538 ( \19881 , \9237 , RI986ebc0_33);
and \U$19539 ( \19882 , RI986ecb0_35, \9235 );
nor \U$19540 ( \19883 , \19881 , \19882 );
and \U$19541 ( \19884 , \19883 , \8836 );
not \U$19542 ( \19885 , \19883 );
and \U$19543 ( \19886 , \19885 , \9241 );
nor \U$19544 ( \19887 , \19884 , \19886 );
xor \U$19545 ( \19888 , \19880 , \19887 );
and \U$19546 ( \19889 , \10424 , RI986f250_47);
and \U$19547 ( \19890 , RI986f160_45, \10422 );
nor \U$19548 ( \19891 , \19889 , \19890 );
and \U$19549 ( \19892 , \19891 , \10428 );
not \U$19550 ( \19893 , \19891 );
and \U$19551 ( \19894 , \19893 , \9840 );
nor \U$19552 ( \19895 , \19892 , \19894 );
and \U$19553 ( \19896 , \19888 , \19895 );
and \U$19554 ( \19897 , \19880 , \19887 );
or \U$19555 ( \19898 , \19896 , \19897 );
xor \U$19556 ( \19899 , \19873 , \19898 );
and \U$19557 ( \19900 , \12293 , RI986e710_23);
and \U$19558 ( \19901 , RI986e620_21, \12291 );
nor \U$19559 ( \19902 , \19900 , \19901 );
and \U$19560 ( \19903 , \19902 , \11686 );
not \U$19561 ( \19904 , \19902 );
and \U$19562 ( \19905 , \19904 , \11687 );
nor \U$19563 ( \19906 , \19903 , \19905 );
and \U$19564 ( \19907 , \11696 , RI986e530_19);
and \U$19565 ( \19908 , RI986e440_17, \11694 );
nor \U$19566 ( \19909 , \19907 , \19908 );
and \U$19567 ( \19910 , \19909 , \11702 );
not \U$19568 ( \19911 , \19909 );
and \U$19569 ( \19912 , \19911 , \10965 );
nor \U$19570 ( \19913 , \19910 , \19912 );
xor \U$19571 ( \19914 , \19906 , \19913 );
and \U$19572 ( \19915 , \13045 , RI986f7f0_59);
and \U$19573 ( \19916 , RI986f700_57, \13043 );
nor \U$19574 ( \19917 , \19915 , \19916 );
and \U$19575 ( \19918 , \19917 , \12619 );
not \U$19576 ( \19919 , \19917 );
and \U$19577 ( \19920 , \19919 , \13047 );
nor \U$19578 ( \19921 , \19918 , \19920 );
and \U$19579 ( \19922 , \19914 , \19921 );
and \U$19580 ( \19923 , \19906 , \19913 );
or \U$19581 ( \19924 , \19922 , \19923 );
and \U$19582 ( \19925 , \19899 , \19924 );
and \U$19583 ( \19926 , \19873 , \19898 );
nor \U$19584 ( \19927 , \19925 , \19926 );
xor \U$19585 ( \19928 , \19847 , \19927 );
and \U$19586 ( \19929 , \4710 , RI9871230_115);
and \U$19587 ( \19930 , RI9871140_113, \4708 );
nor \U$19588 ( \19931 , \19929 , \19930 );
not \U$19589 ( \19932 , \19931 );
not \U$19590 ( \19933 , \4519 );
and \U$19591 ( \19934 , \19932 , \19933 );
and \U$19592 ( \19935 , \19931 , \4521 );
nor \U$19593 ( \19936 , \19934 , \19935 );
and \U$19594 ( \19937 , \3683 , RI9870e70_107);
and \U$19595 ( \19938 , RI9870ba0_101, \3681 );
nor \U$19596 ( \19939 , \19937 , \19938 );
not \U$19597 ( \19940 , \19939 );
not \U$19598 ( \19941 , \3412 );
and \U$19599 ( \19942 , \19940 , \19941 );
and \U$19600 ( \19943 , \19939 , \3412 );
nor \U$19601 ( \19944 , \19942 , \19943 );
xor \U$19602 ( \19945 , \19936 , \19944 );
and \U$19603 ( \19946 , \4203 , RI9871050_111);
and \U$19604 ( \19947 , RI9870c90_103, \4201 );
nor \U$19605 ( \19948 , \19946 , \19947 );
and \U$19606 ( \19949 , \19948 , \3922 );
not \U$19607 ( \19950 , \19948 );
and \U$19608 ( \19951 , \19950 , \4207 );
nor \U$19609 ( \19952 , \19949 , \19951 );
and \U$19610 ( \19953 , \19945 , \19952 );
and \U$19611 ( \19954 , \19936 , \19944 );
or \U$19612 ( \19955 , \19953 , \19954 );
and \U$19613 ( \19956 , \7079 , RI986ead0_31);
and \U$19614 ( \19957 , RI986e9e0_29, \7077 );
nor \U$19615 ( \19958 , \19956 , \19957 );
and \U$19616 ( \19959 , \19958 , \6709 );
not \U$19617 ( \19960 , \19958 );
and \U$19618 ( \19961 , \19960 , \6710 );
nor \U$19619 ( \19962 , \19959 , \19961 );
not \U$19620 ( \19963 , \19962 );
and \U$19621 ( \19964 , \8486 , RI986ee90_39);
and \U$19622 ( \19965 , RI986eda0_37, \8484 );
nor \U$19623 ( \19966 , \19964 , \19965 );
and \U$19624 ( \19967 , \19966 , \8051 );
not \U$19625 ( \19968 , \19966 );
and \U$19626 ( \19969 , \19968 , \8050 );
nor \U$19627 ( \19970 , \19967 , \19969 );
not \U$19628 ( \19971 , \19970 );
and \U$19629 ( \19972 , \19963 , \19971 );
and \U$19630 ( \19973 , \19970 , \19962 );
and \U$19631 ( \19974 , \7729 , RI986e8f0_27);
and \U$19632 ( \19975 , RI986e800_25, \7727 );
nor \U$19633 ( \19976 , \19974 , \19975 );
and \U$19634 ( \19977 , \19976 , \7733 );
not \U$19635 ( \19978 , \19976 );
and \U$19636 ( \19979 , \19978 , \7480 );
nor \U$19637 ( \19980 , \19977 , \19979 );
nor \U$19638 ( \19981 , \19973 , \19980 );
nor \U$19639 ( \19982 , \19972 , \19981 );
xor \U$19640 ( \19983 , \19955 , \19982 );
and \U$19641 ( \19984 , \5881 , RI98716e0_125);
and \U$19642 ( \19985 , RI98717d0_127, \5879 );
nor \U$19643 ( \19986 , \19984 , \19985 );
and \U$19644 ( \19987 , \19986 , \5594 );
not \U$19645 ( \19988 , \19986 );
and \U$19646 ( \19989 , \19988 , \5885 );
nor \U$19647 ( \19990 , \19987 , \19989 );
and \U$19648 ( \19991 , \6453 , RI9871500_121);
and \U$19649 ( \19992 , RI98715f0_123, \6451 );
nor \U$19650 ( \19993 , \19991 , \19992 );
and \U$19651 ( \19994 , \19993 , \6190 );
not \U$19652 ( \19995 , \19993 );
and \U$19653 ( \19996 , \19995 , \6180 );
nor \U$19654 ( \19997 , \19994 , \19996 );
xor \U$19655 ( \19998 , \19990 , \19997 );
and \U$19656 ( \19999 , \5318 , RI9871320_117);
and \U$19657 ( \20000 , RI9871410_119, \5316 );
nor \U$19658 ( \20001 , \19999 , \20000 );
and \U$19659 ( \20002 , \20001 , \5052 );
not \U$19660 ( \20003 , \20001 );
and \U$19661 ( \20004 , \20003 , \5322 );
nor \U$19662 ( \20005 , \20002 , \20004 );
and \U$19663 ( \20006 , \19998 , \20005 );
and \U$19664 ( \20007 , \19990 , \19997 );
nor \U$19665 ( \20008 , \20006 , \20007 );
and \U$19666 ( \20009 , \19983 , \20008 );
and \U$19667 ( \20010 , \19955 , \19982 );
nor \U$19668 ( \20011 , \20009 , \20010 );
and \U$19669 ( \20012 , \19928 , \20011 );
and \U$19670 ( \20013 , \19847 , \19927 );
or \U$19671 ( \20014 , \20012 , \20013 );
xor \U$19672 ( \20015 , \19763 , \20014 );
xor \U$19673 ( \20016 , \18602 , \18609 );
xor \U$19674 ( \20017 , \20016 , \18617 );
xor \U$19675 ( \20018 , \19567 , \19572 );
xor \U$19676 ( \20019 , \20017 , \20018 );
xor \U$19677 ( \20020 , \19551 , \19553 );
xor \U$19678 ( \20021 , \20020 , \19556 );
and \U$19679 ( \20022 , \20019 , \20021 );
xor \U$19680 ( \20023 , \18791 , \18798 );
xor \U$19681 ( \20024 , \20023 , \18806 );
xor \U$19682 ( \20025 , \19625 , \19630 );
xor \U$19683 ( \20026 , \20024 , \20025 );
xor \U$19684 ( \20027 , \19551 , \19553 );
xor \U$19685 ( \20028 , \20027 , \19556 );
and \U$19686 ( \20029 , \20026 , \20028 );
and \U$19687 ( \20030 , \20019 , \20026 );
or \U$19688 ( \20031 , \20022 , \20029 , \20030 );
and \U$19689 ( \20032 , \20015 , \20031 );
and \U$19690 ( \20033 , \19763 , \20014 );
or \U$19691 ( \20034 , \20032 , \20033 );
xor \U$19692 ( \20035 , \19020 , \487 );
xor \U$19693 ( \20036 , \20035 , \19028 );
xor \U$19694 ( \20037 , \19546 , \19559 );
xor \U$19695 ( \20038 , \20036 , \20037 );
xor \U$19696 ( \20039 , \19385 , \19460 );
xor \U$19697 ( \20040 , \20039 , \19541 );
xor \U$19698 ( \20041 , \20038 , \20040 );
xor \U$19699 ( \20042 , \19577 , \19622 );
xor \U$19700 ( \20043 , \20042 , \19635 );
and \U$19701 ( \20044 , \20041 , \20043 );
and \U$19702 ( \20045 , \20038 , \20040 );
or \U$19703 ( \20046 , \20044 , \20045 );
xor \U$19704 ( \20047 , \20034 , \20046 );
xor \U$19705 ( \20048 , \18783 , \18809 );
xor \U$19706 ( \20049 , \20048 , \18836 );
xor \U$19707 ( \20050 , \19644 , \19649 );
xor \U$19708 ( \20051 , \20049 , \20050 );
not \U$19709 ( \20052 , \19383 );
not \U$19710 ( \20053 , \19322 );
or \U$19711 ( \20054 , \20052 , \20053 );
or \U$19712 ( \20055 , \19322 , \19383 );
nand \U$19713 ( \20056 , \20054 , \20055 );
not \U$19714 ( \20057 , \20056 );
not \U$19715 ( \20058 , \19351 );
and \U$19716 ( \20059 , \20057 , \20058 );
and \U$19717 ( \20060 , \20056 , \19351 );
nor \U$19718 ( \20061 , \20059 , \20060 );
xor \U$19719 ( \20062 , \19487 , \19512 );
xor \U$19720 ( \20063 , \20062 , \19538 );
or \U$19721 ( \20064 , \20061 , \20063 );
not \U$19722 ( \20065 , \20063 );
not \U$19723 ( \20066 , \20061 );
or \U$19724 ( \20067 , \20065 , \20066 );
xor \U$19725 ( \20068 , \19585 , \19593 );
xor \U$19726 ( \20069 , \20068 , \19619 );
nand \U$19727 ( \20070 , \20067 , \20069 );
nand \U$19728 ( \20071 , \20064 , \20070 );
xor \U$19729 ( \20072 , \20051 , \20071 );
xor \U$19730 ( \20073 , \18928 , \18934 );
xor \U$19731 ( \20074 , \20073 , \18937 );
xor \U$19732 ( \20075 , \19665 , \19672 );
xor \U$19733 ( \20076 , \20074 , \20075 );
and \U$19734 ( \20077 , \20072 , \20076 );
and \U$19735 ( \20078 , \20051 , \20071 );
or \U$19736 ( \20079 , \20077 , \20078 );
and \U$19737 ( \20080 , \20047 , \20079 );
and \U$19738 ( \20081 , \20034 , \20046 );
or \U$19739 ( \20082 , \20080 , \20081 );
xor \U$19740 ( \20083 , \18926 , \18940 );
xor \U$19741 ( \20084 , \20083 , \18979 );
xor \U$19742 ( \20085 , \18676 , \18756 );
xor \U$19743 ( \20086 , \20085 , \18839 );
xor \U$19744 ( \20087 , \20084 , \20086 );
xor \U$19745 ( \20088 , \18581 , \18583 );
xor \U$19746 ( \20089 , \20088 , \18592 );
xor \U$19747 ( \20090 , \19284 , \19291 );
xor \U$19748 ( \20091 , \20089 , \20090 );
and \U$19749 ( \20092 , \20087 , \20091 );
and \U$19750 ( \20093 , \20084 , \20086 );
or \U$19751 ( \20094 , \20092 , \20093 );
xor \U$19752 ( \20095 , \20082 , \20094 );
xor \U$19753 ( \20096 , \18565 , \18567 );
xor \U$19754 ( \20097 , \20096 , \18576 );
xor \U$19755 ( \20098 , \19270 , \19277 );
xor \U$19756 ( \20099 , \20097 , \20098 );
and \U$19757 ( \20100 , \20095 , \20099 );
and \U$19758 ( \20101 , \20082 , \20094 );
or \U$19759 ( \20102 , \20100 , \20101 );
and \U$19760 ( \20103 , \19715 , \20102 );
and \U$19761 ( \20104 , \19712 , \19714 );
nor \U$19762 ( \20105 , \20103 , \20104 );
not \U$19763 ( \20106 , \20105 );
xor \U$19764 ( \20107 , \19174 , \19176 );
xor \U$19765 ( \20108 , \20107 , \19195 );
xor \U$19766 ( \20109 , \19690 , \19695 );
xor \U$19767 ( \20110 , \20108 , \20109 );
nand \U$19768 ( \20111 , \20106 , \20110 );
or \U$19769 ( \20112 , \19710 , \20111 );
xnor \U$19770 ( \20113 , \20111 , \19710 );
xor \U$19771 ( \20114 , \19873 , \19898 );
xor \U$19772 ( \20115 , \20114 , \19924 );
not \U$19773 ( \20116 , \20115 );
not \U$19774 ( \20117 , \1301 );
and \U$19775 ( \20118 , \1293 , RI9870600_89);
and \U$19776 ( \20119 , RI98708d0_95, \1291 );
nor \U$19777 ( \20120 , \20118 , \20119 );
not \U$19778 ( \20121 , \20120 );
or \U$19779 ( \20122 , \20117 , \20121 );
or \U$19780 ( \20123 , \20120 , \1301 );
nand \U$19781 ( \20124 , \20122 , \20123 );
and \U$19782 ( \20125 , \1329 , RI98707e0_93);
and \U$19783 ( \20126 , RI986fac0_65, \1327 );
nor \U$19784 ( \20127 , \20125 , \20126 );
and \U$19785 ( \20128 , \20127 , \1336 );
not \U$19786 ( \20129 , \20127 );
and \U$19787 ( \20130 , \20129 , \1337 );
nor \U$19788 ( \20131 , \20128 , \20130 );
xor \U$19789 ( \20132 , \20124 , \20131 );
and \U$19790 ( \20133 , \776 , RI9870240_81);
and \U$19791 ( \20134 , RI98706f0_91, \774 );
nor \U$19792 ( \20135 , \20133 , \20134 );
and \U$19793 ( \20136 , \20135 , \474 );
not \U$19794 ( \20137 , \20135 );
and \U$19795 ( \20138 , \20137 , \451 );
nor \U$19796 ( \20139 , \20136 , \20138 );
and \U$19797 ( \20140 , \20132 , \20139 );
and \U$19798 ( \20141 , \20124 , \20131 );
nor \U$19799 ( \20142 , \20140 , \20141 );
and \U$19800 ( \20143 , \2464 , RI9870150_79);
and \U$19801 ( \20144 , RI9870f60_109, \2462 );
nor \U$19802 ( \20145 , \20143 , \20144 );
and \U$19803 ( \20146 , \20145 , \2263 );
not \U$19804 ( \20147 , \20145 );
and \U$19805 ( \20148 , \20147 , \2468 );
nor \U$19806 ( \20149 , \20146 , \20148 );
and \U$19807 ( \20150 , \3254 , RI9870ab0_99);
and \U$19808 ( \20151 , RI9870d80_105, \3252 );
nor \U$19809 ( \20152 , \20150 , \20151 );
not \U$19810 ( \20153 , \20152 );
not \U$19811 ( \20154 , \2935 );
and \U$19812 ( \20155 , \20153 , \20154 );
and \U$19813 ( \20156 , \20152 , \2935 );
nor \U$19814 ( \20157 , \20155 , \20156 );
xor \U$19815 ( \20158 , \20149 , \20157 );
and \U$19816 ( \20159 , \3683 , RI98709c0_97);
and \U$19817 ( \20160 , RI9870e70_107, \3681 );
nor \U$19818 ( \20161 , \20159 , \20160 );
not \U$19819 ( \20162 , \20161 );
not \U$19820 ( \20163 , \3412 );
and \U$19821 ( \20164 , \20162 , \20163 );
and \U$19822 ( \20165 , \20161 , \3412 );
nor \U$19823 ( \20166 , \20164 , \20165 );
and \U$19824 ( \20167 , \20158 , \20166 );
and \U$19825 ( \20168 , \20149 , \20157 );
or \U$19826 ( \20169 , \20167 , \20168 );
xor \U$19827 ( \20170 , \20142 , \20169 );
and \U$19828 ( \20171 , \1311 , RI986fbb0_67);
and \U$19829 ( \20172 , RI986fd90_71, \1309 );
nor \U$19830 ( \20173 , \20171 , \20172 );
and \U$19831 ( \20174 , \20173 , \1318 );
not \U$19832 ( \20175 , \20173 );
and \U$19833 ( \20176 , \20175 , \1458 );
nor \U$19834 ( \20177 , \20174 , \20176 );
and \U$19835 ( \20178 , \2042 , RI986fca0_69);
and \U$19836 ( \20179 , RI986ff70_75, \2040 );
nor \U$19837 ( \20180 , \20178 , \20179 );
not \U$19838 ( \20181 , \20180 );
not \U$19839 ( \20182 , \2034 );
and \U$19840 ( \20183 , \20181 , \20182 );
and \U$19841 ( \20184 , \20180 , \2034 );
nor \U$19842 ( \20185 , \20183 , \20184 );
xor \U$19843 ( \20186 , \20177 , \20185 );
and \U$19844 ( \20187 , \2274 , RI986fe80_73);
and \U$19845 ( \20188 , RI9870060_77, \2272 );
nor \U$19846 ( \20189 , \20187 , \20188 );
and \U$19847 ( \20190 , \20189 , \2031 );
not \U$19848 ( \20191 , \20189 );
and \U$19849 ( \20192 , \20191 , \2030 );
nor \U$19850 ( \20193 , \20190 , \20192 );
and \U$19851 ( \20194 , \20186 , \20193 );
and \U$19852 ( \20195 , \20177 , \20185 );
or \U$19853 ( \20196 , \20194 , \20195 );
xor \U$19854 ( \20197 , \20170 , \20196 );
and \U$19855 ( \20198 , \7079 , RI98715f0_123);
and \U$19856 ( \20199 , RI986ead0_31, \7077 );
nor \U$19857 ( \20200 , \20198 , \20199 );
and \U$19858 ( \20201 , \20200 , \6710 );
not \U$19859 ( \20202 , \20200 );
and \U$19860 ( \20203 , \20202 , \6709 );
nor \U$19861 ( \20204 , \20201 , \20203 );
and \U$19862 ( \20205 , \5881 , RI9871410_119);
and \U$19863 ( \20206 , RI98716e0_125, \5879 );
nor \U$19864 ( \20207 , \20205 , \20206 );
and \U$19865 ( \20208 , \20207 , \5594 );
not \U$19866 ( \20209 , \20207 );
and \U$19867 ( \20210 , \20209 , \5885 );
nor \U$19868 ( \20211 , \20208 , \20210 );
xor \U$19869 ( \20212 , \20204 , \20211 );
and \U$19870 ( \20213 , \6453 , RI98717d0_127);
and \U$19871 ( \20214 , RI9871500_121, \6451 );
nor \U$19872 ( \20215 , \20213 , \20214 );
and \U$19873 ( \20216 , \20215 , \6190 );
not \U$19874 ( \20217 , \20215 );
and \U$19875 ( \20218 , \20217 , \6705 );
nor \U$19876 ( \20219 , \20216 , \20218 );
and \U$19877 ( \20220 , \20212 , \20219 );
and \U$19878 ( \20221 , \20204 , \20211 );
or \U$19879 ( \20222 , \20220 , \20221 );
not \U$19880 ( \20223 , \20222 );
and \U$19881 ( \20224 , \4203 , RI9870ba0_101);
and \U$19882 ( \20225 , RI9871050_111, \4201 );
nor \U$19883 ( \20226 , \20224 , \20225 );
and \U$19884 ( \20227 , \20226 , \3922 );
not \U$19885 ( \20228 , \20226 );
and \U$19886 ( \20229 , \20228 , \4207 );
nor \U$19887 ( \20230 , \20227 , \20229 );
and \U$19888 ( \20231 , \4710 , RI9870c90_103);
and \U$19889 ( \20232 , RI9871230_115, \4708 );
nor \U$19890 ( \20233 , \20231 , \20232 );
not \U$19891 ( \20234 , \20233 );
not \U$19892 ( \20235 , \4519 );
and \U$19893 ( \20236 , \20234 , \20235 );
and \U$19894 ( \20237 , \20233 , \4521 );
nor \U$19895 ( \20238 , \20236 , \20237 );
xor \U$19896 ( \20239 , \20230 , \20238 );
and \U$19897 ( \20240 , \5318 , RI9871140_113);
and \U$19898 ( \20241 , RI9871320_117, \5316 );
nor \U$19899 ( \20242 , \20240 , \20241 );
and \U$19900 ( \20243 , \20242 , \5322 );
not \U$19901 ( \20244 , \20242 );
and \U$19902 ( \20245 , \20244 , \5052 );
nor \U$19903 ( \20246 , \20243 , \20245 );
and \U$19904 ( \20247 , \20239 , \20246 );
and \U$19905 ( \20248 , \20230 , \20238 );
or \U$19906 ( \20249 , \20247 , \20248 );
not \U$19907 ( \20250 , \20249 );
or \U$19908 ( \20251 , \20223 , \20250 );
or \U$19909 ( \20252 , \20249 , \20222 );
nand \U$19910 ( \20253 , \20251 , \20252 );
not \U$19911 ( \20254 , \20253 );
and \U$19912 ( \20255 , \8486 , RI986e800_25);
and \U$19913 ( \20256 , RI986ee90_39, \8484 );
nor \U$19914 ( \20257 , \20255 , \20256 );
and \U$19915 ( \20258 , \20257 , \8050 );
not \U$19916 ( \20259 , \20257 );
and \U$19917 ( \20260 , \20259 , \8051 );
nor \U$19918 ( \20261 , \20258 , \20260 );
and \U$19919 ( \20262 , \9237 , RI986eda0_37);
and \U$19920 ( \20263 , RI986ebc0_33, \9235 );
nor \U$19921 ( \20264 , \20262 , \20263 );
and \U$19922 ( \20265 , \20264 , \9241 );
not \U$19923 ( \20266 , \20264 );
and \U$19924 ( \20267 , \20266 , \8836 );
nor \U$19925 ( \20268 , \20265 , \20267 );
xor \U$19926 ( \20269 , \20261 , \20268 );
and \U$19927 ( \20270 , \7729 , RI986e9e0_29);
and \U$19928 ( \20271 , RI986e8f0_27, \7727 );
nor \U$19929 ( \20272 , \20270 , \20271 );
and \U$19930 ( \20273 , \20272 , \7480 );
not \U$19931 ( \20274 , \20272 );
and \U$19932 ( \20275 , \20274 , \7733 );
nor \U$19933 ( \20276 , \20273 , \20275 );
and \U$19934 ( \20277 , \20269 , \20276 );
and \U$19935 ( \20278 , \20261 , \20268 );
nor \U$19936 ( \20279 , \20277 , \20278 );
not \U$19937 ( \20280 , \20279 );
and \U$19938 ( \20281 , \20254 , \20280 );
and \U$19939 ( \20282 , \20253 , \20279 );
nor \U$19940 ( \20283 , \20281 , \20282 );
xor \U$19941 ( \20284 , \20197 , \20283 );
and \U$19942 ( \20285 , \465 , RI9870420_85);
and \U$19943 ( \20286 , RI9870510_87, \463 );
nor \U$19944 ( \20287 , \20285 , \20286 );
not \U$19945 ( \20288 , \20287 );
not \U$19946 ( \20289 , \456 );
and \U$19947 ( \20290 , \20288 , \20289 );
and \U$19948 ( \20291 , \20287 , \454 );
nor \U$19949 ( \20292 , \20290 , \20291 );
not \U$19950 ( \20293 , \20292 );
xor \U$19951 ( \20294 , \19827 , \19834 );
xor \U$19952 ( \20295 , \20294 , \19842 );
not \U$19953 ( \20296 , \20295 );
or \U$19954 ( \20297 , \20293 , \20296 );
or \U$19955 ( \20298 , \20295 , \20292 );
nand \U$19956 ( \20299 , \20297 , \20298 );
not \U$19957 ( \20300 , \20299 );
xor \U$19958 ( \20301 , \19771 , \19778 );
xor \U$19959 ( \20302 , \20301 , \19786 );
not \U$19960 ( \20303 , \20302 );
and \U$19961 ( \20304 , \20300 , \20303 );
and \U$19962 ( \20305 , \20299 , \20302 );
nor \U$19963 ( \20306 , \20304 , \20305 );
and \U$19964 ( \20307 , \20284 , \20306 );
and \U$19965 ( \20308 , \20197 , \20283 );
nor \U$19966 ( \20309 , \20307 , \20308 );
not \U$19967 ( \20310 , \20309 );
or \U$19968 ( \20311 , \20116 , \20310 );
or \U$19969 ( \20312 , \20309 , \20115 );
nand \U$19970 ( \20313 , \20311 , \20312 );
not \U$19971 ( \20314 , \20313 );
xor \U$19972 ( \20315 , \19955 , \19982 );
xor \U$19973 ( \20316 , \20315 , \20008 );
not \U$19974 ( \20317 , \19845 );
not \U$19975 ( \20318 , \19789 );
or \U$19976 ( \20319 , \20317 , \20318 );
or \U$19977 ( \20320 , \19789 , \19845 );
nand \U$19978 ( \20321 , \20319 , \20320 );
not \U$19979 ( \20322 , \20321 );
not \U$19980 ( \20323 , \19815 );
and \U$19981 ( \20324 , \20322 , \20323 );
and \U$19982 ( \20325 , \20321 , \19815 );
nor \U$19983 ( \20326 , \20324 , \20325 );
xor \U$19984 ( \20327 , \20316 , \20326 );
not \U$19985 ( \20328 , \19741 );
not \U$19986 ( \20329 , \19747 );
or \U$19987 ( \20330 , \20328 , \20329 );
or \U$19988 ( \20331 , \19747 , \19741 );
nand \U$19989 ( \20332 , \20330 , \20331 );
not \U$19990 ( \20333 , \20332 );
not \U$19991 ( \20334 , \19731 );
and \U$19992 ( \20335 , \20333 , \20334 );
and \U$19993 ( \20336 , \20332 , \19731 );
nor \U$19994 ( \20337 , \20335 , \20336 );
xor \U$19995 ( \20338 , \20327 , \20337 );
not \U$19996 ( \20339 , \20338 );
and \U$19997 ( \20340 , \20314 , \20339 );
and \U$19998 ( \20341 , \20313 , \20338 );
nor \U$19999 ( \20342 , \20340 , \20341 );
and \U$20000 ( \20343 , \2274 , RI986ff70_75);
and \U$20001 ( \20344 , RI986fe80_73, \2272 );
nor \U$20002 ( \20345 , \20343 , \20344 );
and \U$20003 ( \20346 , \20345 , \2030 );
not \U$20004 ( \20347 , \20345 );
and \U$20005 ( \20348 , \20347 , \2031 );
nor \U$20006 ( \20349 , \20346 , \20348 );
and \U$20007 ( \20350 , \2464 , RI9870060_77);
and \U$20008 ( \20351 , RI9870150_79, \2462 );
nor \U$20009 ( \20352 , \20350 , \20351 );
and \U$20010 ( \20353 , \20352 , \2468 );
not \U$20011 ( \20354 , \20352 );
and \U$20012 ( \20355 , \20354 , \2263 );
nor \U$20013 ( \20356 , \20353 , \20355 );
xor \U$20014 ( \20357 , \20349 , \20356 );
not \U$20015 ( \20358 , \2935 );
and \U$20016 ( \20359 , \3254 , RI9870f60_109);
and \U$20017 ( \20360 , RI9870ab0_99, \3252 );
nor \U$20018 ( \20361 , \20359 , \20360 );
not \U$20019 ( \20362 , \20361 );
or \U$20020 ( \20363 , \20358 , \20362 );
or \U$20021 ( \20364 , \20361 , \2935 );
nand \U$20022 ( \20365 , \20363 , \20364 );
and \U$20023 ( \20366 , \20357 , \20365 );
and \U$20024 ( \20367 , \20349 , \20356 );
or \U$20025 ( \20368 , \20366 , \20367 );
and \U$20026 ( \20369 , \438 , RI9870420_85);
and \U$20027 ( \20370 , RI9870510_87, \436 );
nor \U$20028 ( \20371 , \20369 , \20370 );
and \U$20029 ( \20372 , \20371 , \444 );
not \U$20030 ( \20373 , \20371 );
and \U$20031 ( \20374 , \20373 , \443 );
nor \U$20032 ( \20375 , \20372 , \20374 );
and \U$20033 ( \20376 , \776 , RI9870330_83);
and \U$20034 ( \20377 , RI9870240_81, \774 );
nor \U$20035 ( \20378 , \20376 , \20377 );
and \U$20036 ( \20379 , \20378 , \474 );
not \U$20037 ( \20380 , \20378 );
and \U$20038 ( \20381 , \20380 , \451 );
nor \U$20039 ( \20382 , \20379 , \20381 );
xor \U$20040 ( \20383 , \20375 , \20382 );
not \U$20041 ( \20384 , \1301 );
and \U$20042 ( \20385 , \1293 , RI98706f0_91);
and \U$20043 ( \20386 , RI9870600_89, \1291 );
nor \U$20044 ( \20387 , \20385 , \20386 );
not \U$20045 ( \20388 , \20387 );
or \U$20046 ( \20389 , \20384 , \20388 );
or \U$20047 ( \20390 , \20387 , \1301 );
nand \U$20048 ( \20391 , \20389 , \20390 );
and \U$20049 ( \20392 , \20383 , \20391 );
and \U$20050 ( \20393 , \20375 , \20382 );
or \U$20051 ( \20394 , \20392 , \20393 );
xor \U$20052 ( \20395 , \20368 , \20394 );
and \U$20053 ( \20396 , \1329 , RI98708d0_95);
and \U$20054 ( \20397 , RI98707e0_93, \1327 );
nor \U$20055 ( \20398 , \20396 , \20397 );
and \U$20056 ( \20399 , \20398 , \1336 );
not \U$20057 ( \20400 , \20398 );
and \U$20058 ( \20401 , \20400 , \1337 );
nor \U$20059 ( \20402 , \20399 , \20401 );
and \U$20060 ( \20403 , \1311 , RI986fac0_65);
and \U$20061 ( \20404 , RI986fbb0_67, \1309 );
nor \U$20062 ( \20405 , \20403 , \20404 );
and \U$20063 ( \20406 , \20405 , \1458 );
not \U$20064 ( \20407 , \20405 );
and \U$20065 ( \20408 , \20407 , \1318 );
nor \U$20066 ( \20409 , \20406 , \20408 );
xor \U$20067 ( \20410 , \20402 , \20409 );
not \U$20068 ( \20411 , \2034 );
and \U$20069 ( \20412 , \2042 , RI986fd90_71);
and \U$20070 ( \20413 , RI986fca0_69, \2040 );
nor \U$20071 ( \20414 , \20412 , \20413 );
not \U$20072 ( \20415 , \20414 );
or \U$20073 ( \20416 , \20411 , \20415 );
or \U$20074 ( \20417 , \20414 , \1462 );
nand \U$20075 ( \20418 , \20416 , \20417 );
and \U$20076 ( \20419 , \20410 , \20418 );
and \U$20077 ( \20420 , \20402 , \20409 );
or \U$20078 ( \20421 , \20419 , \20420 );
and \U$20079 ( \20422 , \20395 , \20421 );
and \U$20080 ( \20423 , \20368 , \20394 );
nor \U$20081 ( \20424 , \20422 , \20423 );
and \U$20082 ( \20425 , \11696 , RI986f250_47);
and \U$20083 ( \20426 , RI986f160_45, \11694 );
nor \U$20084 ( \20427 , \20425 , \20426 );
and \U$20085 ( \20428 , \20427 , \10965 );
not \U$20086 ( \20429 , \20427 );
and \U$20087 ( \20430 , \20429 , \11702 );
nor \U$20088 ( \20431 , \20428 , \20430 );
and \U$20089 ( \20432 , \12293 , RI986e530_19);
and \U$20090 ( \20433 , RI986e440_17, \12291 );
nor \U$20091 ( \20434 , \20432 , \20433 );
and \U$20092 ( \20435 , \20434 , \11687 );
not \U$20093 ( \20436 , \20434 );
and \U$20094 ( \20437 , \20436 , \11686 );
nor \U$20095 ( \20438 , \20435 , \20437 );
xor \U$20096 ( \20439 , \20431 , \20438 );
and \U$20097 ( \20440 , \13045 , RI986e710_23);
and \U$20098 ( \20441 , RI986e620_21, \13043 );
nor \U$20099 ( \20442 , \20440 , \20441 );
and \U$20100 ( \20443 , \20442 , \13047 );
not \U$20101 ( \20444 , \20442 );
and \U$20102 ( \20445 , \20444 , \12619 );
nor \U$20103 ( \20446 , \20443 , \20445 );
and \U$20104 ( \20447 , \20439 , \20446 );
and \U$20105 ( \20448 , \20431 , \20438 );
or \U$20106 ( \20449 , \20447 , \20448 );
and \U$20107 ( \20450 , \9237 , RI986ee90_39);
and \U$20108 ( \20451 , RI986eda0_37, \9235 );
nor \U$20109 ( \20452 , \20450 , \20451 );
and \U$20110 ( \20453 , \20452 , \9241 );
not \U$20111 ( \20454 , \20452 );
and \U$20112 ( \20455 , \20454 , \8836 );
nor \U$20113 ( \20456 , \20453 , \20455 );
and \U$20114 ( \20457 , \9505 , RI986ebc0_33);
and \U$20115 ( \20458 , RI986ecb0_35, \9503 );
nor \U$20116 ( \20459 , \20457 , \20458 );
and \U$20117 ( \20460 , \20459 , \9510 );
not \U$20118 ( \20461 , \20459 );
and \U$20119 ( \20462 , \20461 , \9513 );
nor \U$20120 ( \20463 , \20460 , \20462 );
xor \U$20121 ( \20464 , \20456 , \20463 );
and \U$20122 ( \20465 , \10424 , RI986f070_43);
and \U$20123 ( \20466 , RI986ef80_41, \10422 );
nor \U$20124 ( \20467 , \20465 , \20466 );
and \U$20125 ( \20468 , \20467 , \9840 );
not \U$20126 ( \20469 , \20467 );
and \U$20127 ( \20470 , \20469 , \10428 );
nor \U$20128 ( \20471 , \20468 , \20470 );
and \U$20129 ( \20472 , \20464 , \20471 );
and \U$20130 ( \20473 , \20456 , \20463 );
or \U$20131 ( \20474 , \20472 , \20473 );
xor \U$20132 ( \20475 , \20449 , \20474 );
and \U$20133 ( \20476 , \13882 , RI986f7f0_59);
and \U$20134 ( \20477 , RI986f700_57, \13880 );
nor \U$20135 ( \20478 , \20476 , \20477 );
and \U$20136 ( \20479 , \20478 , \13358 );
not \U$20137 ( \20480 , \20478 );
and \U$20138 ( \20481 , \20480 , \13359 );
nor \U$20139 ( \20482 , \20479 , \20481 );
not \U$20140 ( \20483 , RI9873558_190);
and \U$20141 ( \20484 , \15780 , RI986f430_51);
and \U$20142 ( \20485 , RI9873648_192, RI986f340_49);
nor \U$20143 ( \20486 , \20484 , \20485 );
not \U$20144 ( \20487 , \20486 );
or \U$20145 ( \20488 , \20483 , \20487 );
or \U$20146 ( \20489 , \20486 , RI9873558_190);
nand \U$20147 ( \20490 , \20488 , \20489 );
xor \U$20148 ( \20491 , \20482 , \20490 );
and \U$20149 ( \20492 , \14937 , RI986f9d0_63);
and \U$20150 ( \20493 , RI986f8e0_61, \14935 );
nor \U$20151 ( \20494 , \20492 , \20493 );
and \U$20152 ( \20495 , \20494 , \14539 );
not \U$20153 ( \20496 , \20494 );
and \U$20154 ( \20497 , \20496 , \14538 );
nor \U$20155 ( \20498 , \20495 , \20497 );
and \U$20156 ( \20499 , \20491 , \20498 );
and \U$20157 ( \20500 , \20482 , \20490 );
or \U$20158 ( \20501 , \20499 , \20500 );
and \U$20159 ( \20502 , \20475 , \20501 );
and \U$20160 ( \20503 , \20449 , \20474 );
nor \U$20161 ( \20504 , \20502 , \20503 );
xor \U$20162 ( \20505 , \20424 , \20504 );
and \U$20163 ( \20506 , \5318 , RI9871230_115);
and \U$20164 ( \20507 , RI9871140_113, \5316 );
nor \U$20165 ( \20508 , \20506 , \20507 );
and \U$20166 ( \20509 , \20508 , \5052 );
not \U$20167 ( \20510 , \20508 );
and \U$20168 ( \20511 , \20510 , \5322 );
nor \U$20169 ( \20512 , \20509 , \20511 );
and \U$20170 ( \20513 , \5881 , RI9871320_117);
and \U$20171 ( \20514 , RI9871410_119, \5879 );
nor \U$20172 ( \20515 , \20513 , \20514 );
and \U$20173 ( \20516 , \20515 , \5594 );
not \U$20174 ( \20517 , \20515 );
and \U$20175 ( \20518 , \20517 , \5885 );
nor \U$20176 ( \20519 , \20516 , \20518 );
xor \U$20177 ( \20520 , \20512 , \20519 );
and \U$20178 ( \20521 , \6453 , RI98716e0_125);
and \U$20179 ( \20522 , RI98717d0_127, \6451 );
nor \U$20180 ( \20523 , \20521 , \20522 );
and \U$20181 ( \20524 , \20523 , \6190 );
not \U$20182 ( \20525 , \20523 );
and \U$20183 ( \20526 , \20525 , \6180 );
nor \U$20184 ( \20527 , \20524 , \20526 );
and \U$20185 ( \20528 , \20520 , \20527 );
and \U$20186 ( \20529 , \20512 , \20519 );
or \U$20187 ( \20530 , \20528 , \20529 );
not \U$20188 ( \20531 , \3412 );
and \U$20189 ( \20532 , \3683 , RI9870d80_105);
and \U$20190 ( \20533 , RI98709c0_97, \3681 );
nor \U$20191 ( \20534 , \20532 , \20533 );
not \U$20192 ( \20535 , \20534 );
or \U$20193 ( \20536 , \20531 , \20535 );
or \U$20194 ( \20537 , \20534 , \3918 );
nand \U$20195 ( \20538 , \20536 , \20537 );
and \U$20196 ( \20539 , \4203 , RI9870e70_107);
and \U$20197 ( \20540 , RI9870ba0_101, \4201 );
nor \U$20198 ( \20541 , \20539 , \20540 );
and \U$20199 ( \20542 , \20541 , \4207 );
not \U$20200 ( \20543 , \20541 );
and \U$20201 ( \20544 , \20543 , \3922 );
nor \U$20202 ( \20545 , \20542 , \20544 );
xor \U$20203 ( \20546 , \20538 , \20545 );
not \U$20204 ( \20547 , \4521 );
and \U$20205 ( \20548 , \4710 , RI9871050_111);
and \U$20206 ( \20549 , RI9870c90_103, \4708 );
nor \U$20207 ( \20550 , \20548 , \20549 );
not \U$20208 ( \20551 , \20550 );
or \U$20209 ( \20552 , \20547 , \20551 );
or \U$20210 ( \20553 , \20550 , \4519 );
nand \U$20211 ( \20554 , \20552 , \20553 );
and \U$20212 ( \20555 , \20546 , \20554 );
and \U$20213 ( \20556 , \20538 , \20545 );
or \U$20214 ( \20557 , \20555 , \20556 );
xor \U$20215 ( \20558 , \20530 , \20557 );
and \U$20216 ( \20559 , \7079 , RI9871500_121);
and \U$20217 ( \20560 , RI98715f0_123, \7077 );
nor \U$20218 ( \20561 , \20559 , \20560 );
and \U$20219 ( \20562 , \20561 , \6710 );
not \U$20220 ( \20563 , \20561 );
and \U$20221 ( \20564 , \20563 , \6709 );
nor \U$20222 ( \20565 , \20562 , \20564 );
and \U$20223 ( \20566 , \7729 , RI986ead0_31);
and \U$20224 ( \20567 , RI986e9e0_29, \7727 );
nor \U$20225 ( \20568 , \20566 , \20567 );
and \U$20226 ( \20569 , \20568 , \7480 );
not \U$20227 ( \20570 , \20568 );
and \U$20228 ( \20571 , \20570 , \7733 );
nor \U$20229 ( \20572 , \20569 , \20571 );
xor \U$20230 ( \20573 , \20565 , \20572 );
and \U$20231 ( \20574 , \8486 , RI986e8f0_27);
and \U$20232 ( \20575 , RI986e800_25, \8484 );
nor \U$20233 ( \20576 , \20574 , \20575 );
and \U$20234 ( \20577 , \20576 , \8050 );
not \U$20235 ( \20578 , \20576 );
and \U$20236 ( \20579 , \20578 , \8051 );
nor \U$20237 ( \20580 , \20577 , \20579 );
and \U$20238 ( \20581 , \20573 , \20580 );
and \U$20239 ( \20582 , \20565 , \20572 );
or \U$20240 ( \20583 , \20581 , \20582 );
and \U$20241 ( \20584 , \20558 , \20583 );
and \U$20242 ( \20585 , \20530 , \20557 );
nor \U$20243 ( \20586 , \20584 , \20585 );
and \U$20244 ( \20587 , \20505 , \20586 );
and \U$20245 ( \20588 , \20424 , \20504 );
or \U$20246 ( \20589 , \20587 , \20588 );
xor \U$20247 ( \20590 , \20177 , \20185 );
xor \U$20248 ( \20591 , \20590 , \20193 );
not \U$20249 ( \20592 , \20591 );
xor \U$20250 ( \20593 , \20230 , \20238 );
xor \U$20251 ( \20594 , \20593 , \20246 );
not \U$20252 ( \20595 , \20594 );
and \U$20253 ( \20596 , \20592 , \20595 );
and \U$20254 ( \20597 , \20594 , \20591 );
xor \U$20255 ( \20598 , \20149 , \20157 );
xor \U$20256 ( \20599 , \20598 , \20166 );
nor \U$20257 ( \20600 , \20597 , \20599 );
nor \U$20258 ( \20601 , \20596 , \20600 );
nand \U$20259 ( \20602 , RI9870420_85, \463 );
not \U$20260 ( \20603 , \20602 );
not \U$20261 ( \20604 , \454 );
or \U$20262 ( \20605 , \20603 , \20604 );
or \U$20263 ( \20606 , \454 , \20602 );
nand \U$20264 ( \20607 , \20605 , \20606 );
and \U$20265 ( \20608 , \438 , RI9870510_87);
and \U$20266 ( \20609 , RI9870330_83, \436 );
nor \U$20267 ( \20610 , \20608 , \20609 );
and \U$20268 ( \20611 , \20610 , \444 );
not \U$20269 ( \20612 , \20610 );
and \U$20270 ( \20613 , \20612 , \443 );
nor \U$20271 ( \20614 , \20611 , \20613 );
xor \U$20272 ( \20615 , \20607 , \20614 );
xor \U$20273 ( \20616 , \20124 , \20131 );
xor \U$20274 ( \20617 , \20616 , \20139 );
and \U$20275 ( \20618 , \20615 , \20617 );
and \U$20276 ( \20619 , \20607 , \20614 );
nor \U$20277 ( \20620 , \20618 , \20619 );
xor \U$20278 ( \20621 , \20601 , \20620 );
xor \U$20279 ( \20622 , \20204 , \20211 );
xor \U$20280 ( \20623 , \20622 , \20219 );
and \U$20281 ( \20624 , \11696 , RI986f160_45);
and \U$20282 ( \20625 , RI986e530_19, \11694 );
nor \U$20283 ( \20626 , \20624 , \20625 );
and \U$20284 ( \20627 , \20626 , \10965 );
not \U$20285 ( \20628 , \20626 );
and \U$20286 ( \20629 , \20628 , \11702 );
nor \U$20287 ( \20630 , \20627 , \20629 );
and \U$20288 ( \20631 , \9505 , RI986ecb0_35);
and \U$20289 ( \20632 , RI986f070_43, \9503 );
nor \U$20290 ( \20633 , \20631 , \20632 );
and \U$20291 ( \20634 , \20633 , \9510 );
not \U$20292 ( \20635 , \20633 );
and \U$20293 ( \20636 , \20635 , \9513 );
nor \U$20294 ( \20637 , \20634 , \20636 );
xor \U$20295 ( \20638 , \20630 , \20637 );
and \U$20296 ( \20639 , \10424 , RI986ef80_41);
and \U$20297 ( \20640 , RI986f250_47, \10422 );
nor \U$20298 ( \20641 , \20639 , \20640 );
and \U$20299 ( \20642 , \20641 , \9840 );
not \U$20300 ( \20643 , \20641 );
and \U$20301 ( \20644 , \20643 , \10428 );
nor \U$20302 ( \20645 , \20642 , \20644 );
xor \U$20303 ( \20646 , \20638 , \20645 );
and \U$20304 ( \20647 , \20623 , \20646 );
xor \U$20305 ( \20648 , \20261 , \20268 );
xor \U$20306 ( \20649 , \20648 , \20276 );
xor \U$20307 ( \20650 , \20630 , \20637 );
xor \U$20308 ( \20651 , \20650 , \20645 );
and \U$20309 ( \20652 , \20649 , \20651 );
and \U$20310 ( \20653 , \20623 , \20649 );
or \U$20311 ( \20654 , \20647 , \20652 , \20653 );
not \U$20312 ( \20655 , \20654 );
and \U$20313 ( \20656 , \20621 , \20655 );
and \U$20314 ( \20657 , \20601 , \20620 );
or \U$20315 ( \20658 , \20656 , \20657 );
xor \U$20316 ( \20659 , \20589 , \20658 );
xor \U$20317 ( \20660 , \19936 , \19944 );
xor \U$20318 ( \20661 , \20660 , \19952 );
not \U$20319 ( \20662 , \20661 );
xor \U$20320 ( \20663 , \19990 , \19997 );
xor \U$20321 ( \20664 , \20663 , \20005 );
not \U$20322 ( \20665 , \20664 );
or \U$20323 ( \20666 , \20662 , \20665 );
or \U$20324 ( \20667 , \20661 , \20664 );
nand \U$20325 ( \20668 , \20666 , \20667 );
not \U$20326 ( \20669 , \20668 );
xor \U$20327 ( \20670 , \19797 , \19804 );
xor \U$20328 ( \20671 , \20670 , \19812 );
not \U$20329 ( \20672 , \20671 );
and \U$20330 ( \20673 , \20669 , \20672 );
and \U$20331 ( \20674 , \20668 , \20671 );
nor \U$20332 ( \20675 , \20673 , \20674 );
xor \U$20333 ( \20676 , \19854 , \19862 );
xor \U$20334 ( \20677 , \20676 , \19870 );
xor \U$20335 ( \20678 , \20675 , \20677 );
xor \U$20336 ( \20679 , \19880 , \19887 );
xor \U$20337 ( \20680 , \20679 , \19895 );
not \U$20338 ( \20681 , \20680 );
not \U$20339 ( \20682 , \19962 );
xor \U$20340 ( \20683 , \19980 , \19970 );
not \U$20341 ( \20684 , \20683 );
or \U$20342 ( \20685 , \20682 , \20684 );
or \U$20343 ( \20686 , \20683 , \19962 );
nand \U$20344 ( \20687 , \20685 , \20686 );
not \U$20345 ( \20688 , \20687 );
or \U$20346 ( \20689 , \20681 , \20688 );
or \U$20347 ( \20690 , \20680 , \20687 );
nand \U$20348 ( \20691 , \20689 , \20690 );
not \U$20349 ( \20692 , \20691 );
xor \U$20350 ( \20693 , \19906 , \19913 );
xor \U$20351 ( \20694 , \20693 , \19921 );
not \U$20352 ( \20695 , \20694 );
and \U$20353 ( \20696 , \20692 , \20695 );
and \U$20354 ( \20697 , \20691 , \20694 );
nor \U$20355 ( \20698 , \20696 , \20697 );
and \U$20356 ( \20699 , \20678 , \20698 );
and \U$20357 ( \20700 , \20675 , \20677 );
or \U$20358 ( \20701 , \20699 , \20700 );
xor \U$20359 ( \20702 , \20659 , \20701 );
or \U$20360 ( \20703 , \20342 , \20702 );
not \U$20361 ( \20704 , \20702 );
not \U$20362 ( \20705 , \20342 );
or \U$20363 ( \20706 , \20704 , \20705 );
or \U$20364 ( \20707 , \20671 , \20661 );
not \U$20365 ( \20708 , \20661 );
not \U$20366 ( \20709 , \20671 );
or \U$20367 ( \20710 , \20708 , \20709 );
nand \U$20368 ( \20711 , \20710 , \20664 );
nand \U$20369 ( \20712 , \20707 , \20711 );
or \U$20370 ( \20713 , \20302 , \20292 );
not \U$20371 ( \20714 , \20292 );
not \U$20372 ( \20715 , \20302 );
or \U$20373 ( \20716 , \20714 , \20715 );
nand \U$20374 ( \20717 , \20716 , \20295 );
nand \U$20375 ( \20718 , \20713 , \20717 );
xor \U$20376 ( \20719 , \20712 , \20718 );
or \U$20377 ( \20720 , \20680 , \20694 );
not \U$20378 ( \20721 , \20694 );
not \U$20379 ( \20722 , \20680 );
or \U$20380 ( \20723 , \20721 , \20722 );
nand \U$20381 ( \20724 , \20723 , \20687 );
nand \U$20382 ( \20725 , \20720 , \20724 );
xor \U$20383 ( \20726 , \20719 , \20725 );
xor \U$20384 ( \20727 , \20142 , \20169 );
and \U$20385 ( \20728 , \20727 , \20196 );
and \U$20386 ( \20729 , \20142 , \20169 );
nor \U$20387 ( \20730 , \20728 , \20729 );
xor \U$20388 ( \20731 , \20630 , \20637 );
and \U$20389 ( \20732 , \20731 , \20645 );
and \U$20390 ( \20733 , \20630 , \20637 );
or \U$20391 ( \20734 , \20732 , \20733 );
not \U$20392 ( \20735 , RI9873558_190);
and \U$20393 ( \20736 , \15780 , RI986f340_49);
and \U$20394 ( \20737 , RI9873648_192, RI986f520_53);
nor \U$20395 ( \20738 , \20736 , \20737 );
not \U$20396 ( \20739 , \20738 );
or \U$20397 ( \20740 , \20735 , \20739 );
or \U$20398 ( \20741 , \20738 , RI9873558_190);
nand \U$20399 ( \20742 , \20740 , \20741 );
xor \U$20400 ( \20743 , \20742 , \456 );
and \U$20401 ( \20744 , \14937 , RI986f8e0_61);
and \U$20402 ( \20745 , RI986f430_51, \14935 );
nor \U$20403 ( \20746 , \20744 , \20745 );
and \U$20404 ( \20747 , \20746 , \14539 );
not \U$20405 ( \20748 , \20746 );
and \U$20406 ( \20749 , \20748 , \14538 );
nor \U$20407 ( \20750 , \20747 , \20749 );
and \U$20408 ( \20751 , \20743 , \20750 );
and \U$20409 ( \20752 , \20742 , \456 );
or \U$20410 ( \20753 , \20751 , \20752 );
xor \U$20411 ( \20754 , \20734 , \20753 );
and \U$20412 ( \20755 , \12293 , RI986e440_17);
and \U$20413 ( \20756 , RI986e710_23, \12291 );
nor \U$20414 ( \20757 , \20755 , \20756 );
and \U$20415 ( \20758 , \20757 , \11687 );
not \U$20416 ( \20759 , \20757 );
and \U$20417 ( \20760 , \20759 , \11686 );
nor \U$20418 ( \20761 , \20758 , \20760 );
and \U$20419 ( \20762 , \13045 , RI986e620_21);
and \U$20420 ( \20763 , RI986f7f0_59, \13043 );
nor \U$20421 ( \20764 , \20762 , \20763 );
and \U$20422 ( \20765 , \20764 , \13047 );
not \U$20423 ( \20766 , \20764 );
and \U$20424 ( \20767 , \20766 , \12619 );
nor \U$20425 ( \20768 , \20765 , \20767 );
xor \U$20426 ( \20769 , \20761 , \20768 );
and \U$20427 ( \20770 , \13882 , RI986f700_57);
and \U$20428 ( \20771 , RI986f9d0_63, \13880 );
nor \U$20429 ( \20772 , \20770 , \20771 );
and \U$20430 ( \20773 , \20772 , \13358 );
not \U$20431 ( \20774 , \20772 );
and \U$20432 ( \20775 , \20774 , \13359 );
nor \U$20433 ( \20776 , \20773 , \20775 );
and \U$20434 ( \20777 , \20769 , \20776 );
and \U$20435 ( \20778 , \20761 , \20768 );
or \U$20436 ( \20779 , \20777 , \20778 );
and \U$20437 ( \20780 , \20754 , \20779 );
and \U$20438 ( \20781 , \20734 , \20753 );
or \U$20439 ( \20782 , \20780 , \20781 );
xor \U$20440 ( \20783 , \20730 , \20782 );
or \U$20441 ( \20784 , \20249 , \20279 );
not \U$20442 ( \20785 , \20249 );
not \U$20443 ( \20786 , \20279 );
or \U$20444 ( \20787 , \20785 , \20786 );
nand \U$20445 ( \20788 , \20787 , \20222 );
nand \U$20446 ( \20789 , \20784 , \20788 );
xor \U$20447 ( \20790 , \20783 , \20789 );
xor \U$20448 ( \20791 , \19752 , \19754 );
xor \U$20449 ( \20792 , \20791 , \19757 );
xor \U$20450 ( \20793 , \19393 , \367 );
xor \U$20451 ( \20794 , \20793 , \19401 );
xor \U$20452 ( \20795 , \19717 , \19723 );
xor \U$20453 ( \20796 , \20795 , \19726 );
xor \U$20454 ( \20797 , \20794 , \20796 );
xor \U$20455 ( \20798 , \20792 , \20797 );
xor \U$20456 ( \20799 , \20790 , \20798 );
xor \U$20457 ( \20800 , \20726 , \20799 );
nand \U$20458 ( \20801 , \20706 , \20800 );
nand \U$20459 ( \20802 , \20703 , \20801 );
xor \U$20460 ( \20803 , \20761 , \20768 );
xor \U$20461 ( \20804 , \20803 , \20776 );
xor \U$20462 ( \20805 , \20742 , \456 );
xor \U$20463 ( \20806 , \20805 , \20750 );
and \U$20464 ( \20807 , \20804 , \20806 );
xor \U$20465 ( \20808 , \20630 , \20637 );
xor \U$20466 ( \20809 , \20808 , \20645 );
xor \U$20467 ( \20810 , \20623 , \20649 );
xor \U$20468 ( \20811 , \20809 , \20810 );
xor \U$20469 ( \20812 , \20742 , \456 );
xor \U$20470 ( \20813 , \20812 , \20750 );
and \U$20471 ( \20814 , \20811 , \20813 );
and \U$20472 ( \20815 , \20804 , \20811 );
or \U$20473 ( \20816 , \20807 , \20814 , \20815 );
and \U$20474 ( \20817 , \7729 , RI98715f0_123);
and \U$20475 ( \20818 , RI986ead0_31, \7727 );
nor \U$20476 ( \20819 , \20817 , \20818 );
and \U$20477 ( \20820 , \20819 , \7480 );
not \U$20478 ( \20821 , \20819 );
and \U$20479 ( \20822 , \20821 , \7733 );
nor \U$20480 ( \20823 , \20820 , \20822 );
and \U$20481 ( \20824 , \8486 , RI986e9e0_29);
and \U$20482 ( \20825 , RI986e8f0_27, \8484 );
nor \U$20483 ( \20826 , \20824 , \20825 );
and \U$20484 ( \20827 , \20826 , \8050 );
not \U$20485 ( \20828 , \20826 );
and \U$20486 ( \20829 , \20828 , \8051 );
nor \U$20487 ( \20830 , \20827 , \20829 );
xor \U$20488 ( \20831 , \20823 , \20830 );
and \U$20489 ( \20832 , \9237 , RI986e800_25);
and \U$20490 ( \20833 , RI986ee90_39, \9235 );
nor \U$20491 ( \20834 , \20832 , \20833 );
and \U$20492 ( \20835 , \20834 , \9241 );
not \U$20493 ( \20836 , \20834 );
and \U$20494 ( \20837 , \20836 , \8836 );
nor \U$20495 ( \20838 , \20835 , \20837 );
and \U$20496 ( \20839 , \20831 , \20838 );
and \U$20497 ( \20840 , \20823 , \20830 );
or \U$20498 ( \20841 , \20839 , \20840 );
not \U$20499 ( \20842 , \4521 );
and \U$20500 ( \20843 , \4710 , RI9870ba0_101);
and \U$20501 ( \20844 , RI9871050_111, \4708 );
nor \U$20502 ( \20845 , \20843 , \20844 );
not \U$20503 ( \20846 , \20845 );
or \U$20504 ( \20847 , \20842 , \20846 );
or \U$20505 ( \20848 , \20845 , \4519 );
nand \U$20506 ( \20849 , \20847 , \20848 );
and \U$20507 ( \20850 , \4203 , RI98709c0_97);
and \U$20508 ( \20851 , RI9870e70_107, \4201 );
nor \U$20509 ( \20852 , \20850 , \20851 );
and \U$20510 ( \20853 , \20852 , \4207 );
not \U$20511 ( \20854 , \20852 );
and \U$20512 ( \20855 , \20854 , \3922 );
nor \U$20513 ( \20856 , \20853 , \20855 );
xor \U$20514 ( \20857 , \20849 , \20856 );
and \U$20515 ( \20858 , \5318 , RI9870c90_103);
and \U$20516 ( \20859 , RI9871230_115, \5316 );
nor \U$20517 ( \20860 , \20858 , \20859 );
and \U$20518 ( \20861 , \20860 , \5052 );
not \U$20519 ( \20862 , \20860 );
and \U$20520 ( \20863 , \20862 , \5322 );
nor \U$20521 ( \20864 , \20861 , \20863 );
and \U$20522 ( \20865 , \20857 , \20864 );
and \U$20523 ( \20866 , \20849 , \20856 );
or \U$20524 ( \20867 , \20865 , \20866 );
xor \U$20525 ( \20868 , \20841 , \20867 );
and \U$20526 ( \20869 , \5881 , RI9871140_113);
and \U$20527 ( \20870 , RI9871320_117, \5879 );
nor \U$20528 ( \20871 , \20869 , \20870 );
and \U$20529 ( \20872 , \20871 , \5594 );
not \U$20530 ( \20873 , \20871 );
and \U$20531 ( \20874 , \20873 , \5885 );
nor \U$20532 ( \20875 , \20872 , \20874 );
and \U$20533 ( \20876 , \6453 , RI9871410_119);
and \U$20534 ( \20877 , RI98716e0_125, \6451 );
nor \U$20535 ( \20878 , \20876 , \20877 );
and \U$20536 ( \20879 , \20878 , \6190 );
not \U$20537 ( \20880 , \20878 );
and \U$20538 ( \20881 , \20880 , \6705 );
nor \U$20539 ( \20882 , \20879 , \20881 );
xor \U$20540 ( \20883 , \20875 , \20882 );
and \U$20541 ( \20884 , \7079 , RI98717d0_127);
and \U$20542 ( \20885 , RI9871500_121, \7077 );
nor \U$20543 ( \20886 , \20884 , \20885 );
and \U$20544 ( \20887 , \20886 , \6710 );
not \U$20545 ( \20888 , \20886 );
and \U$20546 ( \20889 , \20888 , \6709 );
nor \U$20547 ( \20890 , \20887 , \20889 );
and \U$20548 ( \20891 , \20883 , \20890 );
and \U$20549 ( \20892 , \20875 , \20882 );
or \U$20550 ( \20893 , \20891 , \20892 );
and \U$20551 ( \20894 , \20868 , \20893 );
and \U$20552 ( \20895 , \20841 , \20867 );
or \U$20553 ( \20896 , \20894 , \20895 );
and \U$20554 ( \20897 , \13045 , RI986e440_17);
and \U$20555 ( \20898 , RI986e710_23, \13043 );
nor \U$20556 ( \20899 , \20897 , \20898 );
and \U$20557 ( \20900 , \20899 , \13047 );
not \U$20558 ( \20901 , \20899 );
and \U$20559 ( \20902 , \20901 , \12619 );
nor \U$20560 ( \20903 , \20900 , \20902 );
and \U$20561 ( \20904 , \12293 , RI986f160_45);
and \U$20562 ( \20905 , RI986e530_19, \12291 );
nor \U$20563 ( \20906 , \20904 , \20905 );
and \U$20564 ( \20907 , \20906 , \11687 );
not \U$20565 ( \20908 , \20906 );
and \U$20566 ( \20909 , \20908 , \11686 );
nor \U$20567 ( \20910 , \20907 , \20909 );
xor \U$20568 ( \20911 , \20903 , \20910 );
and \U$20569 ( \20912 , \13882 , RI986e620_21);
and \U$20570 ( \20913 , RI986f7f0_59, \13880 );
nor \U$20571 ( \20914 , \20912 , \20913 );
and \U$20572 ( \20915 , \20914 , \13358 );
not \U$20573 ( \20916 , \20914 );
and \U$20574 ( \20917 , \20916 , \13359 );
nor \U$20575 ( \20918 , \20915 , \20917 );
and \U$20576 ( \20919 , \20911 , \20918 );
and \U$20577 ( \20920 , \20903 , \20910 );
or \U$20578 ( \20921 , \20919 , \20920 );
not \U$20579 ( \20922 , RI9873558_190);
and \U$20580 ( \20923 , \15780 , RI986f8e0_61);
and \U$20581 ( \20924 , RI9873648_192, RI986f430_51);
nor \U$20582 ( \20925 , \20923 , \20924 );
not \U$20583 ( \20926 , \20925 );
or \U$20584 ( \20927 , \20922 , \20926 );
or \U$20585 ( \20928 , \20925 , RI9873558_190);
nand \U$20586 ( \20929 , \20927 , \20928 );
xor \U$20587 ( \20930 , \20929 , \443 );
and \U$20588 ( \20931 , \14937 , RI986f700_57);
and \U$20589 ( \20932 , RI986f9d0_63, \14935 );
nor \U$20590 ( \20933 , \20931 , \20932 );
and \U$20591 ( \20934 , \20933 , \14539 );
not \U$20592 ( \20935 , \20933 );
and \U$20593 ( \20936 , \20935 , \14538 );
nor \U$20594 ( \20937 , \20934 , \20936 );
and \U$20595 ( \20938 , \20930 , \20937 );
and \U$20596 ( \20939 , \20929 , \443 );
or \U$20597 ( \20940 , \20938 , \20939 );
xor \U$20598 ( \20941 , \20921 , \20940 );
and \U$20599 ( \20942 , \10424 , RI986ecb0_35);
and \U$20600 ( \20943 , RI986f070_43, \10422 );
nor \U$20601 ( \20944 , \20942 , \20943 );
and \U$20602 ( \20945 , \20944 , \9840 );
not \U$20603 ( \20946 , \20944 );
and \U$20604 ( \20947 , \20946 , \10428 );
nor \U$20605 ( \20948 , \20945 , \20947 );
and \U$20606 ( \20949 , \9505 , RI986eda0_37);
and \U$20607 ( \20950 , RI986ebc0_33, \9503 );
nor \U$20608 ( \20951 , \20949 , \20950 );
and \U$20609 ( \20952 , \20951 , \9510 );
not \U$20610 ( \20953 , \20951 );
and \U$20611 ( \20954 , \20953 , \9513 );
nor \U$20612 ( \20955 , \20952 , \20954 );
xor \U$20613 ( \20956 , \20948 , \20955 );
and \U$20614 ( \20957 , \11696 , RI986ef80_41);
and \U$20615 ( \20958 , RI986f250_47, \11694 );
nor \U$20616 ( \20959 , \20957 , \20958 );
and \U$20617 ( \20960 , \20959 , \10965 );
not \U$20618 ( \20961 , \20959 );
and \U$20619 ( \20962 , \20961 , \11702 );
nor \U$20620 ( \20963 , \20960 , \20962 );
and \U$20621 ( \20964 , \20956 , \20963 );
and \U$20622 ( \20965 , \20948 , \20955 );
or \U$20623 ( \20966 , \20964 , \20965 );
and \U$20624 ( \20967 , \20941 , \20966 );
and \U$20625 ( \20968 , \20921 , \20940 );
or \U$20626 ( \20969 , \20967 , \20968 );
xor \U$20627 ( \20970 , \20896 , \20969 );
and \U$20628 ( \20971 , \2274 , RI986fca0_69);
and \U$20629 ( \20972 , RI986ff70_75, \2272 );
nor \U$20630 ( \20973 , \20971 , \20972 );
and \U$20631 ( \20974 , \20973 , \2030 );
not \U$20632 ( \20975 , \20973 );
and \U$20633 ( \20976 , \20975 , \2031 );
nor \U$20634 ( \20977 , \20974 , \20976 );
and \U$20635 ( \20978 , \1311 , RI98707e0_93);
and \U$20636 ( \20979 , RI986fac0_65, \1309 );
nor \U$20637 ( \20980 , \20978 , \20979 );
and \U$20638 ( \20981 , \20980 , \1458 );
not \U$20639 ( \20982 , \20980 );
and \U$20640 ( \20983 , \20982 , \1318 );
nor \U$20641 ( \20984 , \20981 , \20983 );
xor \U$20642 ( \20985 , \20977 , \20984 );
not \U$20643 ( \20986 , \2034 );
and \U$20644 ( \20987 , \2042 , RI986fbb0_67);
and \U$20645 ( \20988 , RI986fd90_71, \2040 );
nor \U$20646 ( \20989 , \20987 , \20988 );
not \U$20647 ( \20990 , \20989 );
or \U$20648 ( \20991 , \20986 , \20990 );
or \U$20649 ( \20992 , \20989 , \1462 );
nand \U$20650 ( \20993 , \20991 , \20992 );
and \U$20651 ( \20994 , \20985 , \20993 );
and \U$20652 ( \20995 , \20977 , \20984 );
or \U$20653 ( \20996 , \20994 , \20995 );
and \U$20654 ( \20997 , \776 , RI9870510_87);
and \U$20655 ( \20998 , RI9870330_83, \774 );
nor \U$20656 ( \20999 , \20997 , \20998 );
and \U$20657 ( \21000 , \20999 , \474 );
not \U$20658 ( \21001 , \20999 );
and \U$20659 ( \21002 , \21001 , \451 );
nor \U$20660 ( \21003 , \21000 , \21002 );
not \U$20661 ( \21004 , \1128 );
and \U$20662 ( \21005 , \1293 , RI9870240_81);
and \U$20663 ( \21006 , RI98706f0_91, \1291 );
nor \U$20664 ( \21007 , \21005 , \21006 );
not \U$20665 ( \21008 , \21007 );
or \U$20666 ( \21009 , \21004 , \21008 );
or \U$20667 ( \21010 , \21007 , \1301 );
nand \U$20668 ( \21011 , \21009 , \21010 );
xor \U$20669 ( \21012 , \21003 , \21011 );
and \U$20670 ( \21013 , \1329 , RI9870600_89);
and \U$20671 ( \21014 , RI98708d0_95, \1327 );
nor \U$20672 ( \21015 , \21013 , \21014 );
and \U$20673 ( \21016 , \21015 , \1336 );
not \U$20674 ( \21017 , \21015 );
and \U$20675 ( \21018 , \21017 , \1337 );
nor \U$20676 ( \21019 , \21016 , \21018 );
and \U$20677 ( \21020 , \21012 , \21019 );
and \U$20678 ( \21021 , \21003 , \21011 );
or \U$20679 ( \21022 , \21020 , \21021 );
xor \U$20680 ( \21023 , \20996 , \21022 );
not \U$20681 ( \21024 , \3918 );
and \U$20682 ( \21025 , \3683 , RI9870ab0_99);
and \U$20683 ( \21026 , RI9870d80_105, \3681 );
nor \U$20684 ( \21027 , \21025 , \21026 );
not \U$20685 ( \21028 , \21027 );
or \U$20686 ( \21029 , \21024 , \21028 );
or \U$20687 ( \21030 , \21027 , \3918 );
nand \U$20688 ( \21031 , \21029 , \21030 );
and \U$20689 ( \21032 , \2464 , RI986fe80_73);
and \U$20690 ( \21033 , RI9870060_77, \2462 );
nor \U$20691 ( \21034 , \21032 , \21033 );
and \U$20692 ( \21035 , \21034 , \2468 );
not \U$20693 ( \21036 , \21034 );
and \U$20694 ( \21037 , \21036 , \2263 );
nor \U$20695 ( \21038 , \21035 , \21037 );
xor \U$20696 ( \21039 , \21031 , \21038 );
not \U$20697 ( \21040 , \3406 );
and \U$20698 ( \21041 , \3254 , RI9870150_79);
and \U$20699 ( \21042 , RI9870f60_109, \3252 );
nor \U$20700 ( \21043 , \21041 , \21042 );
not \U$20701 ( \21044 , \21043 );
or \U$20702 ( \21045 , \21040 , \21044 );
or \U$20703 ( \21046 , \21043 , \3406 );
nand \U$20704 ( \21047 , \21045 , \21046 );
and \U$20705 ( \21048 , \21039 , \21047 );
and \U$20706 ( \21049 , \21031 , \21038 );
or \U$20707 ( \21050 , \21048 , \21049 );
and \U$20708 ( \21051 , \21023 , \21050 );
and \U$20709 ( \21052 , \20996 , \21022 );
or \U$20710 ( \21053 , \21051 , \21052 );
and \U$20711 ( \21054 , \20970 , \21053 );
and \U$20712 ( \21055 , \20896 , \20969 );
or \U$20713 ( \21056 , \21054 , \21055 );
xor \U$20714 ( \21057 , \20816 , \21056 );
xor \U$20715 ( \21058 , \20431 , \20438 );
xor \U$20716 ( \21059 , \21058 , \20446 );
xor \U$20717 ( \21060 , \20482 , \20490 );
xor \U$20718 ( \21061 , \21060 , \20498 );
xor \U$20719 ( \21062 , \21059 , \21061 );
xor \U$20720 ( \21063 , \20456 , \20463 );
xor \U$20721 ( \21064 , \21063 , \20471 );
and \U$20722 ( \21065 , \21062 , \21064 );
and \U$20723 ( \21066 , \21059 , \21061 );
or \U$20724 ( \21067 , \21065 , \21066 );
xor \U$20725 ( \21068 , \20402 , \20409 );
xor \U$20726 ( \21069 , \21068 , \20418 );
xor \U$20727 ( \21070 , \20375 , \20382 );
xor \U$20728 ( \21071 , \21070 , \20391 );
and \U$20729 ( \21072 , \21069 , \21071 );
xor \U$20730 ( \21073 , \20349 , \20356 );
xor \U$20731 ( \21074 , \21073 , \20365 );
xor \U$20732 ( \21075 , \20375 , \20382 );
xor \U$20733 ( \21076 , \21075 , \20391 );
and \U$20734 ( \21077 , \21074 , \21076 );
and \U$20735 ( \21078 , \21069 , \21074 );
or \U$20736 ( \21079 , \21072 , \21077 , \21078 );
xor \U$20737 ( \21080 , \21067 , \21079 );
xor \U$20738 ( \21081 , \20538 , \20545 );
xor \U$20739 ( \21082 , \21081 , \20554 );
xor \U$20740 ( \21083 , \20565 , \20572 );
xor \U$20741 ( \21084 , \21083 , \20580 );
and \U$20742 ( \21085 , \21082 , \21084 );
xor \U$20743 ( \21086 , \20512 , \20519 );
xor \U$20744 ( \21087 , \21086 , \20527 );
xor \U$20745 ( \21088 , \20565 , \20572 );
xor \U$20746 ( \21089 , \21088 , \20580 );
and \U$20747 ( \21090 , \21087 , \21089 );
and \U$20748 ( \21091 , \21082 , \21087 );
or \U$20749 ( \21092 , \21085 , \21090 , \21091 );
and \U$20750 ( \21093 , \21080 , \21092 );
and \U$20751 ( \21094 , \21067 , \21079 );
or \U$20752 ( \21095 , \21093 , \21094 );
and \U$20753 ( \21096 , \21057 , \21095 );
and \U$20754 ( \21097 , \20816 , \21056 );
or \U$20755 ( \21098 , \21096 , \21097 );
xor \U$20756 ( \21099 , \20734 , \20753 );
xor \U$20757 ( \21100 , \21099 , \20779 );
not \U$20758 ( \21101 , \21100 );
xor \U$20759 ( \21102 , \20530 , \20557 );
xor \U$20760 ( \21103 , \21102 , \20583 );
xor \U$20761 ( \21104 , \20449 , \20474 );
xor \U$20762 ( \21105 , \21104 , \20501 );
and \U$20763 ( \21106 , \21103 , \21105 );
not \U$20764 ( \21107 , \21106 );
or \U$20765 ( \21108 , \21101 , \21107 );
or \U$20766 ( \21109 , \21106 , \21100 );
xor \U$20767 ( \21110 , \20368 , \20394 );
xor \U$20768 ( \21111 , \21110 , \20421 );
xor \U$20769 ( \21112 , \20607 , \20614 );
xor \U$20770 ( \21113 , \21112 , \20617 );
xor \U$20771 ( \21114 , \21111 , \21113 );
not \U$20772 ( \21115 , \20591 );
xor \U$20773 ( \21116 , \20599 , \20594 );
not \U$20774 ( \21117 , \21116 );
or \U$20775 ( \21118 , \21115 , \21117 );
or \U$20776 ( \21119 , \21116 , \20591 );
nand \U$20777 ( \21120 , \21118 , \21119 );
and \U$20778 ( \21121 , \21114 , \21120 );
and \U$20779 ( \21122 , \21111 , \21113 );
or \U$20780 ( \21123 , \21121 , \21122 );
nand \U$20781 ( \21124 , \21109 , \21123 );
nand \U$20782 ( \21125 , \21108 , \21124 );
xor \U$20783 ( \21126 , \21098 , \21125 );
xor \U$20784 ( \21127 , \20601 , \20620 );
xor \U$20785 ( \21128 , \21127 , \20655 );
xor \U$20786 ( \21129 , \20197 , \20283 );
xor \U$20787 ( \21130 , \21129 , \20306 );
xor \U$20788 ( \21131 , \21128 , \21130 );
xor \U$20789 ( \21132 , \20675 , \20677 );
xor \U$20790 ( \21133 , \21132 , \20698 );
and \U$20791 ( \21134 , \21131 , \21133 );
and \U$20792 ( \21135 , \21128 , \21130 );
nor \U$20793 ( \21136 , \21134 , \21135 );
and \U$20794 ( \21137 , \21126 , \21136 );
and \U$20795 ( \21138 , \21098 , \21125 );
or \U$20796 ( \21139 , \21137 , \21138 );
xor \U$20797 ( \21140 , \20802 , \21139 );
not \U$20798 ( \21141 , \20069 );
not \U$20799 ( \21142 , \20063 );
or \U$20800 ( \21143 , \21141 , \21142 );
or \U$20801 ( \21144 , \20063 , \20069 );
nand \U$20802 ( \21145 , \21143 , \21144 );
not \U$20803 ( \21146 , \21145 );
not \U$20804 ( \21147 , \20061 );
and \U$20805 ( \21148 , \21146 , \21147 );
and \U$20806 ( \21149 , \21145 , \20061 );
nor \U$20807 ( \21150 , \21148 , \21149 );
not \U$20808 ( \21151 , \21150 );
xnor \U$20809 ( \21152 , \19430 , \19458 );
not \U$20810 ( \21153 , \21152 );
not \U$20811 ( \21154 , \19404 );
and \U$20812 ( \21155 , \21153 , \21154 );
and \U$20813 ( \21156 , \21152 , \19404 );
nor \U$20814 ( \21157 , \21155 , \21156 );
xor \U$20815 ( \21158 , \20316 , \20326 );
and \U$20816 ( \21159 , \21158 , \20337 );
and \U$20817 ( \21160 , \20316 , \20326 );
or \U$20818 ( \21161 , \21159 , \21160 );
xor \U$20819 ( \21162 , \21157 , \21161 );
not \U$20820 ( \21163 , \21162 );
or \U$20821 ( \21164 , \21151 , \21163 );
or \U$20822 ( \21165 , \21162 , \21150 );
nand \U$20823 ( \21166 , \21164 , \21165 );
xor \U$20824 ( \21167 , \20712 , \20718 );
and \U$20825 ( \21168 , \21167 , \20725 );
and \U$20826 ( \21169 , \20712 , \20718 );
or \U$20827 ( \21170 , \21168 , \21169 );
xor \U$20828 ( \21171 , \20730 , \20782 );
and \U$20829 ( \21172 , \21171 , \20789 );
and \U$20830 ( \21173 , \20730 , \20782 );
or \U$20831 ( \21174 , \21172 , \21173 );
xor \U$20832 ( \21175 , \21170 , \21174 );
xor \U$20833 ( \21176 , \19752 , \19754 );
xor \U$20834 ( \21177 , \21176 , \19757 );
and \U$20835 ( \21178 , \20794 , \21177 );
xor \U$20836 ( \21179 , \19752 , \19754 );
xor \U$20837 ( \21180 , \21179 , \19757 );
and \U$20838 ( \21181 , \20796 , \21180 );
and \U$20839 ( \21182 , \20794 , \20796 );
or \U$20840 ( \21183 , \21178 , \21181 , \21182 );
xor \U$20841 ( \21184 , \21175 , \21183 );
xor \U$20842 ( \21185 , \21166 , \21184 );
xor \U$20843 ( \21186 , \19729 , \19749 );
xor \U$20844 ( \21187 , \21186 , \19760 );
xor \U$20845 ( \21188 , \19847 , \19927 );
xor \U$20846 ( \21189 , \21188 , \20011 );
xor \U$20847 ( \21190 , \19551 , \19553 );
xor \U$20848 ( \21191 , \21190 , \19556 );
xor \U$20849 ( \21192 , \20019 , \20026 );
xor \U$20850 ( \21193 , \21191 , \21192 );
xor \U$20851 ( \21194 , \21189 , \21193 );
xor \U$20852 ( \21195 , \21187 , \21194 );
xor \U$20853 ( \21196 , \21185 , \21195 );
xor \U$20854 ( \21197 , \21140 , \21196 );
or \U$20855 ( \21198 , \20338 , \20115 );
not \U$20856 ( \21199 , \20115 );
not \U$20857 ( \21200 , \20338 );
or \U$20858 ( \21201 , \21199 , \21200 );
nand \U$20859 ( \21202 , \21201 , \20309 );
nand \U$20860 ( \21203 , \21198 , \21202 );
xor \U$20861 ( \21204 , \20589 , \20658 );
and \U$20862 ( \21205 , \21204 , \20701 );
and \U$20863 ( \21206 , \20589 , \20658 );
nor \U$20864 ( \21207 , \21205 , \21206 );
xor \U$20865 ( \21208 , \21203 , \21207 );
xor \U$20866 ( \21209 , \20712 , \20718 );
xor \U$20867 ( \21210 , \21209 , \20725 );
and \U$20868 ( \21211 , \20790 , \21210 );
xor \U$20869 ( \21212 , \20712 , \20718 );
xor \U$20870 ( \21213 , \21212 , \20725 );
and \U$20871 ( \21214 , \20798 , \21213 );
and \U$20872 ( \21215 , \20790 , \20798 );
or \U$20873 ( \21216 , \21211 , \21214 , \21215 );
xor \U$20874 ( \21217 , \21208 , \21216 );
xor \U$20875 ( \21218 , \21197 , \21217 );
xnor \U$20876 ( \21219 , \20702 , \20342 );
not \U$20877 ( \21220 , \21219 );
not \U$20878 ( \21221 , \20800 );
and \U$20879 ( \21222 , \21220 , \21221 );
and \U$20880 ( \21223 , \21219 , \20800 );
nor \U$20881 ( \21224 , \21222 , \21223 );
xnor \U$20882 ( \21225 , \21123 , \21106 );
not \U$20883 ( \21226 , \21225 );
not \U$20884 ( \21227 , \21100 );
and \U$20885 ( \21228 , \21226 , \21227 );
and \U$20886 ( \21229 , \21225 , \21100 );
nor \U$20887 ( \21230 , \21228 , \21229 );
xor \U$20888 ( \21231 , \20424 , \20504 );
xor \U$20889 ( \21232 , \21231 , \20586 );
xor \U$20890 ( \21233 , \21230 , \21232 );
xor \U$20891 ( \21234 , \21128 , \21130 );
xor \U$20892 ( \21235 , \21234 , \21133 );
and \U$20893 ( \21236 , \21233 , \21235 );
and \U$20894 ( \21237 , \21230 , \21232 );
or \U$20895 ( \21238 , \21236 , \21237 );
or \U$20896 ( \21239 , \21224 , \21238 );
not \U$20897 ( \21240 , \21238 );
not \U$20898 ( \21241 , \21224 );
or \U$20899 ( \21242 , \21240 , \21241 );
xor \U$20900 ( \21243 , \20896 , \20969 );
xor \U$20901 ( \21244 , \21243 , \21053 );
xor \U$20902 ( \21245 , \20742 , \456 );
xor \U$20903 ( \21246 , \21245 , \20750 );
xor \U$20904 ( \21247 , \20804 , \20811 );
xor \U$20905 ( \21248 , \21246 , \21247 );
xor \U$20906 ( \21249 , \21244 , \21248 );
xor \U$20907 ( \21250 , \21067 , \21079 );
xor \U$20908 ( \21251 , \21250 , \21092 );
and \U$20909 ( \21252 , \21249 , \21251 );
and \U$20910 ( \21253 , \21244 , \21248 );
or \U$20911 ( \21254 , \21252 , \21253 );
xor \U$20912 ( \21255 , \20849 , \20856 );
xor \U$20913 ( \21256 , \21255 , \20864 );
xor \U$20914 ( \21257 , \21031 , \21038 );
xor \U$20915 ( \21258 , \21257 , \21047 );
xor \U$20916 ( \21259 , \21256 , \21258 );
xor \U$20917 ( \21260 , \20875 , \20882 );
xor \U$20918 ( \21261 , \21260 , \20890 );
and \U$20919 ( \21262 , \21259 , \21261 );
and \U$20920 ( \21263 , \21256 , \21258 );
or \U$20921 ( \21264 , \21262 , \21263 );
nand \U$20922 ( \21265 , RI9870420_85, \436 );
and \U$20923 ( \21266 , \21265 , \444 );
not \U$20924 ( \21267 , \21265 );
and \U$20925 ( \21268 , \21267 , \443 );
nor \U$20926 ( \21269 , \21266 , \21268 );
xor \U$20927 ( \21270 , \20977 , \20984 );
xor \U$20928 ( \21271 , \21270 , \20993 );
and \U$20929 ( \21272 , \21269 , \21271 );
xor \U$20930 ( \21273 , \21003 , \21011 );
xor \U$20931 ( \21274 , \21273 , \21019 );
xor \U$20932 ( \21275 , \20977 , \20984 );
xor \U$20933 ( \21276 , \21275 , \20993 );
and \U$20934 ( \21277 , \21274 , \21276 );
and \U$20935 ( \21278 , \21269 , \21274 );
or \U$20936 ( \21279 , \21272 , \21277 , \21278 );
xor \U$20937 ( \21280 , \21264 , \21279 );
xor \U$20938 ( \21281 , \20823 , \20830 );
xor \U$20939 ( \21282 , \21281 , \20838 );
xor \U$20940 ( \21283 , \20903 , \20910 );
xor \U$20941 ( \21284 , \21283 , \20918 );
and \U$20942 ( \21285 , \21282 , \21284 );
xor \U$20943 ( \21286 , \20948 , \20955 );
xor \U$20944 ( \21287 , \21286 , \20963 );
xor \U$20945 ( \21288 , \20903 , \20910 );
xor \U$20946 ( \21289 , \21288 , \20918 );
and \U$20947 ( \21290 , \21287 , \21289 );
and \U$20948 ( \21291 , \21282 , \21287 );
or \U$20949 ( \21292 , \21285 , \21290 , \21291 );
and \U$20950 ( \21293 , \21280 , \21292 );
and \U$20951 ( \21294 , \21264 , \21279 );
or \U$20952 ( \21295 , \21293 , \21294 );
and \U$20953 ( \21296 , \9237 , RI986e8f0_27);
and \U$20954 ( \21297 , RI986e800_25, \9235 );
nor \U$20955 ( \21298 , \21296 , \21297 );
and \U$20956 ( \21299 , \21298 , \9241 );
not \U$20957 ( \21300 , \21298 );
and \U$20958 ( \21301 , \21300 , \8836 );
nor \U$20959 ( \21302 , \21299 , \21301 );
and \U$20960 ( \21303 , \9505 , RI986ee90_39);
and \U$20961 ( \21304 , RI986eda0_37, \9503 );
nor \U$20962 ( \21305 , \21303 , \21304 );
and \U$20963 ( \21306 , \21305 , \9510 );
not \U$20964 ( \21307 , \21305 );
and \U$20965 ( \21308 , \21307 , \9513 );
nor \U$20966 ( \21309 , \21306 , \21308 );
xor \U$20967 ( \21310 , \21302 , \21309 );
and \U$20968 ( \21311 , \10424 , RI986ebc0_33);
and \U$20969 ( \21312 , RI986ecb0_35, \10422 );
nor \U$20970 ( \21313 , \21311 , \21312 );
and \U$20971 ( \21314 , \21313 , \9840 );
not \U$20972 ( \21315 , \21313 );
and \U$20973 ( \21316 , \21315 , \10428 );
nor \U$20974 ( \21317 , \21314 , \21316 );
and \U$20975 ( \21318 , \21310 , \21317 );
and \U$20976 ( \21319 , \21302 , \21309 );
or \U$20977 ( \21320 , \21318 , \21319 );
and \U$20978 ( \21321 , \14937 , RI986f7f0_59);
and \U$20979 ( \21322 , RI986f700_57, \14935 );
nor \U$20980 ( \21323 , \21321 , \21322 );
and \U$20981 ( \21324 , \21323 , \14539 );
not \U$20982 ( \21325 , \21323 );
and \U$20983 ( \21326 , \21325 , \14538 );
nor \U$20984 ( \21327 , \21324 , \21326 );
not \U$20985 ( \21328 , RI9873558_190);
and \U$20986 ( \21329 , \15780 , RI986f9d0_63);
and \U$20987 ( \21330 , RI9873648_192, RI986f8e0_61);
nor \U$20988 ( \21331 , \21329 , \21330 );
not \U$20989 ( \21332 , \21331 );
or \U$20990 ( \21333 , \21328 , \21332 );
or \U$20991 ( \21334 , \21331 , RI9873558_190);
nand \U$20992 ( \21335 , \21333 , \21334 );
xor \U$20993 ( \21336 , \21327 , \21335 );
and \U$20994 ( \21337 , \13882 , RI986e710_23);
and \U$20995 ( \21338 , RI986e620_21, \13880 );
nor \U$20996 ( \21339 , \21337 , \21338 );
and \U$20997 ( \21340 , \21339 , \13358 );
not \U$20998 ( \21341 , \21339 );
and \U$20999 ( \21342 , \21341 , \13359 );
nor \U$21000 ( \21343 , \21340 , \21342 );
and \U$21001 ( \21344 , \21336 , \21343 );
and \U$21002 ( \21345 , \21327 , \21335 );
or \U$21003 ( \21346 , \21344 , \21345 );
xor \U$21004 ( \21347 , \21320 , \21346 );
and \U$21005 ( \21348 , \11696 , RI986f070_43);
and \U$21006 ( \21349 , RI986ef80_41, \11694 );
nor \U$21007 ( \21350 , \21348 , \21349 );
and \U$21008 ( \21351 , \21350 , \10965 );
not \U$21009 ( \21352 , \21350 );
and \U$21010 ( \21353 , \21352 , \11702 );
nor \U$21011 ( \21354 , \21351 , \21353 );
and \U$21012 ( \21355 , \12293 , RI986f250_47);
and \U$21013 ( \21356 , RI986f160_45, \12291 );
nor \U$21014 ( \21357 , \21355 , \21356 );
and \U$21015 ( \21358 , \21357 , \11687 );
not \U$21016 ( \21359 , \21357 );
and \U$21017 ( \21360 , \21359 , \11686 );
nor \U$21018 ( \21361 , \21358 , \21360 );
xor \U$21019 ( \21362 , \21354 , \21361 );
and \U$21020 ( \21363 , \13045 , RI986e530_19);
and \U$21021 ( \21364 , RI986e440_17, \13043 );
nor \U$21022 ( \21365 , \21363 , \21364 );
and \U$21023 ( \21366 , \21365 , \13047 );
not \U$21024 ( \21367 , \21365 );
and \U$21025 ( \21368 , \21367 , \12619 );
nor \U$21026 ( \21369 , \21366 , \21368 );
and \U$21027 ( \21370 , \21362 , \21369 );
and \U$21028 ( \21371 , \21354 , \21361 );
or \U$21029 ( \21372 , \21370 , \21371 );
and \U$21030 ( \21373 , \21347 , \21372 );
and \U$21031 ( \21374 , \21320 , \21346 );
or \U$21032 ( \21375 , \21373 , \21374 );
and \U$21033 ( \21376 , \1329 , RI98706f0_91);
and \U$21034 ( \21377 , RI9870600_89, \1327 );
nor \U$21035 ( \21378 , \21376 , \21377 );
and \U$21036 ( \21379 , \21378 , \1336 );
not \U$21037 ( \21380 , \21378 );
and \U$21038 ( \21381 , \21380 , \1337 );
nor \U$21039 ( \21382 , \21379 , \21381 );
and \U$21040 ( \21383 , \1311 , RI98708d0_95);
and \U$21041 ( \21384 , RI98707e0_93, \1309 );
nor \U$21042 ( \21385 , \21383 , \21384 );
and \U$21043 ( \21386 , \21385 , \1458 );
not \U$21044 ( \21387 , \21385 );
and \U$21045 ( \21388 , \21387 , \1318 );
nor \U$21046 ( \21389 , \21386 , \21388 );
xor \U$21047 ( \21390 , \21382 , \21389 );
not \U$21048 ( \21391 , \1462 );
and \U$21049 ( \21392 , \2042 , RI986fac0_65);
and \U$21050 ( \21393 , RI986fbb0_67, \2040 );
nor \U$21051 ( \21394 , \21392 , \21393 );
not \U$21052 ( \21395 , \21394 );
or \U$21053 ( \21396 , \21391 , \21395 );
or \U$21054 ( \21397 , \21394 , \2034 );
nand \U$21055 ( \21398 , \21396 , \21397 );
and \U$21056 ( \21399 , \21390 , \21398 );
and \U$21057 ( \21400 , \21382 , \21389 );
or \U$21058 ( \21401 , \21399 , \21400 );
not \U$21059 ( \21402 , \1301 );
and \U$21060 ( \21403 , \1293 , RI9870330_83);
and \U$21061 ( \21404 , RI9870240_81, \1291 );
nor \U$21062 ( \21405 , \21403 , \21404 );
not \U$21063 ( \21406 , \21405 );
or \U$21064 ( \21407 , \21402 , \21406 );
or \U$21065 ( \21408 , \21405 , \1128 );
nand \U$21066 ( \21409 , \21407 , \21408 );
and \U$21067 ( \21410 , \776 , RI9870420_85);
and \U$21068 ( \21411 , RI9870510_87, \774 );
nor \U$21069 ( \21412 , \21410 , \21411 );
and \U$21070 ( \21413 , \21412 , \474 );
not \U$21071 ( \21414 , \21412 );
and \U$21072 ( \21415 , \21414 , \451 );
nor \U$21073 ( \21416 , \21413 , \21415 );
and \U$21074 ( \21417 , \21409 , \21416 );
xor \U$21075 ( \21418 , \21401 , \21417 );
and \U$21076 ( \21419 , \2274 , RI986fd90_71);
and \U$21077 ( \21420 , RI986fca0_69, \2272 );
nor \U$21078 ( \21421 , \21419 , \21420 );
and \U$21079 ( \21422 , \21421 , \2030 );
not \U$21080 ( \21423 , \21421 );
and \U$21081 ( \21424 , \21423 , \2031 );
nor \U$21082 ( \21425 , \21422 , \21424 );
and \U$21083 ( \21426 , \2464 , RI986ff70_75);
and \U$21084 ( \21427 , RI986fe80_73, \2462 );
nor \U$21085 ( \21428 , \21426 , \21427 );
and \U$21086 ( \21429 , \21428 , \2468 );
not \U$21087 ( \21430 , \21428 );
and \U$21088 ( \21431 , \21430 , \2263 );
nor \U$21089 ( \21432 , \21429 , \21431 );
xor \U$21090 ( \21433 , \21425 , \21432 );
not \U$21091 ( \21434 , \2935 );
and \U$21092 ( \21435 , \3254 , RI9870060_77);
and \U$21093 ( \21436 , RI9870150_79, \3252 );
nor \U$21094 ( \21437 , \21435 , \21436 );
not \U$21095 ( \21438 , \21437 );
or \U$21096 ( \21439 , \21434 , \21438 );
or \U$21097 ( \21440 , \21437 , \3406 );
nand \U$21098 ( \21441 , \21439 , \21440 );
and \U$21099 ( \21442 , \21433 , \21441 );
and \U$21100 ( \21443 , \21425 , \21432 );
or \U$21101 ( \21444 , \21442 , \21443 );
and \U$21102 ( \21445 , \21418 , \21444 );
and \U$21103 ( \21446 , \21401 , \21417 );
or \U$21104 ( \21447 , \21445 , \21446 );
xor \U$21105 ( \21448 , \21375 , \21447 );
and \U$21106 ( \21449 , \7079 , RI98716e0_125);
and \U$21107 ( \21450 , RI98717d0_127, \7077 );
nor \U$21108 ( \21451 , \21449 , \21450 );
and \U$21109 ( \21452 , \21451 , \6710 );
not \U$21110 ( \21453 , \21451 );
and \U$21111 ( \21454 , \21453 , \6709 );
nor \U$21112 ( \21455 , \21452 , \21454 );
and \U$21113 ( \21456 , \7729 , RI9871500_121);
and \U$21114 ( \21457 , RI98715f0_123, \7727 );
nor \U$21115 ( \21458 , \21456 , \21457 );
and \U$21116 ( \21459 , \21458 , \7480 );
not \U$21117 ( \21460 , \21458 );
and \U$21118 ( \21461 , \21460 , \7733 );
nor \U$21119 ( \21462 , \21459 , \21461 );
xor \U$21120 ( \21463 , \21455 , \21462 );
and \U$21121 ( \21464 , \8486 , RI986ead0_31);
and \U$21122 ( \21465 , RI986e9e0_29, \8484 );
nor \U$21123 ( \21466 , \21464 , \21465 );
and \U$21124 ( \21467 , \21466 , \8050 );
not \U$21125 ( \21468 , \21466 );
and \U$21126 ( \21469 , \21468 , \8051 );
nor \U$21127 ( \21470 , \21467 , \21469 );
and \U$21128 ( \21471 , \21463 , \21470 );
and \U$21129 ( \21472 , \21455 , \21462 );
or \U$21130 ( \21473 , \21471 , \21472 );
and \U$21131 ( \21474 , \5318 , RI9871050_111);
and \U$21132 ( \21475 , RI9870c90_103, \5316 );
nor \U$21133 ( \21476 , \21474 , \21475 );
and \U$21134 ( \21477 , \21476 , \5052 );
not \U$21135 ( \21478 , \21476 );
and \U$21136 ( \21479 , \21478 , \5322 );
nor \U$21137 ( \21480 , \21477 , \21479 );
and \U$21138 ( \21481 , \5881 , RI9871230_115);
and \U$21139 ( \21482 , RI9871140_113, \5879 );
nor \U$21140 ( \21483 , \21481 , \21482 );
and \U$21141 ( \21484 , \21483 , \5594 );
not \U$21142 ( \21485 , \21483 );
and \U$21143 ( \21486 , \21485 , \5885 );
nor \U$21144 ( \21487 , \21484 , \21486 );
xor \U$21145 ( \21488 , \21480 , \21487 );
and \U$21146 ( \21489 , \6453 , RI9871320_117);
and \U$21147 ( \21490 , RI9871410_119, \6451 );
nor \U$21148 ( \21491 , \21489 , \21490 );
and \U$21149 ( \21492 , \21491 , \6190 );
not \U$21150 ( \21493 , \21491 );
and \U$21151 ( \21494 , \21493 , \6705 );
nor \U$21152 ( \21495 , \21492 , \21494 );
and \U$21153 ( \21496 , \21488 , \21495 );
and \U$21154 ( \21497 , \21480 , \21487 );
or \U$21155 ( \21498 , \21496 , \21497 );
xor \U$21156 ( \21499 , \21473 , \21498 );
not \U$21157 ( \21500 , \3918 );
and \U$21158 ( \21501 , \3683 , RI9870f60_109);
and \U$21159 ( \21502 , RI9870ab0_99, \3681 );
nor \U$21160 ( \21503 , \21501 , \21502 );
not \U$21161 ( \21504 , \21503 );
or \U$21162 ( \21505 , \21500 , \21504 );
or \U$21163 ( \21506 , \21503 , \3412 );
nand \U$21164 ( \21507 , \21505 , \21506 );
and \U$21165 ( \21508 , \4203 , RI9870d80_105);
and \U$21166 ( \21509 , RI98709c0_97, \4201 );
nor \U$21167 ( \21510 , \21508 , \21509 );
and \U$21168 ( \21511 , \21510 , \4207 );
not \U$21169 ( \21512 , \21510 );
and \U$21170 ( \21513 , \21512 , \3923 );
nor \U$21171 ( \21514 , \21511 , \21513 );
xor \U$21172 ( \21515 , \21507 , \21514 );
not \U$21173 ( \21516 , \4519 );
and \U$21174 ( \21517 , \4710 , RI9870e70_107);
and \U$21175 ( \21518 , RI9870ba0_101, \4708 );
nor \U$21176 ( \21519 , \21517 , \21518 );
not \U$21177 ( \21520 , \21519 );
or \U$21178 ( \21521 , \21516 , \21520 );
or \U$21179 ( \21522 , \21519 , \4521 );
nand \U$21180 ( \21523 , \21521 , \21522 );
and \U$21181 ( \21524 , \21515 , \21523 );
and \U$21182 ( \21525 , \21507 , \21514 );
or \U$21183 ( \21526 , \21524 , \21525 );
and \U$21184 ( \21527 , \21499 , \21526 );
and \U$21185 ( \21528 , \21473 , \21498 );
or \U$21186 ( \21529 , \21527 , \21528 );
and \U$21187 ( \21530 , \21448 , \21529 );
and \U$21188 ( \21531 , \21375 , \21447 );
or \U$21189 ( \21532 , \21530 , \21531 );
xor \U$21190 ( \21533 , \21295 , \21532 );
xor \U$21191 ( \21534 , \20375 , \20382 );
xor \U$21192 ( \21535 , \21534 , \20391 );
xor \U$21193 ( \21536 , \21069 , \21074 );
xor \U$21194 ( \21537 , \21535 , \21536 );
xor \U$21195 ( \21538 , \21059 , \21061 );
xor \U$21196 ( \21539 , \21538 , \21064 );
and \U$21197 ( \21540 , \21537 , \21539 );
xor \U$21198 ( \21541 , \20565 , \20572 );
xor \U$21199 ( \21542 , \21541 , \20580 );
xor \U$21200 ( \21543 , \21082 , \21087 );
xor \U$21201 ( \21544 , \21542 , \21543 );
xor \U$21202 ( \21545 , \21059 , \21061 );
xor \U$21203 ( \21546 , \21545 , \21064 );
and \U$21204 ( \21547 , \21544 , \21546 );
and \U$21205 ( \21548 , \21537 , \21544 );
or \U$21206 ( \21549 , \21540 , \21547 , \21548 );
and \U$21207 ( \21550 , \21533 , \21549 );
and \U$21208 ( \21551 , \21295 , \21532 );
or \U$21209 ( \21552 , \21550 , \21551 );
xor \U$21210 ( \21553 , \21254 , \21552 );
xor \U$21211 ( \21554 , \20996 , \21022 );
xor \U$21212 ( \21555 , \21554 , \21050 );
xor \U$21213 ( \21556 , \20921 , \20940 );
xor \U$21214 ( \21557 , \21556 , \20966 );
xor \U$21215 ( \21558 , \21555 , \21557 );
xor \U$21216 ( \21559 , \20841 , \20867 );
xor \U$21217 ( \21560 , \21559 , \20893 );
and \U$21218 ( \21561 , \21558 , \21560 );
and \U$21219 ( \21562 , \21555 , \21557 );
or \U$21220 ( \21563 , \21561 , \21562 );
xor \U$21221 ( \21564 , \21103 , \21105 );
xor \U$21222 ( \21565 , \21563 , \21564 );
xor \U$21223 ( \21566 , \21111 , \21113 );
xor \U$21224 ( \21567 , \21566 , \21120 );
and \U$21225 ( \21568 , \21565 , \21567 );
and \U$21226 ( \21569 , \21563 , \21564 );
or \U$21227 ( \21570 , \21568 , \21569 );
and \U$21228 ( \21571 , \21553 , \21570 );
and \U$21229 ( \21572 , \21254 , \21552 );
or \U$21230 ( \21573 , \21571 , \21572 );
nand \U$21231 ( \21574 , \21242 , \21573 );
nand \U$21232 ( \21575 , \21239 , \21574 );
xor \U$21233 ( \21576 , \21218 , \21575 );
not \U$21234 ( \21577 , \21576 );
xor \U$21235 ( \21578 , \21098 , \21125 );
xor \U$21236 ( \21579 , \21578 , \21136 );
not \U$21237 ( \21580 , \21579 );
xor \U$21238 ( \21581 , \21230 , \21232 );
xor \U$21239 ( \21582 , \21581 , \21235 );
not \U$21240 ( \21583 , \21582 );
xor \U$21241 ( \21584 , \21254 , \21552 );
xor \U$21242 ( \21585 , \21584 , \21570 );
nand \U$21243 ( \21586 , \21583 , \21585 );
nand \U$21244 ( \21587 , \21580 , \21586 );
xor \U$21245 ( \21588 , \21327 , \21335 );
xor \U$21246 ( \21589 , \21588 , \21343 );
xor \U$21247 ( \21590 , \21302 , \21309 );
xor \U$21248 ( \21591 , \21590 , \21317 );
xor \U$21249 ( \21592 , \21589 , \21591 );
xor \U$21250 ( \21593 , \21354 , \21361 );
xor \U$21251 ( \21594 , \21593 , \21369 );
and \U$21252 ( \21595 , \21592 , \21594 );
and \U$21253 ( \21596 , \21589 , \21591 );
or \U$21254 ( \21597 , \21595 , \21596 );
xor \U$21255 ( \21598 , \21409 , \21416 );
xor \U$21256 ( \21599 , \21425 , \21432 );
xor \U$21257 ( \21600 , \21599 , \21441 );
and \U$21258 ( \21601 , \21598 , \21600 );
xor \U$21259 ( \21602 , \21382 , \21389 );
xor \U$21260 ( \21603 , \21602 , \21398 );
xor \U$21261 ( \21604 , \21425 , \21432 );
xor \U$21262 ( \21605 , \21604 , \21441 );
and \U$21263 ( \21606 , \21603 , \21605 );
and \U$21264 ( \21607 , \21598 , \21603 );
or \U$21265 ( \21608 , \21601 , \21606 , \21607 );
xor \U$21266 ( \21609 , \21597 , \21608 );
xor \U$21267 ( \21610 , \21507 , \21514 );
xor \U$21268 ( \21611 , \21610 , \21523 );
xor \U$21269 ( \21612 , \21455 , \21462 );
xor \U$21270 ( \21613 , \21612 , \21470 );
and \U$21271 ( \21614 , \21611 , \21613 );
xor \U$21272 ( \21615 , \21480 , \21487 );
xor \U$21273 ( \21616 , \21615 , \21495 );
xor \U$21274 ( \21617 , \21455 , \21462 );
xor \U$21275 ( \21618 , \21617 , \21470 );
and \U$21276 ( \21619 , \21616 , \21618 );
and \U$21277 ( \21620 , \21611 , \21616 );
or \U$21278 ( \21621 , \21614 , \21619 , \21620 );
and \U$21279 ( \21622 , \21609 , \21621 );
and \U$21280 ( \21623 , \21597 , \21608 );
or \U$21281 ( \21624 , \21622 , \21623 );
and \U$21282 ( \21625 , \2464 , RI986fca0_69);
and \U$21283 ( \21626 , RI986ff70_75, \2462 );
nor \U$21284 ( \21627 , \21625 , \21626 );
and \U$21285 ( \21628 , \21627 , \2468 );
not \U$21286 ( \21629 , \21627 );
and \U$21287 ( \21630 , \21629 , \2263 );
nor \U$21288 ( \21631 , \21628 , \21630 );
not \U$21289 ( \21632 , \3406 );
and \U$21290 ( \21633 , \3254 , RI986fe80_73);
and \U$21291 ( \21634 , RI9870060_77, \3252 );
nor \U$21292 ( \21635 , \21633 , \21634 );
not \U$21293 ( \21636 , \21635 );
or \U$21294 ( \21637 , \21632 , \21636 );
or \U$21295 ( \21638 , \21635 , \2935 );
nand \U$21296 ( \21639 , \21637 , \21638 );
xor \U$21297 ( \21640 , \21631 , \21639 );
not \U$21298 ( \21641 , \3412 );
and \U$21299 ( \21642 , \3683 , RI9870150_79);
and \U$21300 ( \21643 , RI9870f60_109, \3681 );
nor \U$21301 ( \21644 , \21642 , \21643 );
not \U$21302 ( \21645 , \21644 );
or \U$21303 ( \21646 , \21641 , \21645 );
or \U$21304 ( \21647 , \21644 , \3412 );
nand \U$21305 ( \21648 , \21646 , \21647 );
and \U$21306 ( \21649 , \21640 , \21648 );
and \U$21307 ( \21650 , \21631 , \21639 );
or \U$21308 ( \21651 , \21649 , \21650 );
and \U$21309 ( \21652 , \1329 , RI9870240_81);
and \U$21310 ( \21653 , RI98706f0_91, \1327 );
nor \U$21311 ( \21654 , \21652 , \21653 );
and \U$21312 ( \21655 , \21654 , \1336 );
not \U$21313 ( \21656 , \21654 );
and \U$21314 ( \21657 , \21656 , \1337 );
nor \U$21315 ( \21658 , \21655 , \21657 );
nand \U$21316 ( \21659 , RI9870420_85, \774 );
and \U$21317 ( \21660 , \21659 , \474 );
not \U$21318 ( \21661 , \21659 );
and \U$21319 ( \21662 , \21661 , \451 );
nor \U$21320 ( \21663 , \21660 , \21662 );
xor \U$21321 ( \21664 , \21658 , \21663 );
not \U$21322 ( \21665 , \1301 );
and \U$21323 ( \21666 , \1293 , RI9870510_87);
and \U$21324 ( \21667 , RI9870330_83, \1291 );
nor \U$21325 ( \21668 , \21666 , \21667 );
not \U$21326 ( \21669 , \21668 );
or \U$21327 ( \21670 , \21665 , \21669 );
or \U$21328 ( \21671 , \21668 , \1301 );
nand \U$21329 ( \21672 , \21670 , \21671 );
and \U$21330 ( \21673 , \21664 , \21672 );
and \U$21331 ( \21674 , \21658 , \21663 );
or \U$21332 ( \21675 , \21673 , \21674 );
xor \U$21333 ( \21676 , \21651 , \21675 );
and \U$21334 ( \21677 , \1311 , RI9870600_89);
and \U$21335 ( \21678 , RI98708d0_95, \1309 );
nor \U$21336 ( \21679 , \21677 , \21678 );
and \U$21337 ( \21680 , \21679 , \1458 );
not \U$21338 ( \21681 , \21679 );
and \U$21339 ( \21682 , \21681 , \1318 );
nor \U$21340 ( \21683 , \21680 , \21682 );
not \U$21341 ( \21684 , \1462 );
and \U$21342 ( \21685 , \2042 , RI98707e0_93);
and \U$21343 ( \21686 , RI986fac0_65, \2040 );
nor \U$21344 ( \21687 , \21685 , \21686 );
not \U$21345 ( \21688 , \21687 );
or \U$21346 ( \21689 , \21684 , \21688 );
or \U$21347 ( \21690 , \21687 , \2034 );
nand \U$21348 ( \21691 , \21689 , \21690 );
xor \U$21349 ( \21692 , \21683 , \21691 );
and \U$21350 ( \21693 , \2274 , RI986fbb0_67);
and \U$21351 ( \21694 , RI986fd90_71, \2272 );
nor \U$21352 ( \21695 , \21693 , \21694 );
and \U$21353 ( \21696 , \21695 , \2030 );
not \U$21354 ( \21697 , \21695 );
and \U$21355 ( \21698 , \21697 , \2031 );
nor \U$21356 ( \21699 , \21696 , \21698 );
and \U$21357 ( \21700 , \21692 , \21699 );
and \U$21358 ( \21701 , \21683 , \21691 );
or \U$21359 ( \21702 , \21700 , \21701 );
and \U$21360 ( \21703 , \21676 , \21702 );
and \U$21361 ( \21704 , \21651 , \21675 );
or \U$21362 ( \21705 , \21703 , \21704 );
and \U$21363 ( \21706 , \12293 , RI986ef80_41);
and \U$21364 ( \21707 , RI986f250_47, \12291 );
nor \U$21365 ( \21708 , \21706 , \21707 );
and \U$21366 ( \21709 , \21708 , \11686 );
not \U$21367 ( \21710 , \21708 );
and \U$21368 ( \21711 , \21710 , \11687 );
nor \U$21369 ( \21712 , \21709 , \21711 );
and \U$21370 ( \21713 , \13882 , RI986e440_17);
and \U$21371 ( \21714 , RI986e710_23, \13880 );
nor \U$21372 ( \21715 , \21713 , \21714 );
and \U$21373 ( \21716 , \21715 , \13359 );
not \U$21374 ( \21717 , \21715 );
and \U$21375 ( \21718 , \21717 , \13358 );
nor \U$21376 ( \21719 , \21716 , \21718 );
or \U$21377 ( \21720 , \21712 , \21719 );
not \U$21378 ( \21721 , \21719 );
not \U$21379 ( \21722 , \21712 );
or \U$21380 ( \21723 , \21721 , \21722 );
and \U$21381 ( \21724 , \13045 , RI986f160_45);
and \U$21382 ( \21725 , RI986e530_19, \13043 );
nor \U$21383 ( \21726 , \21724 , \21725 );
and \U$21384 ( \21727 , \21726 , \13047 );
not \U$21385 ( \21728 , \21726 );
and \U$21386 ( \21729 , \21728 , \12619 );
nor \U$21387 ( \21730 , \21727 , \21729 );
nand \U$21388 ( \21731 , \21723 , \21730 );
nand \U$21389 ( \21732 , \21720 , \21731 );
not \U$21390 ( \21733 , RI9873558_190);
and \U$21391 ( \21734 , \15780 , RI986f700_57);
and \U$21392 ( \21735 , RI9873648_192, RI986f9d0_63);
nor \U$21393 ( \21736 , \21734 , \21735 );
not \U$21394 ( \21737 , \21736 );
or \U$21395 ( \21738 , \21733 , \21737 );
or \U$21396 ( \21739 , \21736 , RI9873558_190);
nand \U$21397 ( \21740 , \21738 , \21739 );
xor \U$21398 ( \21741 , \21740 , \451 );
and \U$21399 ( \21742 , \14937 , RI986e620_21);
and \U$21400 ( \21743 , RI986f7f0_59, \14935 );
nor \U$21401 ( \21744 , \21742 , \21743 );
and \U$21402 ( \21745 , \21744 , \14539 );
not \U$21403 ( \21746 , \21744 );
and \U$21404 ( \21747 , \21746 , \14538 );
nor \U$21405 ( \21748 , \21745 , \21747 );
and \U$21406 ( \21749 , \21741 , \21748 );
and \U$21407 ( \21750 , \21740 , \451 );
or \U$21408 ( \21751 , \21749 , \21750 );
xor \U$21409 ( \21752 , \21732 , \21751 );
and \U$21410 ( \21753 , \9505 , RI986e800_25);
and \U$21411 ( \21754 , RI986ee90_39, \9503 );
nor \U$21412 ( \21755 , \21753 , \21754 );
and \U$21413 ( \21756 , \21755 , \9513 );
not \U$21414 ( \21757 , \21755 );
and \U$21415 ( \21758 , \21757 , \9510 );
nor \U$21416 ( \21759 , \21756 , \21758 );
and \U$21417 ( \21760 , \11696 , RI986ecb0_35);
and \U$21418 ( \21761 , RI986f070_43, \11694 );
nor \U$21419 ( \21762 , \21760 , \21761 );
and \U$21420 ( \21763 , \21762 , \11702 );
not \U$21421 ( \21764 , \21762 );
and \U$21422 ( \21765 , \21764 , \10965 );
nor \U$21423 ( \21766 , \21763 , \21765 );
or \U$21424 ( \21767 , \21759 , \21766 );
not \U$21425 ( \21768 , \21766 );
not \U$21426 ( \21769 , \21759 );
or \U$21427 ( \21770 , \21768 , \21769 );
and \U$21428 ( \21771 , \10424 , RI986eda0_37);
and \U$21429 ( \21772 , RI986ebc0_33, \10422 );
nor \U$21430 ( \21773 , \21771 , \21772 );
and \U$21431 ( \21774 , \21773 , \9840 );
not \U$21432 ( \21775 , \21773 );
and \U$21433 ( \21776 , \21775 , \10428 );
nor \U$21434 ( \21777 , \21774 , \21776 );
nand \U$21435 ( \21778 , \21770 , \21777 );
nand \U$21436 ( \21779 , \21767 , \21778 );
and \U$21437 ( \21780 , \21752 , \21779 );
and \U$21438 ( \21781 , \21732 , \21751 );
or \U$21439 ( \21782 , \21780 , \21781 );
xor \U$21440 ( \21783 , \21705 , \21782 );
and \U$21441 ( \21784 , \8486 , RI98715f0_123);
and \U$21442 ( \21785 , RI986ead0_31, \8484 );
nor \U$21443 ( \21786 , \21784 , \21785 );
and \U$21444 ( \21787 , \21786 , \8051 );
not \U$21445 ( \21788 , \21786 );
and \U$21446 ( \21789 , \21788 , \8050 );
nor \U$21447 ( \21790 , \21787 , \21789 );
and \U$21448 ( \21791 , \9237 , RI986e9e0_29);
and \U$21449 ( \21792 , RI986e8f0_27, \9235 );
nor \U$21450 ( \21793 , \21791 , \21792 );
and \U$21451 ( \21794 , \21793 , \8836 );
not \U$21452 ( \21795 , \21793 );
and \U$21453 ( \21796 , \21795 , \9241 );
nor \U$21454 ( \21797 , \21794 , \21796 );
xor \U$21455 ( \21798 , \21790 , \21797 );
and \U$21456 ( \21799 , \7729 , RI98717d0_127);
and \U$21457 ( \21800 , RI9871500_121, \7727 );
nor \U$21458 ( \21801 , \21799 , \21800 );
and \U$21459 ( \21802 , \21801 , \7733 );
not \U$21460 ( \21803 , \21801 );
and \U$21461 ( \21804 , \21803 , \7480 );
nor \U$21462 ( \21805 , \21802 , \21804 );
and \U$21463 ( \21806 , \21798 , \21805 );
and \U$21464 ( \21807 , \21790 , \21797 );
nor \U$21465 ( \21808 , \21806 , \21807 );
and \U$21466 ( \21809 , \6453 , RI9871140_113);
and \U$21467 ( \21810 , RI9871320_117, \6451 );
nor \U$21468 ( \21811 , \21809 , \21810 );
and \U$21469 ( \21812 , \21811 , \6180 );
not \U$21470 ( \21813 , \21811 );
and \U$21471 ( \21814 , \21813 , \6190 );
nor \U$21472 ( \21815 , \21812 , \21814 );
and \U$21473 ( \21816 , \7079 , RI9871410_119);
and \U$21474 ( \21817 , RI98716e0_125, \7077 );
nor \U$21475 ( \21818 , \21816 , \21817 );
and \U$21476 ( \21819 , \21818 , \6709 );
not \U$21477 ( \21820 , \21818 );
and \U$21478 ( \21821 , \21820 , \6710 );
nor \U$21479 ( \21822 , \21819 , \21821 );
xor \U$21480 ( \21823 , \21815 , \21822 );
and \U$21481 ( \21824 , \5881 , RI9870c90_103);
and \U$21482 ( \21825 , RI9871230_115, \5879 );
nor \U$21483 ( \21826 , \21824 , \21825 );
and \U$21484 ( \21827 , \21826 , \5885 );
not \U$21485 ( \21828 , \21826 );
and \U$21486 ( \21829 , \21828 , \5594 );
nor \U$21487 ( \21830 , \21827 , \21829 );
and \U$21488 ( \21831 , \21823 , \21830 );
and \U$21489 ( \21832 , \21815 , \21822 );
nor \U$21490 ( \21833 , \21831 , \21832 );
xor \U$21491 ( \21834 , \21808 , \21833 );
and \U$21492 ( \21835 , \4203 , RI9870ab0_99);
and \U$21493 ( \21836 , RI9870d80_105, \4201 );
nor \U$21494 ( \21837 , \21835 , \21836 );
and \U$21495 ( \21838 , \21837 , \4207 );
not \U$21496 ( \21839 , \21837 );
and \U$21497 ( \21840 , \21839 , \3923 );
nor \U$21498 ( \21841 , \21838 , \21840 );
not \U$21499 ( \21842 , \4521 );
and \U$21500 ( \21843 , \4710 , RI98709c0_97);
and \U$21501 ( \21844 , RI9870e70_107, \4708 );
nor \U$21502 ( \21845 , \21843 , \21844 );
not \U$21503 ( \21846 , \21845 );
or \U$21504 ( \21847 , \21842 , \21846 );
or \U$21505 ( \21848 , \21845 , \4519 );
nand \U$21506 ( \21849 , \21847 , \21848 );
xor \U$21507 ( \21850 , \21841 , \21849 );
and \U$21508 ( \21851 , \5318 , RI9870ba0_101);
and \U$21509 ( \21852 , RI9871050_111, \5316 );
nor \U$21510 ( \21853 , \21851 , \21852 );
and \U$21511 ( \21854 , \21853 , \5052 );
not \U$21512 ( \21855 , \21853 );
and \U$21513 ( \21856 , \21855 , \5322 );
nor \U$21514 ( \21857 , \21854 , \21856 );
and \U$21515 ( \21858 , \21850 , \21857 );
and \U$21516 ( \21859 , \21841 , \21849 );
or \U$21517 ( \21860 , \21858 , \21859 );
and \U$21518 ( \21861 , \21834 , \21860 );
and \U$21519 ( \21862 , \21808 , \21833 );
or \U$21520 ( \21863 , \21861 , \21862 );
and \U$21521 ( \21864 , \21783 , \21863 );
and \U$21522 ( \21865 , \21705 , \21782 );
or \U$21523 ( \21866 , \21864 , \21865 );
xor \U$21524 ( \21867 , \21624 , \21866 );
xor \U$21525 ( \21868 , \20929 , \443 );
xor \U$21526 ( \21869 , \21868 , \20937 );
xor \U$21527 ( \21870 , \21256 , \21258 );
xor \U$21528 ( \21871 , \21870 , \21261 );
and \U$21529 ( \21872 , \21869 , \21871 );
xor \U$21530 ( \21873 , \20903 , \20910 );
xor \U$21531 ( \21874 , \21873 , \20918 );
xor \U$21532 ( \21875 , \21282 , \21287 );
xor \U$21533 ( \21876 , \21874 , \21875 );
xor \U$21534 ( \21877 , \21256 , \21258 );
xor \U$21535 ( \21878 , \21877 , \21261 );
and \U$21536 ( \21879 , \21876 , \21878 );
and \U$21537 ( \21880 , \21869 , \21876 );
or \U$21538 ( \21881 , \21872 , \21879 , \21880 );
and \U$21539 ( \21882 , \21867 , \21881 );
and \U$21540 ( \21883 , \21624 , \21866 );
or \U$21541 ( \21884 , \21882 , \21883 );
xor \U$21542 ( \21885 , \21375 , \21447 );
xor \U$21543 ( \21886 , \21885 , \21529 );
xor \U$21544 ( \21887 , \21264 , \21279 );
xor \U$21545 ( \21888 , \21887 , \21292 );
and \U$21546 ( \21889 , \21886 , \21888 );
xor \U$21547 ( \21890 , \21884 , \21889 );
xor \U$21548 ( \21891 , \21401 , \21417 );
xor \U$21549 ( \21892 , \21891 , \21444 );
xor \U$21550 ( \21893 , \21473 , \21498 );
xor \U$21551 ( \21894 , \21893 , \21526 );
and \U$21552 ( \21895 , \21892 , \21894 );
xor \U$21553 ( \21896 , \20977 , \20984 );
xor \U$21554 ( \21897 , \21896 , \20993 );
xor \U$21555 ( \21898 , \21269 , \21274 );
xor \U$21556 ( \21899 , \21897 , \21898 );
xor \U$21557 ( \21900 , \21473 , \21498 );
xor \U$21558 ( \21901 , \21900 , \21526 );
and \U$21559 ( \21902 , \21899 , \21901 );
and \U$21560 ( \21903 , \21892 , \21899 );
or \U$21561 ( \21904 , \21895 , \21902 , \21903 );
xor \U$21562 ( \21905 , \21555 , \21557 );
xor \U$21563 ( \21906 , \21905 , \21560 );
and \U$21564 ( \21907 , \21904 , \21906 );
xor \U$21565 ( \21908 , \21059 , \21061 );
xor \U$21566 ( \21909 , \21908 , \21064 );
xor \U$21567 ( \21910 , \21537 , \21544 );
xor \U$21568 ( \21911 , \21909 , \21910 );
xor \U$21569 ( \21912 , \21555 , \21557 );
xor \U$21570 ( \21913 , \21912 , \21560 );
and \U$21571 ( \21914 , \21911 , \21913 );
and \U$21572 ( \21915 , \21904 , \21911 );
or \U$21573 ( \21916 , \21907 , \21914 , \21915 );
and \U$21574 ( \21917 , \21890 , \21916 );
and \U$21575 ( \21918 , \21884 , \21889 );
or \U$21576 ( \21919 , \21917 , \21918 );
xor \U$21577 ( \21920 , \20816 , \21056 );
xor \U$21578 ( \21921 , \21920 , \21095 );
xor \U$21579 ( \21922 , \21919 , \21921 );
xor \U$21580 ( \21923 , \21295 , \21532 );
xor \U$21581 ( \21924 , \21923 , \21549 );
xor \U$21582 ( \21925 , \21244 , \21248 );
xor \U$21583 ( \21926 , \21925 , \21251 );
and \U$21584 ( \21927 , \21924 , \21926 );
xor \U$21585 ( \21928 , \21563 , \21564 );
xor \U$21586 ( \21929 , \21928 , \21567 );
xor \U$21587 ( \21930 , \21244 , \21248 );
xor \U$21588 ( \21931 , \21930 , \21251 );
and \U$21589 ( \21932 , \21929 , \21931 );
and \U$21590 ( \21933 , \21924 , \21929 );
or \U$21591 ( \21934 , \21927 , \21932 , \21933 );
and \U$21592 ( \21935 , \21922 , \21934 );
and \U$21593 ( \21936 , \21919 , \21921 );
or \U$21594 ( \21937 , \21935 , \21936 );
and \U$21595 ( \21938 , \21587 , \21937 );
not \U$21596 ( \21939 , \21586 );
and \U$21597 ( \21940 , \21579 , \21939 );
nor \U$21598 ( \21941 , \21938 , \21940 );
not \U$21599 ( \21942 , \21941 );
and \U$21600 ( \21943 , \21577 , \21942 );
and \U$21601 ( \21944 , \21576 , \21941 );
nor \U$21602 ( \21945 , \21943 , \21944 );
not \U$21603 ( \21946 , \21573 );
not \U$21604 ( \21947 , \21238 );
or \U$21605 ( \21948 , \21946 , \21947 );
or \U$21606 ( \21949 , \21238 , \21573 );
nand \U$21607 ( \21950 , \21948 , \21949 );
not \U$21608 ( \21951 , \21950 );
not \U$21609 ( \21952 , \21224 );
and \U$21610 ( \21953 , \21951 , \21952 );
and \U$21611 ( \21954 , \21950 , \21224 );
nor \U$21612 ( \21955 , \21953 , \21954 );
not \U$21613 ( \21956 , \21955 );
not \U$21614 ( \21957 , \21579 );
not \U$21615 ( \21958 , \21937 );
not \U$21616 ( \21959 , \21586 );
and \U$21617 ( \21960 , \21958 , \21959 );
and \U$21618 ( \21961 , \21937 , \21586 );
nor \U$21619 ( \21962 , \21960 , \21961 );
not \U$21620 ( \21963 , \21962 );
or \U$21621 ( \21964 , \21957 , \21963 );
or \U$21622 ( \21965 , \21962 , \21579 );
nand \U$21623 ( \21966 , \21964 , \21965 );
nand \U$21624 ( \21967 , \21956 , \21966 );
or \U$21625 ( \21968 , \21945 , \21967 );
xnor \U$21626 ( \21969 , \21967 , \21945 );
not \U$21627 ( \21970 , \21955 );
not \U$21628 ( \21971 , \21966 );
or \U$21629 ( \21972 , \21970 , \21971 );
or \U$21630 ( \21973 , \21966 , \21955 );
nand \U$21631 ( \21974 , \21972 , \21973 );
not \U$21632 ( \21975 , \21585 );
not \U$21633 ( \21976 , \21582 );
or \U$21634 ( \21977 , \21975 , \21976 );
or \U$21635 ( \21978 , \21582 , \21585 );
nand \U$21636 ( \21979 , \21977 , \21978 );
not \U$21637 ( \21980 , \21979 );
xor \U$21638 ( \21981 , \21919 , \21921 );
xor \U$21639 ( \21982 , \21981 , \21934 );
not \U$21640 ( \21983 , \21982 );
or \U$21641 ( \21984 , \21980 , \21983 );
or \U$21642 ( \21985 , \21982 , \21979 );
xor \U$21643 ( \21986 , \21705 , \21782 );
xor \U$21644 ( \21987 , \21986 , \21863 );
xor \U$21645 ( \21988 , \21597 , \21608 );
xor \U$21646 ( \21989 , \21988 , \21621 );
and \U$21647 ( \21990 , \21987 , \21989 );
xor \U$21648 ( \21991 , \21256 , \21258 );
xor \U$21649 ( \21992 , \21991 , \21261 );
xor \U$21650 ( \21993 , \21869 , \21876 );
xor \U$21651 ( \21994 , \21992 , \21993 );
xor \U$21652 ( \21995 , \21597 , \21608 );
xor \U$21653 ( \21996 , \21995 , \21621 );
and \U$21654 ( \21997 , \21994 , \21996 );
and \U$21655 ( \21998 , \21987 , \21994 );
or \U$21656 ( \21999 , \21990 , \21997 , \21998 );
xor \U$21657 ( \22000 , \21790 , \21797 );
xor \U$21658 ( \22001 , \22000 , \21805 );
not \U$21659 ( \22002 , \22001 );
not \U$21660 ( \22003 , \21766 );
not \U$21661 ( \22004 , \21777 );
or \U$21662 ( \22005 , \22003 , \22004 );
or \U$21663 ( \22006 , \21766 , \21777 );
nand \U$21664 ( \22007 , \22005 , \22006 );
not \U$21665 ( \22008 , \22007 );
not \U$21666 ( \22009 , \21759 );
and \U$21667 ( \22010 , \22008 , \22009 );
and \U$21668 ( \22011 , \22007 , \21759 );
nor \U$21669 ( \22012 , \22010 , \22011 );
not \U$21670 ( \22013 , \22012 );
and \U$21671 ( \22014 , \22002 , \22013 );
and \U$21672 ( \22015 , \22012 , \22001 );
xor \U$21673 ( \22016 , \21815 , \21822 );
xor \U$21674 ( \22017 , \22016 , \21830 );
nor \U$21675 ( \22018 , \22015 , \22017 );
nor \U$21676 ( \22019 , \22014 , \22018 );
not \U$21677 ( \22020 , \21719 );
not \U$21678 ( \22021 , \21730 );
or \U$21679 ( \22022 , \22020 , \22021 );
or \U$21680 ( \22023 , \21719 , \21730 );
nand \U$21681 ( \22024 , \22022 , \22023 );
not \U$21682 ( \22025 , \22024 );
not \U$21683 ( \22026 , \21712 );
and \U$21684 ( \22027 , \22025 , \22026 );
and \U$21685 ( \22028 , \22024 , \21712 );
nor \U$21686 ( \22029 , \22027 , \22028 );
not \U$21687 ( \22030 , \22029 );
xor \U$21688 ( \22031 , \21740 , \451 );
xor \U$21689 ( \22032 , \22031 , \21748 );
nand \U$21690 ( \22033 , \22030 , \22032 );
or \U$21691 ( \22034 , \22019 , \22033 );
not \U$21692 ( \22035 , \22033 );
not \U$21693 ( \22036 , \22019 );
or \U$21694 ( \22037 , \22035 , \22036 );
xor \U$21695 ( \22038 , \21683 , \21691 );
xor \U$21696 ( \22039 , \22038 , \21699 );
xor \U$21697 ( \22040 , \21631 , \21639 );
xor \U$21698 ( \22041 , \22040 , \21648 );
and \U$21699 ( \22042 , \22039 , \22041 );
xor \U$21700 ( \22043 , \21841 , \21849 );
xor \U$21701 ( \22044 , \22043 , \21857 );
xor \U$21702 ( \22045 , \21631 , \21639 );
xor \U$21703 ( \22046 , \22045 , \21648 );
and \U$21704 ( \22047 , \22044 , \22046 );
and \U$21705 ( \22048 , \22039 , \22044 );
or \U$21706 ( \22049 , \22042 , \22047 , \22048 );
nand \U$21707 ( \22050 , \22037 , \22049 );
nand \U$21708 ( \22051 , \22034 , \22050 );
and \U$21709 ( \22052 , \7079 , RI9871320_117);
and \U$21710 ( \22053 , RI9871410_119, \7077 );
nor \U$21711 ( \22054 , \22052 , \22053 );
and \U$21712 ( \22055 , \22054 , \6710 );
not \U$21713 ( \22056 , \22054 );
and \U$21714 ( \22057 , \22056 , \6709 );
nor \U$21715 ( \22058 , \22055 , \22057 );
and \U$21716 ( \22059 , \7729 , RI98716e0_125);
and \U$21717 ( \22060 , RI98717d0_127, \7727 );
nor \U$21718 ( \22061 , \22059 , \22060 );
and \U$21719 ( \22062 , \22061 , \7480 );
not \U$21720 ( \22063 , \22061 );
and \U$21721 ( \22064 , \22063 , \7733 );
nor \U$21722 ( \22065 , \22062 , \22064 );
xor \U$21723 ( \22066 , \22058 , \22065 );
and \U$21724 ( \22067 , \8486 , RI9871500_121);
and \U$21725 ( \22068 , RI98715f0_123, \8484 );
nor \U$21726 ( \22069 , \22067 , \22068 );
and \U$21727 ( \22070 , \22069 , \8050 );
not \U$21728 ( \22071 , \22069 );
and \U$21729 ( \22072 , \22071 , \8051 );
nor \U$21730 ( \22073 , \22070 , \22072 );
and \U$21731 ( \22074 , \22066 , \22073 );
and \U$21732 ( \22075 , \22058 , \22065 );
or \U$21733 ( \22076 , \22074 , \22075 );
not \U$21734 ( \22077 , \3918 );
and \U$21735 ( \22078 , \3683 , RI9870060_77);
and \U$21736 ( \22079 , RI9870150_79, \3681 );
nor \U$21737 ( \22080 , \22078 , \22079 );
not \U$21738 ( \22081 , \22080 );
or \U$21739 ( \22082 , \22077 , \22081 );
or \U$21740 ( \22083 , \22080 , \3918 );
nand \U$21741 ( \22084 , \22082 , \22083 );
and \U$21742 ( \22085 , \4203 , RI9870f60_109);
and \U$21743 ( \22086 , RI9870ab0_99, \4201 );
nor \U$21744 ( \22087 , \22085 , \22086 );
and \U$21745 ( \22088 , \22087 , \4207 );
not \U$21746 ( \22089 , \22087 );
and \U$21747 ( \22090 , \22089 , \3923 );
nor \U$21748 ( \22091 , \22088 , \22090 );
xor \U$21749 ( \22092 , \22084 , \22091 );
not \U$21750 ( \22093 , \4519 );
and \U$21751 ( \22094 , \4710 , RI9870d80_105);
and \U$21752 ( \22095 , RI98709c0_97, \4708 );
nor \U$21753 ( \22096 , \22094 , \22095 );
not \U$21754 ( \22097 , \22096 );
or \U$21755 ( \22098 , \22093 , \22097 );
or \U$21756 ( \22099 , \22096 , \4519 );
nand \U$21757 ( \22100 , \22098 , \22099 );
and \U$21758 ( \22101 , \22092 , \22100 );
and \U$21759 ( \22102 , \22084 , \22091 );
or \U$21760 ( \22103 , \22101 , \22102 );
xor \U$21761 ( \22104 , \22076 , \22103 );
and \U$21762 ( \22105 , \5881 , RI9871050_111);
and \U$21763 ( \22106 , RI9870c90_103, \5879 );
nor \U$21764 ( \22107 , \22105 , \22106 );
and \U$21765 ( \22108 , \22107 , \5594 );
not \U$21766 ( \22109 , \22107 );
and \U$21767 ( \22110 , \22109 , \5885 );
nor \U$21768 ( \22111 , \22108 , \22110 );
and \U$21769 ( \22112 , \5318 , RI9870e70_107);
and \U$21770 ( \22113 , RI9870ba0_101, \5316 );
nor \U$21771 ( \22114 , \22112 , \22113 );
and \U$21772 ( \22115 , \22114 , \5052 );
not \U$21773 ( \22116 , \22114 );
and \U$21774 ( \22117 , \22116 , \5322 );
nor \U$21775 ( \22118 , \22115 , \22117 );
xor \U$21776 ( \22119 , \22111 , \22118 );
and \U$21777 ( \22120 , \6453 , RI9871230_115);
and \U$21778 ( \22121 , RI9871140_113, \6451 );
nor \U$21779 ( \22122 , \22120 , \22121 );
and \U$21780 ( \22123 , \22122 , \6190 );
not \U$21781 ( \22124 , \22122 );
and \U$21782 ( \22125 , \22124 , \6705 );
nor \U$21783 ( \22126 , \22123 , \22125 );
and \U$21784 ( \22127 , \22119 , \22126 );
and \U$21785 ( \22128 , \22111 , \22118 );
or \U$21786 ( \22129 , \22127 , \22128 );
and \U$21787 ( \22130 , \22104 , \22129 );
and \U$21788 ( \22131 , \22076 , \22103 );
or \U$21789 ( \22132 , \22130 , \22131 );
and \U$21790 ( \22133 , \9237 , RI986ead0_31);
and \U$21791 ( \22134 , RI986e9e0_29, \9235 );
nor \U$21792 ( \22135 , \22133 , \22134 );
and \U$21793 ( \22136 , \22135 , \9241 );
not \U$21794 ( \22137 , \22135 );
and \U$21795 ( \22138 , \22137 , \8836 );
nor \U$21796 ( \22139 , \22136 , \22138 );
and \U$21797 ( \22140 , \9505 , RI986e8f0_27);
and \U$21798 ( \22141 , RI986e800_25, \9503 );
nor \U$21799 ( \22142 , \22140 , \22141 );
and \U$21800 ( \22143 , \22142 , \9510 );
not \U$21801 ( \22144 , \22142 );
and \U$21802 ( \22145 , \22144 , \9513 );
nor \U$21803 ( \22146 , \22143 , \22145 );
xor \U$21804 ( \22147 , \22139 , \22146 );
and \U$21805 ( \22148 , \10424 , RI986ee90_39);
and \U$21806 ( \22149 , RI986eda0_37, \10422 );
nor \U$21807 ( \22150 , \22148 , \22149 );
and \U$21808 ( \22151 , \22150 , \9840 );
not \U$21809 ( \22152 , \22150 );
and \U$21810 ( \22153 , \22152 , \10428 );
nor \U$21811 ( \22154 , \22151 , \22153 );
and \U$21812 ( \22155 , \22147 , \22154 );
and \U$21813 ( \22156 , \22139 , \22146 );
or \U$21814 ( \22157 , \22155 , \22156 );
and \U$21815 ( \22158 , \14937 , RI986e710_23);
and \U$21816 ( \22159 , RI986e620_21, \14935 );
nor \U$21817 ( \22160 , \22158 , \22159 );
and \U$21818 ( \22161 , \22160 , \14539 );
not \U$21819 ( \22162 , \22160 );
and \U$21820 ( \22163 , \22162 , \14538 );
nor \U$21821 ( \22164 , \22161 , \22163 );
not \U$21822 ( \22165 , RI9873558_190);
and \U$21823 ( \22166 , \15780 , RI986f7f0_59);
and \U$21824 ( \22167 , RI9873648_192, RI986f700_57);
nor \U$21825 ( \22168 , \22166 , \22167 );
not \U$21826 ( \22169 , \22168 );
or \U$21827 ( \22170 , \22165 , \22169 );
or \U$21828 ( \22171 , \22168 , RI9873558_190);
nand \U$21829 ( \22172 , \22170 , \22171 );
xor \U$21830 ( \22173 , \22164 , \22172 );
and \U$21831 ( \22174 , \13882 , RI986e530_19);
and \U$21832 ( \22175 , RI986e440_17, \13880 );
nor \U$21833 ( \22176 , \22174 , \22175 );
and \U$21834 ( \22177 , \22176 , \13358 );
not \U$21835 ( \22178 , \22176 );
and \U$21836 ( \22179 , \22178 , \13359 );
nor \U$21837 ( \22180 , \22177 , \22179 );
and \U$21838 ( \22181 , \22173 , \22180 );
and \U$21839 ( \22182 , \22164 , \22172 );
or \U$21840 ( \22183 , \22181 , \22182 );
xor \U$21841 ( \22184 , \22157 , \22183 );
and \U$21842 ( \22185 , \11696 , RI986ebc0_33);
and \U$21843 ( \22186 , RI986ecb0_35, \11694 );
nor \U$21844 ( \22187 , \22185 , \22186 );
and \U$21845 ( \22188 , \22187 , \10965 );
not \U$21846 ( \22189 , \22187 );
and \U$21847 ( \22190 , \22189 , \11702 );
nor \U$21848 ( \22191 , \22188 , \22190 );
and \U$21849 ( \22192 , \12293 , RI986f070_43);
and \U$21850 ( \22193 , RI986ef80_41, \12291 );
nor \U$21851 ( \22194 , \22192 , \22193 );
and \U$21852 ( \22195 , \22194 , \11687 );
not \U$21853 ( \22196 , \22194 );
and \U$21854 ( \22197 , \22196 , \11686 );
nor \U$21855 ( \22198 , \22195 , \22197 );
xor \U$21856 ( \22199 , \22191 , \22198 );
and \U$21857 ( \22200 , \13045 , RI986f250_47);
and \U$21858 ( \22201 , RI986f160_45, \13043 );
nor \U$21859 ( \22202 , \22200 , \22201 );
and \U$21860 ( \22203 , \22202 , \13047 );
not \U$21861 ( \22204 , \22202 );
and \U$21862 ( \22205 , \22204 , \12619 );
nor \U$21863 ( \22206 , \22203 , \22205 );
and \U$21864 ( \22207 , \22199 , \22206 );
and \U$21865 ( \22208 , \22191 , \22198 );
or \U$21866 ( \22209 , \22207 , \22208 );
and \U$21867 ( \22210 , \22184 , \22209 );
and \U$21868 ( \22211 , \22157 , \22183 );
or \U$21869 ( \22212 , \22210 , \22211 );
xor \U$21870 ( \22213 , \22132 , \22212 );
and \U$21871 ( \22214 , \1329 , RI9870330_83);
and \U$21872 ( \22215 , RI9870240_81, \1327 );
nor \U$21873 ( \22216 , \22214 , \22215 );
and \U$21874 ( \22217 , \22216 , \1336 );
not \U$21875 ( \22218 , \22216 );
and \U$21876 ( \22219 , \22218 , \1337 );
nor \U$21877 ( \22220 , \22217 , \22219 );
and \U$21878 ( \22221 , \1311 , RI98706f0_91);
and \U$21879 ( \22222 , RI9870600_89, \1309 );
nor \U$21880 ( \22223 , \22221 , \22222 );
and \U$21881 ( \22224 , \22223 , \1458 );
not \U$21882 ( \22225 , \22223 );
and \U$21883 ( \22226 , \22225 , \1318 );
nor \U$21884 ( \22227 , \22224 , \22226 );
xor \U$21885 ( \22228 , \22220 , \22227 );
not \U$21886 ( \22229 , \1462 );
and \U$21887 ( \22230 , \2042 , RI98708d0_95);
and \U$21888 ( \22231 , RI98707e0_93, \2040 );
nor \U$21889 ( \22232 , \22230 , \22231 );
not \U$21890 ( \22233 , \22232 );
or \U$21891 ( \22234 , \22229 , \22233 );
or \U$21892 ( \22235 , \22232 , \1462 );
nand \U$21893 ( \22236 , \22234 , \22235 );
and \U$21894 ( \22237 , \22228 , \22236 );
and \U$21895 ( \22238 , \22220 , \22227 );
or \U$21896 ( \22239 , \22237 , \22238 );
and \U$21897 ( \22240 , \2274 , RI986fac0_65);
and \U$21898 ( \22241 , RI986fbb0_67, \2272 );
nor \U$21899 ( \22242 , \22240 , \22241 );
and \U$21900 ( \22243 , \22242 , \2030 );
not \U$21901 ( \22244 , \22242 );
and \U$21902 ( \22245 , \22244 , \2031 );
nor \U$21903 ( \22246 , \22243 , \22245 );
and \U$21904 ( \22247 , \2464 , RI986fd90_71);
and \U$21905 ( \22248 , RI986fca0_69, \2462 );
nor \U$21906 ( \22249 , \22247 , \22248 );
and \U$21907 ( \22250 , \22249 , \2468 );
not \U$21908 ( \22251 , \22249 );
and \U$21909 ( \22252 , \22251 , \2263 );
nor \U$21910 ( \22253 , \22250 , \22252 );
xor \U$21911 ( \22254 , \22246 , \22253 );
not \U$21912 ( \22255 , \3406 );
and \U$21913 ( \22256 , \3254 , RI986ff70_75);
and \U$21914 ( \22257 , RI986fe80_73, \3252 );
nor \U$21915 ( \22258 , \22256 , \22257 );
not \U$21916 ( \22259 , \22258 );
or \U$21917 ( \22260 , \22255 , \22259 );
or \U$21918 ( \22261 , \22258 , \3406 );
nand \U$21919 ( \22262 , \22260 , \22261 );
and \U$21920 ( \22263 , \22254 , \22262 );
and \U$21921 ( \22264 , \22246 , \22253 );
or \U$21922 ( \22265 , \22263 , \22264 );
xor \U$21923 ( \22266 , \22239 , \22265 );
xor \U$21924 ( \22267 , \21658 , \21663 );
xor \U$21925 ( \22268 , \22267 , \21672 );
and \U$21926 ( \22269 , \22266 , \22268 );
and \U$21927 ( \22270 , \22239 , \22265 );
or \U$21928 ( \22271 , \22269 , \22270 );
and \U$21929 ( \22272 , \22213 , \22271 );
and \U$21930 ( \22273 , \22132 , \22212 );
or \U$21931 ( \22274 , \22272 , \22273 );
xor \U$21932 ( \22275 , \22051 , \22274 );
xor \U$21933 ( \22276 , \21455 , \21462 );
xor \U$21934 ( \22277 , \22276 , \21470 );
xor \U$21935 ( \22278 , \21611 , \21616 );
xor \U$21936 ( \22279 , \22277 , \22278 );
xor \U$21937 ( \22280 , \21589 , \21591 );
xor \U$21938 ( \22281 , \22280 , \21594 );
and \U$21939 ( \22282 , \22279 , \22281 );
xor \U$21940 ( \22283 , \21425 , \21432 );
xor \U$21941 ( \22284 , \22283 , \21441 );
xor \U$21942 ( \22285 , \21598 , \21603 );
xor \U$21943 ( \22286 , \22284 , \22285 );
xor \U$21944 ( \22287 , \21589 , \21591 );
xor \U$21945 ( \22288 , \22287 , \21594 );
and \U$21946 ( \22289 , \22286 , \22288 );
and \U$21947 ( \22290 , \22279 , \22286 );
or \U$21948 ( \22291 , \22282 , \22289 , \22290 );
and \U$21949 ( \22292 , \22275 , \22291 );
and \U$21950 ( \22293 , \22051 , \22274 );
or \U$21951 ( \22294 , \22292 , \22293 );
xor \U$21952 ( \22295 , \21999 , \22294 );
xor \U$21953 ( \22296 , \21808 , \21833 );
xor \U$21954 ( \22297 , \22296 , \21860 );
xor \U$21955 ( \22298 , \21732 , \21751 );
xor \U$21956 ( \22299 , \22298 , \21779 );
xor \U$21957 ( \22300 , \22297 , \22299 );
xor \U$21958 ( \22301 , \21651 , \21675 );
xor \U$21959 ( \22302 , \22301 , \21702 );
and \U$21960 ( \22303 , \22300 , \22302 );
and \U$21961 ( \22304 , \22297 , \22299 );
or \U$21962 ( \22305 , \22303 , \22304 );
xor \U$21963 ( \22306 , \21320 , \21346 );
xor \U$21964 ( \22307 , \22306 , \21372 );
xor \U$21965 ( \22308 , \22305 , \22307 );
xor \U$21966 ( \22309 , \21473 , \21498 );
xor \U$21967 ( \22310 , \22309 , \21526 );
xor \U$21968 ( \22311 , \21892 , \21899 );
xor \U$21969 ( \22312 , \22310 , \22311 );
and \U$21970 ( \22313 , \22308 , \22312 );
and \U$21971 ( \22314 , \22305 , \22307 );
or \U$21972 ( \22315 , \22313 , \22314 );
and \U$21973 ( \22316 , \22295 , \22315 );
and \U$21974 ( \22317 , \21999 , \22294 );
or \U$21975 ( \22318 , \22316 , \22317 );
xor \U$21976 ( \22319 , \21886 , \21888 );
xor \U$21977 ( \22320 , \21624 , \21866 );
xor \U$21978 ( \22321 , \22320 , \21881 );
and \U$21979 ( \22322 , \22319 , \22321 );
xor \U$21980 ( \22323 , \21555 , \21557 );
xor \U$21981 ( \22324 , \22323 , \21560 );
xor \U$21982 ( \22325 , \21904 , \21911 );
xor \U$21983 ( \22326 , \22324 , \22325 );
xor \U$21984 ( \22327 , \21624 , \21866 );
xor \U$21985 ( \22328 , \22327 , \21881 );
and \U$21986 ( \22329 , \22326 , \22328 );
and \U$21987 ( \22330 , \22319 , \22326 );
or \U$21988 ( \22331 , \22322 , \22329 , \22330 );
xor \U$21989 ( \22332 , \22318 , \22331 );
xor \U$21990 ( \22333 , \21244 , \21248 );
xor \U$21991 ( \22334 , \22333 , \21251 );
xor \U$21992 ( \22335 , \21924 , \21929 );
xor \U$21993 ( \22336 , \22334 , \22335 );
and \U$21994 ( \22337 , \22332 , \22336 );
and \U$21995 ( \22338 , \22318 , \22331 );
or \U$21996 ( \22339 , \22337 , \22338 );
nand \U$21997 ( \22340 , \21985 , \22339 );
nand \U$21998 ( \22341 , \21984 , \22340 );
and \U$21999 ( \22342 , \21974 , \22341 );
xor \U$22000 ( \22343 , \22341 , \21974 );
xnor \U$22001 ( \22344 , \22339 , \21982 );
not \U$22002 ( \22345 , \22344 );
not \U$22003 ( \22346 , \21979 );
and \U$22004 ( \22347 , \22345 , \22346 );
and \U$22005 ( \22348 , \22344 , \21979 );
nor \U$22006 ( \22349 , \22347 , \22348 );
xor \U$22007 ( \22350 , \22318 , \22331 );
xor \U$22008 ( \22351 , \22350 , \22336 );
xor \U$22009 ( \22352 , \21884 , \21889 );
xor \U$22010 ( \22353 , \22352 , \21916 );
xor \U$22011 ( \22354 , \22351 , \22353 );
xor \U$22012 ( \22355 , \22239 , \22265 );
xor \U$22013 ( \22356 , \22355 , \22268 );
xor \U$22014 ( \22357 , \22076 , \22103 );
xor \U$22015 ( \22358 , \22357 , \22129 );
xor \U$22016 ( \22359 , \22356 , \22358 );
xor \U$22017 ( \22360 , \22157 , \22183 );
xor \U$22018 ( \22361 , \22360 , \22209 );
and \U$22019 ( \22362 , \22359 , \22361 );
and \U$22020 ( \22363 , \22356 , \22358 );
or \U$22021 ( \22364 , \22362 , \22363 );
xor \U$22022 ( \22365 , \22297 , \22299 );
xor \U$22023 ( \22366 , \22365 , \22302 );
and \U$22024 ( \22367 , \22364 , \22366 );
xor \U$22025 ( \22368 , \21589 , \21591 );
xor \U$22026 ( \22369 , \22368 , \21594 );
xor \U$22027 ( \22370 , \22279 , \22286 );
xor \U$22028 ( \22371 , \22369 , \22370 );
xor \U$22029 ( \22372 , \22297 , \22299 );
xor \U$22030 ( \22373 , \22372 , \22302 );
and \U$22031 ( \22374 , \22371 , \22373 );
and \U$22032 ( \22375 , \22364 , \22371 );
or \U$22033 ( \22376 , \22367 , \22374 , \22375 );
xor \U$22034 ( \22377 , \22220 , \22227 );
xor \U$22035 ( \22378 , \22377 , \22236 );
xor \U$22036 ( \22379 , \22084 , \22091 );
xor \U$22037 ( \22380 , \22379 , \22100 );
and \U$22038 ( \22381 , \22378 , \22380 );
xor \U$22039 ( \22382 , \22246 , \22253 );
xor \U$22040 ( \22383 , \22382 , \22262 );
xor \U$22041 ( \22384 , \22084 , \22091 );
xor \U$22042 ( \22385 , \22384 , \22100 );
and \U$22043 ( \22386 , \22383 , \22385 );
and \U$22044 ( \22387 , \22378 , \22383 );
or \U$22045 ( \22388 , \22381 , \22386 , \22387 );
xor \U$22046 ( \22389 , \22191 , \22198 );
xor \U$22047 ( \22390 , \22389 , \22206 );
xor \U$22048 ( \22391 , \22164 , \22172 );
xor \U$22049 ( \22392 , \22391 , \22180 );
and \U$22050 ( \22393 , \22390 , \22392 );
xor \U$22051 ( \22394 , \22388 , \22393 );
xor \U$22052 ( \22395 , \22111 , \22118 );
xor \U$22053 ( \22396 , \22395 , \22126 );
xor \U$22054 ( \22397 , \22058 , \22065 );
xor \U$22055 ( \22398 , \22397 , \22073 );
xor \U$22056 ( \22399 , \22396 , \22398 );
xor \U$22057 ( \22400 , \22139 , \22146 );
xor \U$22058 ( \22401 , \22400 , \22154 );
and \U$22059 ( \22402 , \22399 , \22401 );
and \U$22060 ( \22403 , \22396 , \22398 );
or \U$22061 ( \22404 , \22402 , \22403 );
and \U$22062 ( \22405 , \22394 , \22404 );
and \U$22063 ( \22406 , \22388 , \22393 );
or \U$22064 ( \22407 , \22405 , \22406 );
and \U$22065 ( \22408 , \9505 , RI986e9e0_29);
and \U$22066 ( \22409 , RI986e8f0_27, \9503 );
nor \U$22067 ( \22410 , \22408 , \22409 );
and \U$22068 ( \22411 , \22410 , \9510 );
not \U$22069 ( \22412 , \22410 );
and \U$22070 ( \22413 , \22412 , \9513 );
nor \U$22071 ( \22414 , \22411 , \22413 );
and \U$22072 ( \22415 , \10424 , RI986e800_25);
and \U$22073 ( \22416 , RI986ee90_39, \10422 );
nor \U$22074 ( \22417 , \22415 , \22416 );
and \U$22075 ( \22418 , \22417 , \9840 );
not \U$22076 ( \22419 , \22417 );
and \U$22077 ( \22420 , \22419 , \10428 );
nor \U$22078 ( \22421 , \22418 , \22420 );
xor \U$22079 ( \22422 , \22414 , \22421 );
and \U$22080 ( \22423 , \11696 , RI986eda0_37);
and \U$22081 ( \22424 , RI986ebc0_33, \11694 );
nor \U$22082 ( \22425 , \22423 , \22424 );
and \U$22083 ( \22426 , \22425 , \10965 );
not \U$22084 ( \22427 , \22425 );
and \U$22085 ( \22428 , \22427 , \11702 );
nor \U$22086 ( \22429 , \22426 , \22428 );
and \U$22087 ( \22430 , \22422 , \22429 );
and \U$22088 ( \22431 , \22414 , \22421 );
or \U$22089 ( \22432 , \22430 , \22431 );
not \U$22090 ( \22433 , RI9873558_190);
and \U$22091 ( \22434 , \15780 , RI986e620_21);
and \U$22092 ( \22435 , RI9873648_192, RI986f7f0_59);
nor \U$22093 ( \22436 , \22434 , \22435 );
not \U$22094 ( \22437 , \22436 );
or \U$22095 ( \22438 , \22433 , \22437 );
or \U$22096 ( \22439 , \22436 , RI9873558_190);
nand \U$22097 ( \22440 , \22438 , \22439 );
xor \U$22098 ( \22441 , \22440 , \1128 );
and \U$22099 ( \22442 , \14937 , RI986e440_17);
and \U$22100 ( \22443 , RI986e710_23, \14935 );
nor \U$22101 ( \22444 , \22442 , \22443 );
and \U$22102 ( \22445 , \22444 , \14539 );
not \U$22103 ( \22446 , \22444 );
and \U$22104 ( \22447 , \22446 , \14538 );
nor \U$22105 ( \22448 , \22445 , \22447 );
and \U$22106 ( \22449 , \22441 , \22448 );
and \U$22107 ( \22450 , \22440 , \1128 );
or \U$22108 ( \22451 , \22449 , \22450 );
xor \U$22109 ( \22452 , \22432 , \22451 );
and \U$22110 ( \22453 , \12293 , RI986ecb0_35);
and \U$22111 ( \22454 , RI986f070_43, \12291 );
nor \U$22112 ( \22455 , \22453 , \22454 );
and \U$22113 ( \22456 , \22455 , \11687 );
not \U$22114 ( \22457 , \22455 );
and \U$22115 ( \22458 , \22457 , \11686 );
nor \U$22116 ( \22459 , \22456 , \22458 );
and \U$22117 ( \22460 , \13045 , RI986ef80_41);
and \U$22118 ( \22461 , RI986f250_47, \13043 );
nor \U$22119 ( \22462 , \22460 , \22461 );
and \U$22120 ( \22463 , \22462 , \13047 );
not \U$22121 ( \22464 , \22462 );
and \U$22122 ( \22465 , \22464 , \12619 );
nor \U$22123 ( \22466 , \22463 , \22465 );
xor \U$22124 ( \22467 , \22459 , \22466 );
and \U$22125 ( \22468 , \13882 , RI986f160_45);
and \U$22126 ( \22469 , RI986e530_19, \13880 );
nor \U$22127 ( \22470 , \22468 , \22469 );
and \U$22128 ( \22471 , \22470 , \13358 );
not \U$22129 ( \22472 , \22470 );
and \U$22130 ( \22473 , \22472 , \13359 );
nor \U$22131 ( \22474 , \22471 , \22473 );
and \U$22132 ( \22475 , \22467 , \22474 );
and \U$22133 ( \22476 , \22459 , \22466 );
or \U$22134 ( \22477 , \22475 , \22476 );
and \U$22135 ( \22478 , \22452 , \22477 );
and \U$22136 ( \22479 , \22432 , \22451 );
or \U$22137 ( \22480 , \22478 , \22479 );
not \U$22138 ( \22481 , \3412 );
and \U$22139 ( \22482 , \3683 , RI986fe80_73);
and \U$22140 ( \22483 , RI9870060_77, \3681 );
nor \U$22141 ( \22484 , \22482 , \22483 );
not \U$22142 ( \22485 , \22484 );
or \U$22143 ( \22486 , \22481 , \22485 );
or \U$22144 ( \22487 , \22484 , \3918 );
nand \U$22145 ( \22488 , \22486 , \22487 );
and \U$22146 ( \22489 , \2464 , RI986fbb0_67);
and \U$22147 ( \22490 , RI986fd90_71, \2462 );
nor \U$22148 ( \22491 , \22489 , \22490 );
and \U$22149 ( \22492 , \22491 , \2468 );
not \U$22150 ( \22493 , \22491 );
and \U$22151 ( \22494 , \22493 , \2263 );
nor \U$22152 ( \22495 , \22492 , \22494 );
xor \U$22153 ( \22496 , \22488 , \22495 );
not \U$22154 ( \22497 , \2935 );
and \U$22155 ( \22498 , \3254 , RI986fca0_69);
and \U$22156 ( \22499 , RI986ff70_75, \3252 );
nor \U$22157 ( \22500 , \22498 , \22499 );
not \U$22158 ( \22501 , \22500 );
or \U$22159 ( \22502 , \22497 , \22501 );
or \U$22160 ( \22503 , \22500 , \2935 );
nand \U$22161 ( \22504 , \22502 , \22503 );
and \U$22162 ( \22505 , \22496 , \22504 );
and \U$22163 ( \22506 , \22488 , \22495 );
or \U$22164 ( \22507 , \22505 , \22506 );
not \U$22165 ( \22508 , \1301 );
and \U$22166 ( \22509 , \1293 , RI9870420_85);
and \U$22167 ( \22510 , RI9870510_87, \1291 );
nor \U$22168 ( \22511 , \22509 , \22510 );
not \U$22169 ( \22512 , \22511 );
or \U$22170 ( \22513 , \22508 , \22512 );
or \U$22171 ( \22514 , \22511 , \1128 );
nand \U$22172 ( \22515 , \22513 , \22514 );
xor \U$22173 ( \22516 , \22507 , \22515 );
and \U$22174 ( \22517 , \1311 , RI9870240_81);
and \U$22175 ( \22518 , RI98706f0_91, \1309 );
nor \U$22176 ( \22519 , \22517 , \22518 );
and \U$22177 ( \22520 , \22519 , \1458 );
not \U$22178 ( \22521 , \22519 );
and \U$22179 ( \22522 , \22521 , \1318 );
nor \U$22180 ( \22523 , \22520 , \22522 );
not \U$22181 ( \22524 , \2034 );
and \U$22182 ( \22525 , \2042 , RI9870600_89);
and \U$22183 ( \22526 , RI98708d0_95, \2040 );
nor \U$22184 ( \22527 , \22525 , \22526 );
not \U$22185 ( \22528 , \22527 );
or \U$22186 ( \22529 , \22524 , \22528 );
or \U$22187 ( \22530 , \22527 , \1462 );
nand \U$22188 ( \22531 , \22529 , \22530 );
xor \U$22189 ( \22532 , \22523 , \22531 );
and \U$22190 ( \22533 , \2274 , RI98707e0_93);
and \U$22191 ( \22534 , RI986fac0_65, \2272 );
nor \U$22192 ( \22535 , \22533 , \22534 );
and \U$22193 ( \22536 , \22535 , \2030 );
not \U$22194 ( \22537 , \22535 );
and \U$22195 ( \22538 , \22537 , \2031 );
nor \U$22196 ( \22539 , \22536 , \22538 );
and \U$22197 ( \22540 , \22532 , \22539 );
and \U$22198 ( \22541 , \22523 , \22531 );
or \U$22199 ( \22542 , \22540 , \22541 );
and \U$22200 ( \22543 , \22516 , \22542 );
and \U$22201 ( \22544 , \22507 , \22515 );
or \U$22202 ( \22545 , \22543 , \22544 );
xor \U$22203 ( \22546 , \22480 , \22545 );
and \U$22204 ( \22547 , \7729 , RI9871410_119);
and \U$22205 ( \22548 , RI98716e0_125, \7727 );
nor \U$22206 ( \22549 , \22547 , \22548 );
and \U$22207 ( \22550 , \22549 , \7480 );
not \U$22208 ( \22551 , \22549 );
and \U$22209 ( \22552 , \22551 , \7733 );
nor \U$22210 ( \22553 , \22550 , \22552 );
and \U$22211 ( \22554 , \8486 , RI98717d0_127);
and \U$22212 ( \22555 , RI9871500_121, \8484 );
nor \U$22213 ( \22556 , \22554 , \22555 );
and \U$22214 ( \22557 , \22556 , \8050 );
not \U$22215 ( \22558 , \22556 );
and \U$22216 ( \22559 , \22558 , \8051 );
nor \U$22217 ( \22560 , \22557 , \22559 );
xor \U$22218 ( \22561 , \22553 , \22560 );
and \U$22219 ( \22562 , \9237 , RI98715f0_123);
and \U$22220 ( \22563 , RI986ead0_31, \9235 );
nor \U$22221 ( \22564 , \22562 , \22563 );
and \U$22222 ( \22565 , \22564 , \9241 );
not \U$22223 ( \22566 , \22564 );
and \U$22224 ( \22567 , \22566 , \8836 );
nor \U$22225 ( \22568 , \22565 , \22567 );
and \U$22226 ( \22569 , \22561 , \22568 );
and \U$22227 ( \22570 , \22553 , \22560 );
or \U$22228 ( \22571 , \22569 , \22570 );
and \U$22229 ( \22572 , \5881 , RI9870ba0_101);
and \U$22230 ( \22573 , RI9871050_111, \5879 );
nor \U$22231 ( \22574 , \22572 , \22573 );
and \U$22232 ( \22575 , \22574 , \5594 );
not \U$22233 ( \22576 , \22574 );
and \U$22234 ( \22577 , \22576 , \5885 );
nor \U$22235 ( \22578 , \22575 , \22577 );
and \U$22236 ( \22579 , \6453 , RI9870c90_103);
and \U$22237 ( \22580 , RI9871230_115, \6451 );
nor \U$22238 ( \22581 , \22579 , \22580 );
and \U$22239 ( \22582 , \22581 , \6190 );
not \U$22240 ( \22583 , \22581 );
and \U$22241 ( \22584 , \22583 , \6705 );
nor \U$22242 ( \22585 , \22582 , \22584 );
xor \U$22243 ( \22586 , \22578 , \22585 );
and \U$22244 ( \22587 , \7079 , RI9871140_113);
and \U$22245 ( \22588 , RI9871320_117, \7077 );
nor \U$22246 ( \22589 , \22587 , \22588 );
and \U$22247 ( \22590 , \22589 , \6710 );
not \U$22248 ( \22591 , \22589 );
and \U$22249 ( \22592 , \22591 , \6709 );
nor \U$22250 ( \22593 , \22590 , \22592 );
and \U$22251 ( \22594 , \22586 , \22593 );
and \U$22252 ( \22595 , \22578 , \22585 );
or \U$22253 ( \22596 , \22594 , \22595 );
xor \U$22254 ( \22597 , \22571 , \22596 );
not \U$22255 ( \22598 , \4521 );
and \U$22256 ( \22599 , \4710 , RI9870ab0_99);
and \U$22257 ( \22600 , RI9870d80_105, \4708 );
nor \U$22258 ( \22601 , \22599 , \22600 );
not \U$22259 ( \22602 , \22601 );
or \U$22260 ( \22603 , \22598 , \22602 );
or \U$22261 ( \22604 , \22601 , \4519 );
nand \U$22262 ( \22605 , \22603 , \22604 );
and \U$22263 ( \22606 , \4203 , RI9870150_79);
and \U$22264 ( \22607 , RI9870f60_109, \4201 );
nor \U$22265 ( \22608 , \22606 , \22607 );
and \U$22266 ( \22609 , \22608 , \4207 );
not \U$22267 ( \22610 , \22608 );
and \U$22268 ( \22611 , \22610 , \3923 );
nor \U$22269 ( \22612 , \22609 , \22611 );
xor \U$22270 ( \22613 , \22605 , \22612 );
and \U$22271 ( \22614 , \5318 , RI98709c0_97);
and \U$22272 ( \22615 , RI9870e70_107, \5316 );
nor \U$22273 ( \22616 , \22614 , \22615 );
and \U$22274 ( \22617 , \22616 , \5052 );
not \U$22275 ( \22618 , \22616 );
and \U$22276 ( \22619 , \22618 , \5322 );
nor \U$22277 ( \22620 , \22617 , \22619 );
and \U$22278 ( \22621 , \22613 , \22620 );
and \U$22279 ( \22622 , \22605 , \22612 );
or \U$22280 ( \22623 , \22621 , \22622 );
and \U$22281 ( \22624 , \22597 , \22623 );
and \U$22282 ( \22625 , \22571 , \22596 );
or \U$22283 ( \22626 , \22624 , \22625 );
and \U$22284 ( \22627 , \22546 , \22626 );
and \U$22285 ( \22628 , \22480 , \22545 );
or \U$22286 ( \22629 , \22627 , \22628 );
xor \U$22287 ( \22630 , \22407 , \22629 );
not \U$22288 ( \22631 , \22012 );
xor \U$22289 ( \22632 , \22017 , \22001 );
not \U$22290 ( \22633 , \22632 );
or \U$22291 ( \22634 , \22631 , \22633 );
or \U$22292 ( \22635 , \22632 , \22012 );
nand \U$22293 ( \22636 , \22634 , \22635 );
not \U$22294 ( \22637 , \22029 );
not \U$22295 ( \22638 , \22032 );
or \U$22296 ( \22639 , \22637 , \22638 );
or \U$22297 ( \22640 , \22032 , \22029 );
nand \U$22298 ( \22641 , \22639 , \22640 );
xor \U$22299 ( \22642 , \22636 , \22641 );
xor \U$22300 ( \22643 , \21631 , \21639 );
xor \U$22301 ( \22644 , \22643 , \21648 );
xor \U$22302 ( \22645 , \22039 , \22044 );
xor \U$22303 ( \22646 , \22644 , \22645 );
and \U$22304 ( \22647 , \22642 , \22646 );
and \U$22305 ( \22648 , \22636 , \22641 );
or \U$22306 ( \22649 , \22647 , \22648 );
and \U$22307 ( \22650 , \22630 , \22649 );
and \U$22308 ( \22651 , \22407 , \22629 );
or \U$22309 ( \22652 , \22650 , \22651 );
xor \U$22310 ( \22653 , \22376 , \22652 );
xor \U$22311 ( \22654 , \21597 , \21608 );
xor \U$22312 ( \22655 , \22654 , \21621 );
xor \U$22313 ( \22656 , \21987 , \21994 );
xor \U$22314 ( \22657 , \22655 , \22656 );
and \U$22315 ( \22658 , \22653 , \22657 );
and \U$22316 ( \22659 , \22376 , \22652 );
or \U$22317 ( \22660 , \22658 , \22659 );
xor \U$22318 ( \22661 , \21999 , \22294 );
xor \U$22319 ( \22662 , \22661 , \22315 );
and \U$22320 ( \22663 , \22660 , \22662 );
xor \U$22321 ( \22664 , \21624 , \21866 );
xor \U$22322 ( \22665 , \22664 , \21881 );
xor \U$22323 ( \22666 , \22319 , \22326 );
xor \U$22324 ( \22667 , \22665 , \22666 );
xor \U$22325 ( \22668 , \21999 , \22294 );
xor \U$22326 ( \22669 , \22668 , \22315 );
and \U$22327 ( \22670 , \22667 , \22669 );
and \U$22328 ( \22671 , \22660 , \22667 );
or \U$22329 ( \22672 , \22663 , \22670 , \22671 );
and \U$22330 ( \22673 , \22354 , \22672 );
and \U$22331 ( \22674 , \22351 , \22353 );
nor \U$22332 ( \22675 , \22673 , \22674 );
or \U$22333 ( \22676 , \22349 , \22675 );
xnor \U$22334 ( \22677 , \22675 , \22349 );
xor \U$22335 ( \22678 , \22051 , \22274 );
xor \U$22336 ( \22679 , \22678 , \22291 );
xor \U$22337 ( \22680 , \22376 , \22652 );
xor \U$22338 ( \22681 , \22680 , \22657 );
and \U$22339 ( \22682 , \22679 , \22681 );
xor \U$22340 ( \22683 , \22440 , \1128 );
xor \U$22341 ( \22684 , \22683 , \22448 );
xor \U$22342 ( \22685 , \22414 , \22421 );
xor \U$22343 ( \22686 , \22685 , \22429 );
and \U$22344 ( \22687 , \22684 , \22686 );
xor \U$22345 ( \22688 , \22459 , \22466 );
xor \U$22346 ( \22689 , \22688 , \22474 );
xor \U$22347 ( \22690 , \22414 , \22421 );
xor \U$22348 ( \22691 , \22690 , \22429 );
and \U$22349 ( \22692 , \22689 , \22691 );
and \U$22350 ( \22693 , \22684 , \22689 );
or \U$22351 ( \22694 , \22687 , \22692 , \22693 );
xor \U$22352 ( \22695 , \22488 , \22495 );
xor \U$22353 ( \22696 , \22695 , \22504 );
nand \U$22354 ( \22697 , RI9870420_85, \1291 );
not \U$22355 ( \22698 , \22697 );
not \U$22356 ( \22699 , \1301 );
or \U$22357 ( \22700 , \22698 , \22699 );
or \U$22358 ( \22701 , \1128 , \22697 );
nand \U$22359 ( \22702 , \22700 , \22701 );
xor \U$22360 ( \22703 , \22696 , \22702 );
xor \U$22361 ( \22704 , \22523 , \22531 );
xor \U$22362 ( \22705 , \22704 , \22539 );
and \U$22363 ( \22706 , \22703 , \22705 );
and \U$22364 ( \22707 , \22696 , \22702 );
or \U$22365 ( \22708 , \22706 , \22707 );
xor \U$22366 ( \22709 , \22694 , \22708 );
xor \U$22367 ( \22710 , \22605 , \22612 );
xor \U$22368 ( \22711 , \22710 , \22620 );
xor \U$22369 ( \22712 , \22578 , \22585 );
xor \U$22370 ( \22713 , \22712 , \22593 );
and \U$22371 ( \22714 , \22711 , \22713 );
xor \U$22372 ( \22715 , \22553 , \22560 );
xor \U$22373 ( \22716 , \22715 , \22568 );
xor \U$22374 ( \22717 , \22578 , \22585 );
xor \U$22375 ( \22718 , \22717 , \22593 );
and \U$22376 ( \22719 , \22716 , \22718 );
and \U$22377 ( \22720 , \22711 , \22716 );
or \U$22378 ( \22721 , \22714 , \22719 , \22720 );
and \U$22379 ( \22722 , \22709 , \22721 );
and \U$22380 ( \22723 , \22694 , \22708 );
or \U$22381 ( \22724 , \22722 , \22723 );
and \U$22382 ( \22725 , \11696 , RI986ee90_39);
and \U$22383 ( \22726 , RI986eda0_37, \11694 );
nor \U$22384 ( \22727 , \22725 , \22726 );
and \U$22385 ( \22728 , \22727 , \10965 );
not \U$22386 ( \22729 , \22727 );
and \U$22387 ( \22730 , \22729 , \11702 );
nor \U$22388 ( \22731 , \22728 , \22730 );
and \U$22389 ( \22732 , \12293 , RI986ebc0_33);
and \U$22390 ( \22733 , RI986ecb0_35, \12291 );
nor \U$22391 ( \22734 , \22732 , \22733 );
and \U$22392 ( \22735 , \22734 , \11687 );
not \U$22393 ( \22736 , \22734 );
and \U$22394 ( \22737 , \22736 , \11686 );
nor \U$22395 ( \22738 , \22735 , \22737 );
xor \U$22396 ( \22739 , \22731 , \22738 );
and \U$22397 ( \22740 , \13045 , RI986f070_43);
and \U$22398 ( \22741 , RI986ef80_41, \13043 );
nor \U$22399 ( \22742 , \22740 , \22741 );
and \U$22400 ( \22743 , \22742 , \13047 );
not \U$22401 ( \22744 , \22742 );
and \U$22402 ( \22745 , \22744 , \12619 );
nor \U$22403 ( \22746 , \22743 , \22745 );
and \U$22404 ( \22747 , \22739 , \22746 );
and \U$22405 ( \22748 , \22731 , \22738 );
or \U$22406 ( \22749 , \22747 , \22748 );
and \U$22407 ( \22750 , \13882 , RI986f250_47);
and \U$22408 ( \22751 , RI986f160_45, \13880 );
nor \U$22409 ( \22752 , \22750 , \22751 );
and \U$22410 ( \22753 , \22752 , \13358 );
not \U$22411 ( \22754 , \22752 );
and \U$22412 ( \22755 , \22754 , \13359 );
nor \U$22413 ( \22756 , \22753 , \22755 );
not \U$22414 ( \22757 , RI9873558_190);
and \U$22415 ( \22758 , \15780 , RI986e710_23);
and \U$22416 ( \22759 , RI9873648_192, RI986e620_21);
nor \U$22417 ( \22760 , \22758 , \22759 );
not \U$22418 ( \22761 , \22760 );
or \U$22419 ( \22762 , \22757 , \22761 );
or \U$22420 ( \22763 , \22760 , RI9873558_190);
nand \U$22421 ( \22764 , \22762 , \22763 );
xor \U$22422 ( \22765 , \22756 , \22764 );
and \U$22423 ( \22766 , \14937 , RI986e530_19);
and \U$22424 ( \22767 , RI986e440_17, \14935 );
nor \U$22425 ( \22768 , \22766 , \22767 );
and \U$22426 ( \22769 , \22768 , \14539 );
not \U$22427 ( \22770 , \22768 );
and \U$22428 ( \22771 , \22770 , \14538 );
nor \U$22429 ( \22772 , \22769 , \22771 );
and \U$22430 ( \22773 , \22765 , \22772 );
and \U$22431 ( \22774 , \22756 , \22764 );
or \U$22432 ( \22775 , \22773 , \22774 );
xor \U$22433 ( \22776 , \22749 , \22775 );
and \U$22434 ( \22777 , \9237 , RI9871500_121);
and \U$22435 ( \22778 , RI98715f0_123, \9235 );
nor \U$22436 ( \22779 , \22777 , \22778 );
and \U$22437 ( \22780 , \22779 , \9241 );
not \U$22438 ( \22781 , \22779 );
and \U$22439 ( \22782 , \22781 , \8836 );
nor \U$22440 ( \22783 , \22780 , \22782 );
and \U$22441 ( \22784 , \9505 , RI986ead0_31);
and \U$22442 ( \22785 , RI986e9e0_29, \9503 );
nor \U$22443 ( \22786 , \22784 , \22785 );
and \U$22444 ( \22787 , \22786 , \9510 );
not \U$22445 ( \22788 , \22786 );
and \U$22446 ( \22789 , \22788 , \9513 );
nor \U$22447 ( \22790 , \22787 , \22789 );
xor \U$22448 ( \22791 , \22783 , \22790 );
and \U$22449 ( \22792 , \10424 , RI986e8f0_27);
and \U$22450 ( \22793 , RI986e800_25, \10422 );
nor \U$22451 ( \22794 , \22792 , \22793 );
and \U$22452 ( \22795 , \22794 , \9840 );
not \U$22453 ( \22796 , \22794 );
and \U$22454 ( \22797 , \22796 , \10428 );
nor \U$22455 ( \22798 , \22795 , \22797 );
and \U$22456 ( \22799 , \22791 , \22798 );
and \U$22457 ( \22800 , \22783 , \22790 );
or \U$22458 ( \22801 , \22799 , \22800 );
and \U$22459 ( \22802 , \22776 , \22801 );
and \U$22460 ( \22803 , \22749 , \22775 );
or \U$22461 ( \22804 , \22802 , \22803 );
and \U$22462 ( \22805 , \2274 , RI98708d0_95);
and \U$22463 ( \22806 , RI98707e0_93, \2272 );
nor \U$22464 ( \22807 , \22805 , \22806 );
and \U$22465 ( \22808 , \22807 , \2030 );
not \U$22466 ( \22809 , \22807 );
and \U$22467 ( \22810 , \22809 , \2031 );
nor \U$22468 ( \22811 , \22808 , \22810 );
and \U$22469 ( \22812 , \2464 , RI986fac0_65);
and \U$22470 ( \22813 , RI986fbb0_67, \2462 );
nor \U$22471 ( \22814 , \22812 , \22813 );
and \U$22472 ( \22815 , \22814 , \2468 );
not \U$22473 ( \22816 , \22814 );
and \U$22474 ( \22817 , \22816 , \2263 );
nor \U$22475 ( \22818 , \22815 , \22817 );
xor \U$22476 ( \22819 , \22811 , \22818 );
not \U$22477 ( \22820 , \3406 );
and \U$22478 ( \22821 , \3254 , RI986fd90_71);
and \U$22479 ( \22822 , RI986fca0_69, \3252 );
nor \U$22480 ( \22823 , \22821 , \22822 );
not \U$22481 ( \22824 , \22823 );
or \U$22482 ( \22825 , \22820 , \22824 );
or \U$22483 ( \22826 , \22823 , \3406 );
nand \U$22484 ( \22827 , \22825 , \22826 );
and \U$22485 ( \22828 , \22819 , \22827 );
and \U$22486 ( \22829 , \22811 , \22818 );
or \U$22487 ( \22830 , \22828 , \22829 );
and \U$22488 ( \22831 , \1329 , RI9870510_87);
and \U$22489 ( \22832 , RI9870330_83, \1327 );
nor \U$22490 ( \22833 , \22831 , \22832 );
and \U$22491 ( \22834 , \22833 , \1336 );
not \U$22492 ( \22835 , \22833 );
and \U$22493 ( \22836 , \22835 , \1337 );
nor \U$22494 ( \22837 , \22834 , \22836 );
xor \U$22495 ( \22838 , \22830 , \22837 );
and \U$22496 ( \22839 , \1311 , RI9870330_83);
and \U$22497 ( \22840 , RI9870240_81, \1309 );
nor \U$22498 ( \22841 , \22839 , \22840 );
and \U$22499 ( \22842 , \22841 , \1458 );
not \U$22500 ( \22843 , \22841 );
and \U$22501 ( \22844 , \22843 , \1318 );
nor \U$22502 ( \22845 , \22842 , \22844 );
and \U$22503 ( \22846 , \1329 , RI9870420_85);
and \U$22504 ( \22847 , RI9870510_87, \1327 );
nor \U$22505 ( \22848 , \22846 , \22847 );
and \U$22506 ( \22849 , \22848 , \1336 );
not \U$22507 ( \22850 , \22848 );
and \U$22508 ( \22851 , \22850 , \1337 );
nor \U$22509 ( \22852 , \22849 , \22851 );
xor \U$22510 ( \22853 , \22845 , \22852 );
not \U$22511 ( \22854 , \2034 );
and \U$22512 ( \22855 , \2042 , RI98706f0_91);
and \U$22513 ( \22856 , RI9870600_89, \2040 );
nor \U$22514 ( \22857 , \22855 , \22856 );
not \U$22515 ( \22858 , \22857 );
or \U$22516 ( \22859 , \22854 , \22858 );
or \U$22517 ( \22860 , \22857 , \2034 );
nand \U$22518 ( \22861 , \22859 , \22860 );
and \U$22519 ( \22862 , \22853 , \22861 );
and \U$22520 ( \22863 , \22845 , \22852 );
or \U$22521 ( \22864 , \22862 , \22863 );
and \U$22522 ( \22865 , \22838 , \22864 );
and \U$22523 ( \22866 , \22830 , \22837 );
or \U$22524 ( \22867 , \22865 , \22866 );
xor \U$22525 ( \22868 , \22804 , \22867 );
and \U$22526 ( \22869 , \7079 , RI9871230_115);
and \U$22527 ( \22870 , RI9871140_113, \7077 );
nor \U$22528 ( \22871 , \22869 , \22870 );
and \U$22529 ( \22872 , \22871 , \6710 );
not \U$22530 ( \22873 , \22871 );
and \U$22531 ( \22874 , \22873 , \6709 );
nor \U$22532 ( \22875 , \22872 , \22874 );
and \U$22533 ( \22876 , \7729 , RI9871320_117);
and \U$22534 ( \22877 , RI9871410_119, \7727 );
nor \U$22535 ( \22878 , \22876 , \22877 );
and \U$22536 ( \22879 , \22878 , \7480 );
not \U$22537 ( \22880 , \22878 );
and \U$22538 ( \22881 , \22880 , \7733 );
nor \U$22539 ( \22882 , \22879 , \22881 );
xor \U$22540 ( \22883 , \22875 , \22882 );
and \U$22541 ( \22884 , \8486 , RI98716e0_125);
and \U$22542 ( \22885 , RI98717d0_127, \8484 );
nor \U$22543 ( \22886 , \22884 , \22885 );
and \U$22544 ( \22887 , \22886 , \8050 );
not \U$22545 ( \22888 , \22886 );
and \U$22546 ( \22889 , \22888 , \8051 );
nor \U$22547 ( \22890 , \22887 , \22889 );
and \U$22548 ( \22891 , \22883 , \22890 );
and \U$22549 ( \22892 , \22875 , \22882 );
or \U$22550 ( \22893 , \22891 , \22892 );
and \U$22551 ( \22894 , \5318 , RI9870d80_105);
and \U$22552 ( \22895 , RI98709c0_97, \5316 );
nor \U$22553 ( \22896 , \22894 , \22895 );
and \U$22554 ( \22897 , \22896 , \5052 );
not \U$22555 ( \22898 , \22896 );
and \U$22556 ( \22899 , \22898 , \5322 );
nor \U$22557 ( \22900 , \22897 , \22899 );
and \U$22558 ( \22901 , \5881 , RI9870e70_107);
and \U$22559 ( \22902 , RI9870ba0_101, \5879 );
nor \U$22560 ( \22903 , \22901 , \22902 );
and \U$22561 ( \22904 , \22903 , \5594 );
not \U$22562 ( \22905 , \22903 );
and \U$22563 ( \22906 , \22905 , \5885 );
nor \U$22564 ( \22907 , \22904 , \22906 );
xor \U$22565 ( \22908 , \22900 , \22907 );
and \U$22566 ( \22909 , \6453 , RI9871050_111);
and \U$22567 ( \22910 , RI9870c90_103, \6451 );
nor \U$22568 ( \22911 , \22909 , \22910 );
and \U$22569 ( \22912 , \22911 , \6190 );
not \U$22570 ( \22913 , \22911 );
and \U$22571 ( \22914 , \22913 , \6180 );
nor \U$22572 ( \22915 , \22912 , \22914 );
and \U$22573 ( \22916 , \22908 , \22915 );
and \U$22574 ( \22917 , \22900 , \22907 );
or \U$22575 ( \22918 , \22916 , \22917 );
xor \U$22576 ( \22919 , \22893 , \22918 );
not \U$22577 ( \22920 , \3412 );
and \U$22578 ( \22921 , \3683 , RI986ff70_75);
and \U$22579 ( \22922 , RI986fe80_73, \3681 );
nor \U$22580 ( \22923 , \22921 , \22922 );
not \U$22581 ( \22924 , \22923 );
or \U$22582 ( \22925 , \22920 , \22924 );
or \U$22583 ( \22926 , \22923 , \3412 );
nand \U$22584 ( \22927 , \22925 , \22926 );
and \U$22585 ( \22928 , \4203 , RI9870060_77);
and \U$22586 ( \22929 , RI9870150_79, \4201 );
nor \U$22587 ( \22930 , \22928 , \22929 );
and \U$22588 ( \22931 , \22930 , \4207 );
not \U$22589 ( \22932 , \22930 );
and \U$22590 ( \22933 , \22932 , \3923 );
nor \U$22591 ( \22934 , \22931 , \22933 );
xor \U$22592 ( \22935 , \22927 , \22934 );
not \U$22593 ( \22936 , \4519 );
and \U$22594 ( \22937 , \4710 , RI9870f60_109);
and \U$22595 ( \22938 , RI9870ab0_99, \4708 );
nor \U$22596 ( \22939 , \22937 , \22938 );
not \U$22597 ( \22940 , \22939 );
or \U$22598 ( \22941 , \22936 , \22940 );
or \U$22599 ( \22942 , \22939 , \4519 );
nand \U$22600 ( \22943 , \22941 , \22942 );
and \U$22601 ( \22944 , \22935 , \22943 );
and \U$22602 ( \22945 , \22927 , \22934 );
or \U$22603 ( \22946 , \22944 , \22945 );
and \U$22604 ( \22947 , \22919 , \22946 );
and \U$22605 ( \22948 , \22893 , \22918 );
or \U$22606 ( \22949 , \22947 , \22948 );
and \U$22607 ( \22950 , \22868 , \22949 );
and \U$22608 ( \22951 , \22804 , \22867 );
or \U$22609 ( \22952 , \22950 , \22951 );
xor \U$22610 ( \22953 , \22724 , \22952 );
xor \U$22611 ( \22954 , \22390 , \22392 );
xor \U$22612 ( \22955 , \22396 , \22398 );
xor \U$22613 ( \22956 , \22955 , \22401 );
and \U$22614 ( \22957 , \22954 , \22956 );
xor \U$22615 ( \22958 , \22084 , \22091 );
xor \U$22616 ( \22959 , \22958 , \22100 );
xor \U$22617 ( \22960 , \22378 , \22383 );
xor \U$22618 ( \22961 , \22959 , \22960 );
xor \U$22619 ( \22962 , \22396 , \22398 );
xor \U$22620 ( \22963 , \22962 , \22401 );
and \U$22621 ( \22964 , \22961 , \22963 );
and \U$22622 ( \22965 , \22954 , \22961 );
or \U$22623 ( \22966 , \22957 , \22964 , \22965 );
and \U$22624 ( \22967 , \22953 , \22966 );
and \U$22625 ( \22968 , \22724 , \22952 );
nor \U$22626 ( \22969 , \22967 , \22968 );
not \U$22627 ( \22970 , \22049 );
not \U$22628 ( \22971 , \22019 );
or \U$22629 ( \22972 , \22970 , \22971 );
or \U$22630 ( \22973 , \22019 , \22049 );
nand \U$22631 ( \22974 , \22972 , \22973 );
not \U$22632 ( \22975 , \22974 );
not \U$22633 ( \22976 , \22033 );
and \U$22634 ( \22977 , \22975 , \22976 );
and \U$22635 ( \22978 , \22974 , \22033 );
nor \U$22636 ( \22979 , \22977 , \22978 );
or \U$22637 ( \22980 , \22969 , \22979 );
not \U$22638 ( \22981 , \22979 );
not \U$22639 ( \22982 , \22969 );
or \U$22640 ( \22983 , \22981 , \22982 );
xor \U$22641 ( \22984 , \22507 , \22515 );
xor \U$22642 ( \22985 , \22984 , \22542 );
xor \U$22643 ( \22986 , \22432 , \22451 );
xor \U$22644 ( \22987 , \22986 , \22477 );
and \U$22645 ( \22988 , \22985 , \22987 );
xor \U$22646 ( \22989 , \22571 , \22596 );
xor \U$22647 ( \22990 , \22989 , \22623 );
xor \U$22648 ( \22991 , \22432 , \22451 );
xor \U$22649 ( \22992 , \22991 , \22477 );
and \U$22650 ( \22993 , \22990 , \22992 );
and \U$22651 ( \22994 , \22985 , \22990 );
or \U$22652 ( \22995 , \22988 , \22993 , \22994 );
xor \U$22653 ( \22996 , \22356 , \22358 );
xor \U$22654 ( \22997 , \22996 , \22361 );
and \U$22655 ( \22998 , \22995 , \22997 );
xor \U$22656 ( \22999 , \22636 , \22641 );
xor \U$22657 ( \23000 , \22999 , \22646 );
xor \U$22658 ( \23001 , \22356 , \22358 );
xor \U$22659 ( \23002 , \23001 , \22361 );
and \U$22660 ( \23003 , \23000 , \23002 );
and \U$22661 ( \23004 , \22995 , \23000 );
or \U$22662 ( \23005 , \22998 , \23003 , \23004 );
nand \U$22663 ( \23006 , \22983 , \23005 );
nand \U$22664 ( \23007 , \22980 , \23006 );
xor \U$22665 ( \23008 , \22305 , \22307 );
xor \U$22666 ( \23009 , \23008 , \22312 );
xor \U$22667 ( \23010 , \23007 , \23009 );
xor \U$22668 ( \23011 , \22132 , \22212 );
xor \U$22669 ( \23012 , \23011 , \22271 );
xor \U$22670 ( \23013 , \22407 , \22629 );
xor \U$22671 ( \23014 , \23013 , \22649 );
and \U$22672 ( \23015 , \23012 , \23014 );
xor \U$22673 ( \23016 , \22297 , \22299 );
xor \U$22674 ( \23017 , \23016 , \22302 );
xor \U$22675 ( \23018 , \22364 , \22371 );
xor \U$22676 ( \23019 , \23017 , \23018 );
xor \U$22677 ( \23020 , \22407 , \22629 );
xor \U$22678 ( \23021 , \23020 , \22649 );
and \U$22679 ( \23022 , \23019 , \23021 );
and \U$22680 ( \23023 , \23012 , \23019 );
or \U$22681 ( \23024 , \23015 , \23022 , \23023 );
and \U$22682 ( \23025 , \23010 , \23024 );
and \U$22683 ( \23026 , \23007 , \23009 );
or \U$22684 ( \23027 , \23025 , \23026 );
xnor \U$22685 ( \23028 , \22682 , \23027 );
not \U$22686 ( \23029 , \23028 );
xor \U$22687 ( \23030 , \21999 , \22294 );
xor \U$22688 ( \23031 , \23030 , \22315 );
xor \U$22689 ( \23032 , \22660 , \22667 );
xor \U$22690 ( \23033 , \23031 , \23032 );
not \U$22691 ( \23034 , \23033 );
and \U$22692 ( \23035 , \23029 , \23034 );
and \U$22693 ( \23036 , \23028 , \23033 );
nor \U$22694 ( \23037 , \23035 , \23036 );
xor \U$22695 ( \23038 , \22679 , \22681 );
xor \U$22696 ( \23039 , \23007 , \23009 );
xor \U$22697 ( \23040 , \23039 , \23024 );
xor \U$22698 ( \23041 , \23038 , \23040 );
xor \U$22699 ( \23042 , \22724 , \22952 );
xor \U$22700 ( \23043 , \23042 , \22966 );
xor \U$22701 ( \23044 , \22480 , \22545 );
xor \U$22702 ( \23045 , \23044 , \22626 );
xor \U$22703 ( \23046 , \23043 , \23045 );
xor \U$22704 ( \23047 , \22356 , \22358 );
xor \U$22705 ( \23048 , \23047 , \22361 );
xor \U$22706 ( \23049 , \22995 , \23000 );
xor \U$22707 ( \23050 , \23048 , \23049 );
and \U$22708 ( \23051 , \23046 , \23050 );
and \U$22709 ( \23052 , \23043 , \23045 );
or \U$22710 ( \23053 , \23051 , \23052 );
xor \U$22711 ( \23054 , \22927 , \22934 );
xor \U$22712 ( \23055 , \23054 , \22943 );
xor \U$22713 ( \23056 , \22811 , \22818 );
xor \U$22714 ( \23057 , \23056 , \22827 );
and \U$22715 ( \23058 , \23055 , \23057 );
xor \U$22716 ( \23059 , \22900 , \22907 );
xor \U$22717 ( \23060 , \23059 , \22915 );
xor \U$22718 ( \23061 , \22811 , \22818 );
xor \U$22719 ( \23062 , \23061 , \22827 );
and \U$22720 ( \23063 , \23060 , \23062 );
and \U$22721 ( \23064 , \23055 , \23060 );
or \U$22722 ( \23065 , \23058 , \23063 , \23064 );
xor \U$22723 ( \23066 , \22783 , \22790 );
xor \U$22724 ( \23067 , \23066 , \22798 );
xor \U$22725 ( \23068 , \22875 , \22882 );
xor \U$22726 ( \23069 , \23068 , \22890 );
xor \U$22727 ( \23070 , \23067 , \23069 );
xor \U$22728 ( \23071 , \22731 , \22738 );
xor \U$22729 ( \23072 , \23071 , \22746 );
and \U$22730 ( \23073 , \23070 , \23072 );
and \U$22731 ( \23074 , \23067 , \23069 );
or \U$22732 ( \23075 , \23073 , \23074 );
xor \U$22733 ( \23076 , \23065 , \23075 );
xor \U$22734 ( \23077 , \22414 , \22421 );
xor \U$22735 ( \23078 , \23077 , \22429 );
xor \U$22736 ( \23079 , \22684 , \22689 );
xor \U$22737 ( \23080 , \23078 , \23079 );
and \U$22738 ( \23081 , \23076 , \23080 );
and \U$22739 ( \23082 , \23065 , \23075 );
or \U$22740 ( \23083 , \23081 , \23082 );
not \U$22741 ( \23084 , \3406 );
and \U$22742 ( \23085 , \3254 , RI986fbb0_67);
and \U$22743 ( \23086 , RI986fd90_71, \3252 );
nor \U$22744 ( \23087 , \23085 , \23086 );
not \U$22745 ( \23088 , \23087 );
or \U$22746 ( \23089 , \23084 , \23088 );
or \U$22747 ( \23090 , \23087 , \3406 );
nand \U$22748 ( \23091 , \23089 , \23090 );
and \U$22749 ( \23092 , \2464 , RI98707e0_93);
and \U$22750 ( \23093 , RI986fac0_65, \2462 );
nor \U$22751 ( \23094 , \23092 , \23093 );
and \U$22752 ( \23095 , \23094 , \2468 );
not \U$22753 ( \23096 , \23094 );
and \U$22754 ( \23097 , \23096 , \2263 );
nor \U$22755 ( \23098 , \23095 , \23097 );
xor \U$22756 ( \23099 , \23091 , \23098 );
not \U$22757 ( \23100 , \3918 );
and \U$22758 ( \23101 , \3683 , RI986fca0_69);
and \U$22759 ( \23102 , RI986ff70_75, \3681 );
nor \U$22760 ( \23103 , \23101 , \23102 );
not \U$22761 ( \23104 , \23103 );
or \U$22762 ( \23105 , \23100 , \23104 );
or \U$22763 ( \23106 , \23103 , \3918 );
nand \U$22764 ( \23107 , \23105 , \23106 );
and \U$22765 ( \23108 , \23099 , \23107 );
and \U$22766 ( \23109 , \23091 , \23098 );
or \U$22767 ( \23110 , \23108 , \23109 );
and \U$22768 ( \23111 , \1311 , RI9870510_87);
and \U$22769 ( \23112 , RI9870330_83, \1309 );
nor \U$22770 ( \23113 , \23111 , \23112 );
and \U$22771 ( \23114 , \23113 , \1458 );
not \U$22772 ( \23115 , \23113 );
and \U$22773 ( \23116 , \23115 , \1318 );
nor \U$22774 ( \23117 , \23114 , \23116 );
not \U$22775 ( \23118 , \2034 );
and \U$22776 ( \23119 , \2042 , RI9870240_81);
and \U$22777 ( \23120 , RI98706f0_91, \2040 );
nor \U$22778 ( \23121 , \23119 , \23120 );
not \U$22779 ( \23122 , \23121 );
or \U$22780 ( \23123 , \23118 , \23122 );
or \U$22781 ( \23124 , \23121 , \2034 );
nand \U$22782 ( \23125 , \23123 , \23124 );
xor \U$22783 ( \23126 , \23117 , \23125 );
and \U$22784 ( \23127 , \2274 , RI9870600_89);
and \U$22785 ( \23128 , RI98708d0_95, \2272 );
nor \U$22786 ( \23129 , \23127 , \23128 );
and \U$22787 ( \23130 , \23129 , \2030 );
not \U$22788 ( \23131 , \23129 );
and \U$22789 ( \23132 , \23131 , \2031 );
nor \U$22790 ( \23133 , \23130 , \23132 );
and \U$22791 ( \23134 , \23126 , \23133 );
and \U$22792 ( \23135 , \23117 , \23125 );
or \U$22793 ( \23136 , \23134 , \23135 );
xor \U$22794 ( \23137 , \23110 , \23136 );
xor \U$22795 ( \23138 , \22845 , \22852 );
xor \U$22796 ( \23139 , \23138 , \22861 );
and \U$22797 ( \23140 , \23137 , \23139 );
and \U$22798 ( \23141 , \23110 , \23136 );
nor \U$22799 ( \23142 , \23140 , \23141 );
and \U$22800 ( \23143 , \10424 , RI986e9e0_29);
and \U$22801 ( \23144 , RI986e8f0_27, \10422 );
nor \U$22802 ( \23145 , \23143 , \23144 );
and \U$22803 ( \23146 , \23145 , \9840 );
not \U$22804 ( \23147 , \23145 );
and \U$22805 ( \23148 , \23147 , \10428 );
nor \U$22806 ( \23149 , \23146 , \23148 );
and \U$22807 ( \23150 , \11696 , RI986e800_25);
and \U$22808 ( \23151 , RI986ee90_39, \11694 );
nor \U$22809 ( \23152 , \23150 , \23151 );
and \U$22810 ( \23153 , \23152 , \10965 );
not \U$22811 ( \23154 , \23152 );
and \U$22812 ( \23155 , \23154 , \11702 );
nor \U$22813 ( \23156 , \23153 , \23155 );
xor \U$22814 ( \23157 , \23149 , \23156 );
and \U$22815 ( \23158 , \9505 , RI98715f0_123);
and \U$22816 ( \23159 , RI986ead0_31, \9503 );
nor \U$22817 ( \23160 , \23158 , \23159 );
and \U$22818 ( \23161 , \23160 , \9510 );
not \U$22819 ( \23162 , \23160 );
and \U$22820 ( \23163 , \23162 , \9513 );
nor \U$22821 ( \23164 , \23161 , \23163 );
and \U$22822 ( \23165 , \23157 , \23164 );
and \U$22823 ( \23166 , \23149 , \23156 );
nor \U$22824 ( \23167 , \23165 , \23166 );
not \U$22825 ( \23168 , \23167 );
and \U$22826 ( \23169 , \13045 , RI986ecb0_35);
and \U$22827 ( \23170 , RI986f070_43, \13043 );
nor \U$22828 ( \23171 , \23169 , \23170 );
and \U$22829 ( \23172 , \23171 , \13047 );
not \U$22830 ( \23173 , \23171 );
and \U$22831 ( \23174 , \23173 , \12619 );
nor \U$22832 ( \23175 , \23172 , \23174 );
and \U$22833 ( \23176 , \13882 , RI986ef80_41);
and \U$22834 ( \23177 , RI986f250_47, \13880 );
nor \U$22835 ( \23178 , \23176 , \23177 );
and \U$22836 ( \23179 , \23178 , \13358 );
not \U$22837 ( \23180 , \23178 );
and \U$22838 ( \23181 , \23180 , \13359 );
nor \U$22839 ( \23182 , \23179 , \23181 );
xor \U$22840 ( \23183 , \23175 , \23182 );
and \U$22841 ( \23184 , \12293 , RI986eda0_37);
and \U$22842 ( \23185 , RI986ebc0_33, \12291 );
nor \U$22843 ( \23186 , \23184 , \23185 );
and \U$22844 ( \23187 , \23186 , \11687 );
not \U$22845 ( \23188 , \23186 );
and \U$22846 ( \23189 , \23188 , \11686 );
nor \U$22847 ( \23190 , \23187 , \23189 );
and \U$22848 ( \23191 , \23183 , \23190 );
and \U$22849 ( \23192 , \23175 , \23182 );
nor \U$22850 ( \23193 , \23191 , \23192 );
not \U$22851 ( \23194 , \23193 );
and \U$22852 ( \23195 , \23168 , \23194 );
and \U$22853 ( \23196 , \23167 , \23193 );
not \U$22854 ( \23197 , RI9873558_190);
and \U$22855 ( \23198 , \15780 , RI986e440_17);
and \U$22856 ( \23199 , RI9873648_192, RI986e710_23);
nor \U$22857 ( \23200 , \23198 , \23199 );
not \U$22858 ( \23201 , \23200 );
or \U$22859 ( \23202 , \23197 , \23201 );
or \U$22860 ( \23203 , \23200 , RI9873558_190);
nand \U$22861 ( \23204 , \23202 , \23203 );
and \U$22862 ( \23205 , \23204 , \1337 );
not \U$22863 ( \23206 , \23204 );
not \U$22864 ( \23207 , \1337 );
and \U$22865 ( \23208 , \23206 , \23207 );
and \U$22866 ( \23209 , \14937 , RI986f160_45);
and \U$22867 ( \23210 , RI986e530_19, \14935 );
nor \U$22868 ( \23211 , \23209 , \23210 );
and \U$22869 ( \23212 , \23211 , \14538 );
not \U$22870 ( \23213 , \23211 );
and \U$22871 ( \23214 , \23213 , \14539 );
nor \U$22872 ( \23215 , \23212 , \23214 );
nor \U$22873 ( \23216 , \23208 , \23215 );
nor \U$22874 ( \23217 , \23205 , \23216 );
nor \U$22875 ( \23218 , \23196 , \23217 );
nor \U$22876 ( \23219 , \23195 , \23218 );
or \U$22877 ( \23220 , \23142 , \23219 );
not \U$22878 ( \23221 , \23219 );
not \U$22879 ( \23222 , \23142 );
or \U$22880 ( \23223 , \23221 , \23222 );
and \U$22881 ( \23224 , \7729 , RI9871140_113);
and \U$22882 ( \23225 , RI9871320_117, \7727 );
nor \U$22883 ( \23226 , \23224 , \23225 );
and \U$22884 ( \23227 , \23226 , \7480 );
not \U$22885 ( \23228 , \23226 );
and \U$22886 ( \23229 , \23228 , \7733 );
nor \U$22887 ( \23230 , \23227 , \23229 );
and \U$22888 ( \23231 , \8486 , RI9871410_119);
and \U$22889 ( \23232 , RI98716e0_125, \8484 );
nor \U$22890 ( \23233 , \23231 , \23232 );
and \U$22891 ( \23234 , \23233 , \8050 );
not \U$22892 ( \23235 , \23233 );
and \U$22893 ( \23236 , \23235 , \8051 );
nor \U$22894 ( \23237 , \23234 , \23236 );
xor \U$22895 ( \23238 , \23230 , \23237 );
and \U$22896 ( \23239 , \9237 , RI98717d0_127);
and \U$22897 ( \23240 , RI9871500_121, \9235 );
nor \U$22898 ( \23241 , \23239 , \23240 );
and \U$22899 ( \23242 , \23241 , \9241 );
not \U$22900 ( \23243 , \23241 );
and \U$22901 ( \23244 , \23243 , \8836 );
nor \U$22902 ( \23245 , \23242 , \23244 );
and \U$22903 ( \23246 , \23238 , \23245 );
and \U$22904 ( \23247 , \23230 , \23237 );
or \U$22905 ( \23248 , \23246 , \23247 );
not \U$22906 ( \23249 , \4519 );
and \U$22907 ( \23250 , \4710 , RI9870150_79);
and \U$22908 ( \23251 , RI9870f60_109, \4708 );
nor \U$22909 ( \23252 , \23250 , \23251 );
not \U$22910 ( \23253 , \23252 );
or \U$22911 ( \23254 , \23249 , \23253 );
or \U$22912 ( \23255 , \23252 , \4519 );
nand \U$22913 ( \23256 , \23254 , \23255 );
and \U$22914 ( \23257 , \4203 , RI986fe80_73);
and \U$22915 ( \23258 , RI9870060_77, \4201 );
nor \U$22916 ( \23259 , \23257 , \23258 );
and \U$22917 ( \23260 , \23259 , \4207 );
not \U$22918 ( \23261 , \23259 );
and \U$22919 ( \23262 , \23261 , \3922 );
nor \U$22920 ( \23263 , \23260 , \23262 );
xor \U$22921 ( \23264 , \23256 , \23263 );
and \U$22922 ( \23265 , \5318 , RI9870ab0_99);
and \U$22923 ( \23266 , RI9870d80_105, \5316 );
nor \U$22924 ( \23267 , \23265 , \23266 );
and \U$22925 ( \23268 , \23267 , \5052 );
not \U$22926 ( \23269 , \23267 );
and \U$22927 ( \23270 , \23269 , \5322 );
nor \U$22928 ( \23271 , \23268 , \23270 );
and \U$22929 ( \23272 , \23264 , \23271 );
and \U$22930 ( \23273 , \23256 , \23263 );
or \U$22931 ( \23274 , \23272 , \23273 );
xor \U$22932 ( \23275 , \23248 , \23274 );
and \U$22933 ( \23276 , \5881 , RI98709c0_97);
and \U$22934 ( \23277 , RI9870e70_107, \5879 );
nor \U$22935 ( \23278 , \23276 , \23277 );
and \U$22936 ( \23279 , \23278 , \5594 );
not \U$22937 ( \23280 , \23278 );
and \U$22938 ( \23281 , \23280 , \5885 );
nor \U$22939 ( \23282 , \23279 , \23281 );
and \U$22940 ( \23283 , \6453 , RI9870ba0_101);
and \U$22941 ( \23284 , RI9871050_111, \6451 );
nor \U$22942 ( \23285 , \23283 , \23284 );
and \U$22943 ( \23286 , \23285 , \6190 );
not \U$22944 ( \23287 , \23285 );
and \U$22945 ( \23288 , \23287 , \6705 );
nor \U$22946 ( \23289 , \23286 , \23288 );
xor \U$22947 ( \23290 , \23282 , \23289 );
and \U$22948 ( \23291 , \7079 , RI9870c90_103);
and \U$22949 ( \23292 , RI9871230_115, \7077 );
nor \U$22950 ( \23293 , \23291 , \23292 );
and \U$22951 ( \23294 , \23293 , \6710 );
not \U$22952 ( \23295 , \23293 );
and \U$22953 ( \23296 , \23295 , \6709 );
nor \U$22954 ( \23297 , \23294 , \23296 );
and \U$22955 ( \23298 , \23290 , \23297 );
and \U$22956 ( \23299 , \23282 , \23289 );
or \U$22957 ( \23300 , \23298 , \23299 );
and \U$22958 ( \23301 , \23275 , \23300 );
and \U$22959 ( \23302 , \23248 , \23274 );
or \U$22960 ( \23303 , \23301 , \23302 );
nand \U$22961 ( \23304 , \23223 , \23303 );
nand \U$22962 ( \23305 , \23220 , \23304 );
xor \U$22963 ( \23306 , \23083 , \23305 );
xor \U$22964 ( \23307 , \22830 , \22837 );
xor \U$22965 ( \23308 , \23307 , \22864 );
xor \U$22966 ( \23309 , \22696 , \22702 );
xor \U$22967 ( \23310 , \23309 , \22705 );
and \U$22968 ( \23311 , \23308 , \23310 );
xor \U$22969 ( \23312 , \22578 , \22585 );
xor \U$22970 ( \23313 , \23312 , \22593 );
xor \U$22971 ( \23314 , \22711 , \22716 );
xor \U$22972 ( \23315 , \23313 , \23314 );
xor \U$22973 ( \23316 , \22696 , \22702 );
xor \U$22974 ( \23317 , \23316 , \22705 );
and \U$22975 ( \23318 , \23315 , \23317 );
and \U$22976 ( \23319 , \23308 , \23315 );
or \U$22977 ( \23320 , \23311 , \23318 , \23319 );
and \U$22978 ( \23321 , \23306 , \23320 );
and \U$22979 ( \23322 , \23083 , \23305 );
or \U$22980 ( \23323 , \23321 , \23322 );
xor \U$22981 ( \23324 , \22388 , \22393 );
xor \U$22982 ( \23325 , \23324 , \22404 );
xor \U$22983 ( \23326 , \23323 , \23325 );
xor \U$22984 ( \23327 , \22432 , \22451 );
xor \U$22985 ( \23328 , \23327 , \22477 );
xor \U$22986 ( \23329 , \22985 , \22990 );
xor \U$22987 ( \23330 , \23328 , \23329 );
xor \U$22988 ( \23331 , \22694 , \22708 );
xor \U$22989 ( \23332 , \23331 , \22721 );
and \U$22990 ( \23333 , \23330 , \23332 );
xor \U$22991 ( \23334 , \22396 , \22398 );
xor \U$22992 ( \23335 , \23334 , \22401 );
xor \U$22993 ( \23336 , \22954 , \22961 );
xor \U$22994 ( \23337 , \23335 , \23336 );
xor \U$22995 ( \23338 , \22694 , \22708 );
xor \U$22996 ( \23339 , \23338 , \22721 );
and \U$22997 ( \23340 , \23337 , \23339 );
and \U$22998 ( \23341 , \23330 , \23337 );
or \U$22999 ( \23342 , \23333 , \23340 , \23341 );
and \U$23000 ( \23343 , \23326 , \23342 );
and \U$23001 ( \23344 , \23323 , \23325 );
or \U$23002 ( \23345 , \23343 , \23344 );
xor \U$23003 ( \23346 , \23053 , \23345 );
xor \U$23004 ( \23347 , \22407 , \22629 );
xor \U$23005 ( \23348 , \23347 , \22649 );
xor \U$23006 ( \23349 , \23012 , \23019 );
xor \U$23007 ( \23350 , \23348 , \23349 );
and \U$23008 ( \23351 , \23346 , \23350 );
and \U$23009 ( \23352 , \23053 , \23345 );
or \U$23010 ( \23353 , \23351 , \23352 );
and \U$23011 ( \23354 , \23041 , \23353 );
and \U$23012 ( \23355 , \23038 , \23040 );
nor \U$23013 ( \23356 , \23354 , \23355 );
or \U$23014 ( \23357 , \23037 , \23356 );
xnor \U$23015 ( \23358 , \23037 , \23356 );
xor \U$23016 ( \23359 , \23038 , \23040 );
xor \U$23017 ( \23360 , \23359 , \23353 );
xor \U$23018 ( \23361 , \23043 , \23045 );
xor \U$23019 ( \23362 , \23361 , \23050 );
xor \U$23020 ( \23363 , \22804 , \22867 );
xor \U$23021 ( \23364 , \23363 , \22949 );
xor \U$23022 ( \23365 , \23083 , \23305 );
xor \U$23023 ( \23366 , \23365 , \23320 );
and \U$23024 ( \23367 , \23364 , \23366 );
xor \U$23025 ( \23368 , \22694 , \22708 );
xor \U$23026 ( \23369 , \23368 , \22721 );
xor \U$23027 ( \23370 , \23330 , \23337 );
xor \U$23028 ( \23371 , \23369 , \23370 );
xor \U$23029 ( \23372 , \23083 , \23305 );
xor \U$23030 ( \23373 , \23372 , \23320 );
and \U$23031 ( \23374 , \23371 , \23373 );
and \U$23032 ( \23375 , \23364 , \23371 );
or \U$23033 ( \23376 , \23367 , \23374 , \23375 );
and \U$23034 ( \23377 , \23362 , \23376 );
not \U$23035 ( \23378 , \23362 );
not \U$23036 ( \23379 , \23376 );
and \U$23037 ( \23380 , \23378 , \23379 );
xor \U$23038 ( \23381 , \22893 , \22918 );
xor \U$23039 ( \23382 , \23381 , \22946 );
xor \U$23040 ( \23383 , \22749 , \22775 );
xor \U$23041 ( \23384 , \23383 , \22801 );
xor \U$23042 ( \23385 , \23382 , \23384 );
xor \U$23043 ( \23386 , \22696 , \22702 );
xor \U$23044 ( \23387 , \23386 , \22705 );
xor \U$23045 ( \23388 , \23308 , \23315 );
xor \U$23046 ( \23389 , \23387 , \23388 );
and \U$23047 ( \23390 , \23385 , \23389 );
and \U$23048 ( \23391 , \23382 , \23384 );
or \U$23049 ( \23392 , \23390 , \23391 );
not \U$23050 ( \23393 , \23392 );
not \U$23051 ( \23394 , \23393 );
not \U$23052 ( \23395 , \23219 );
not \U$23053 ( \23396 , \23303 );
or \U$23054 ( \23397 , \23395 , \23396 );
or \U$23055 ( \23398 , \23303 , \23219 );
nand \U$23056 ( \23399 , \23397 , \23398 );
not \U$23057 ( \23400 , \23399 );
not \U$23058 ( \23401 , \23142 );
and \U$23059 ( \23402 , \23400 , \23401 );
and \U$23060 ( \23403 , \23399 , \23142 );
nor \U$23061 ( \23404 , \23402 , \23403 );
not \U$23062 ( \23405 , \23404 );
xor \U$23063 ( \23406 , \23065 , \23075 );
xor \U$23064 ( \23407 , \23406 , \23080 );
nand \U$23065 ( \23408 , \23405 , \23407 );
not \U$23066 ( \23409 , \23408 );
and \U$23067 ( \23410 , \23394 , \23409 );
and \U$23068 ( \23411 , \23393 , \23408 );
xor \U$23069 ( \23412 , \23230 , \23237 );
xor \U$23070 ( \23413 , \23412 , \23245 );
xor \U$23071 ( \23414 , \23149 , \23156 );
xor \U$23072 ( \23415 , \23414 , \23164 );
xor \U$23073 ( \23416 , \23413 , \23415 );
xor \U$23074 ( \23417 , \23175 , \23182 );
xor \U$23075 ( \23418 , \23417 , \23190 );
and \U$23076 ( \23419 , \23416 , \23418 );
and \U$23077 ( \23420 , \23413 , \23415 );
or \U$23078 ( \23421 , \23419 , \23420 );
xor \U$23079 ( \23422 , \22756 , \22764 );
xor \U$23080 ( \23423 , \23422 , \22772 );
xor \U$23081 ( \23424 , \23421 , \23423 );
xor \U$23082 ( \23425 , \23091 , \23098 );
xor \U$23083 ( \23426 , \23425 , \23107 );
xor \U$23084 ( \23427 , \23282 , \23289 );
xor \U$23085 ( \23428 , \23427 , \23297 );
and \U$23086 ( \23429 , \23426 , \23428 );
xor \U$23087 ( \23430 , \23256 , \23263 );
xor \U$23088 ( \23431 , \23430 , \23271 );
xor \U$23089 ( \23432 , \23282 , \23289 );
xor \U$23090 ( \23433 , \23432 , \23297 );
and \U$23091 ( \23434 , \23431 , \23433 );
and \U$23092 ( \23435 , \23426 , \23431 );
or \U$23093 ( \23436 , \23429 , \23434 , \23435 );
and \U$23094 ( \23437 , \23424 , \23436 );
and \U$23095 ( \23438 , \23421 , \23423 );
or \U$23096 ( \23439 , \23437 , \23438 );
and \U$23097 ( \23440 , \8486 , RI9871320_117);
and \U$23098 ( \23441 , RI9871410_119, \8484 );
nor \U$23099 ( \23442 , \23440 , \23441 );
and \U$23100 ( \23443 , \23442 , \8050 );
not \U$23101 ( \23444 , \23442 );
and \U$23102 ( \23445 , \23444 , \8051 );
nor \U$23103 ( \23446 , \23443 , \23445 );
and \U$23104 ( \23447 , \7079 , RI9871050_111);
and \U$23105 ( \23448 , RI9870c90_103, \7077 );
nor \U$23106 ( \23449 , \23447 , \23448 );
and \U$23107 ( \23450 , \23449 , \6710 );
not \U$23108 ( \23451 , \23449 );
and \U$23109 ( \23452 , \23451 , \6709 );
nor \U$23110 ( \23453 , \23450 , \23452 );
xor \U$23111 ( \23454 , \23446 , \23453 );
and \U$23112 ( \23455 , \7729 , RI9871230_115);
and \U$23113 ( \23456 , RI9871140_113, \7727 );
nor \U$23114 ( \23457 , \23455 , \23456 );
and \U$23115 ( \23458 , \23457 , \7480 );
not \U$23116 ( \23459 , \23457 );
and \U$23117 ( \23460 , \23459 , \7733 );
nor \U$23118 ( \23461 , \23458 , \23460 );
and \U$23119 ( \23462 , \23454 , \23461 );
and \U$23120 ( \23463 , \23446 , \23453 );
or \U$23121 ( \23464 , \23462 , \23463 );
not \U$23122 ( \23465 , \3918 );
and \U$23123 ( \23466 , \3683 , RI986fd90_71);
and \U$23124 ( \23467 , RI986fca0_69, \3681 );
nor \U$23125 ( \23468 , \23466 , \23467 );
not \U$23126 ( \23469 , \23468 );
or \U$23127 ( \23470 , \23465 , \23469 );
or \U$23128 ( \23471 , \23468 , \3918 );
nand \U$23129 ( \23472 , \23470 , \23471 );
and \U$23130 ( \23473 , \4203 , RI986ff70_75);
and \U$23131 ( \23474 , RI986fe80_73, \4201 );
nor \U$23132 ( \23475 , \23473 , \23474 );
and \U$23133 ( \23476 , \23475 , \4207 );
not \U$23134 ( \23477 , \23475 );
and \U$23135 ( \23478 , \23477 , \3922 );
nor \U$23136 ( \23479 , \23476 , \23478 );
xor \U$23137 ( \23480 , \23472 , \23479 );
not \U$23138 ( \23481 , \4519 );
and \U$23139 ( \23482 , \4710 , RI9870060_77);
and \U$23140 ( \23483 , RI9870150_79, \4708 );
nor \U$23141 ( \23484 , \23482 , \23483 );
not \U$23142 ( \23485 , \23484 );
or \U$23143 ( \23486 , \23481 , \23485 );
or \U$23144 ( \23487 , \23484 , \4519 );
nand \U$23145 ( \23488 , \23486 , \23487 );
and \U$23146 ( \23489 , \23480 , \23488 );
and \U$23147 ( \23490 , \23472 , \23479 );
or \U$23148 ( \23491 , \23489 , \23490 );
xor \U$23149 ( \23492 , \23464 , \23491 );
and \U$23150 ( \23493 , \6453 , RI9870e70_107);
and \U$23151 ( \23494 , RI9870ba0_101, \6451 );
nor \U$23152 ( \23495 , \23493 , \23494 );
and \U$23153 ( \23496 , \23495 , \6190 );
not \U$23154 ( \23497 , \23495 );
and \U$23155 ( \23498 , \23497 , \6180 );
nor \U$23156 ( \23499 , \23496 , \23498 );
and \U$23157 ( \23500 , \5318 , RI9870f60_109);
and \U$23158 ( \23501 , RI9870ab0_99, \5316 );
nor \U$23159 ( \23502 , \23500 , \23501 );
and \U$23160 ( \23503 , \23502 , \5052 );
not \U$23161 ( \23504 , \23502 );
and \U$23162 ( \23505 , \23504 , \5322 );
nor \U$23163 ( \23506 , \23503 , \23505 );
xor \U$23164 ( \23507 , \23499 , \23506 );
and \U$23165 ( \23508 , \5881 , RI9870d80_105);
and \U$23166 ( \23509 , RI98709c0_97, \5879 );
nor \U$23167 ( \23510 , \23508 , \23509 );
and \U$23168 ( \23511 , \23510 , \5594 );
not \U$23169 ( \23512 , \23510 );
and \U$23170 ( \23513 , \23512 , \5885 );
nor \U$23171 ( \23514 , \23511 , \23513 );
and \U$23172 ( \23515 , \23507 , \23514 );
and \U$23173 ( \23516 , \23499 , \23506 );
or \U$23174 ( \23517 , \23515 , \23516 );
and \U$23175 ( \23518 , \23492 , \23517 );
and \U$23176 ( \23519 , \23464 , \23491 );
or \U$23177 ( \23520 , \23518 , \23519 );
and \U$23178 ( \23521 , \11696 , RI986e8f0_27);
and \U$23179 ( \23522 , RI986e800_25, \11694 );
nor \U$23180 ( \23523 , \23521 , \23522 );
and \U$23181 ( \23524 , \23523 , \10965 );
not \U$23182 ( \23525 , \23523 );
and \U$23183 ( \23526 , \23525 , \11702 );
nor \U$23184 ( \23527 , \23524 , \23526 );
and \U$23185 ( \23528 , \12293 , RI986ee90_39);
and \U$23186 ( \23529 , RI986eda0_37, \12291 );
nor \U$23187 ( \23530 , \23528 , \23529 );
and \U$23188 ( \23531 , \23530 , \11687 );
not \U$23189 ( \23532 , \23530 );
and \U$23190 ( \23533 , \23532 , \11686 );
nor \U$23191 ( \23534 , \23531 , \23533 );
xor \U$23192 ( \23535 , \23527 , \23534 );
and \U$23193 ( \23536 , \13045 , RI986ebc0_33);
and \U$23194 ( \23537 , RI986ecb0_35, \13043 );
nor \U$23195 ( \23538 , \23536 , \23537 );
and \U$23196 ( \23539 , \23538 , \13047 );
not \U$23197 ( \23540 , \23538 );
and \U$23198 ( \23541 , \23540 , \12619 );
nor \U$23199 ( \23542 , \23539 , \23541 );
and \U$23200 ( \23543 , \23535 , \23542 );
and \U$23201 ( \23544 , \23527 , \23534 );
or \U$23202 ( \23545 , \23543 , \23544 );
and \U$23203 ( \23546 , \13882 , RI986f070_43);
and \U$23204 ( \23547 , RI986ef80_41, \13880 );
nor \U$23205 ( \23548 , \23546 , \23547 );
and \U$23206 ( \23549 , \23548 , \13358 );
not \U$23207 ( \23550 , \23548 );
and \U$23208 ( \23551 , \23550 , \13359 );
nor \U$23209 ( \23552 , \23549 , \23551 );
not \U$23210 ( \23553 , RI9873558_190);
and \U$23211 ( \23554 , \15780 , RI986e530_19);
and \U$23212 ( \23555 , RI9873648_192, RI986e440_17);
nor \U$23213 ( \23556 , \23554 , \23555 );
not \U$23214 ( \23557 , \23556 );
or \U$23215 ( \23558 , \23553 , \23557 );
or \U$23216 ( \23559 , \23556 , RI9873558_190);
nand \U$23217 ( \23560 , \23558 , \23559 );
xor \U$23218 ( \23561 , \23552 , \23560 );
and \U$23219 ( \23562 , \14937 , RI986f250_47);
and \U$23220 ( \23563 , RI986f160_45, \14935 );
nor \U$23221 ( \23564 , \23562 , \23563 );
and \U$23222 ( \23565 , \23564 , \14539 );
not \U$23223 ( \23566 , \23564 );
and \U$23224 ( \23567 , \23566 , \14538 );
nor \U$23225 ( \23568 , \23565 , \23567 );
and \U$23226 ( \23569 , \23561 , \23568 );
and \U$23227 ( \23570 , \23552 , \23560 );
or \U$23228 ( \23571 , \23569 , \23570 );
xor \U$23229 ( \23572 , \23545 , \23571 );
and \U$23230 ( \23573 , \10424 , RI986ead0_31);
and \U$23231 ( \23574 , RI986e9e0_29, \10422 );
nor \U$23232 ( \23575 , \23573 , \23574 );
and \U$23233 ( \23576 , \23575 , \9840 );
not \U$23234 ( \23577 , \23575 );
and \U$23235 ( \23578 , \23577 , \10428 );
nor \U$23236 ( \23579 , \23576 , \23578 );
and \U$23237 ( \23580 , \9237 , RI98716e0_125);
and \U$23238 ( \23581 , RI98717d0_127, \9235 );
nor \U$23239 ( \23582 , \23580 , \23581 );
and \U$23240 ( \23583 , \23582 , \9241 );
not \U$23241 ( \23584 , \23582 );
and \U$23242 ( \23585 , \23584 , \8836 );
nor \U$23243 ( \23586 , \23583 , \23585 );
xor \U$23244 ( \23587 , \23579 , \23586 );
and \U$23245 ( \23588 , \9505 , RI9871500_121);
and \U$23246 ( \23589 , RI98715f0_123, \9503 );
nor \U$23247 ( \23590 , \23588 , \23589 );
and \U$23248 ( \23591 , \23590 , \9510 );
not \U$23249 ( \23592 , \23590 );
and \U$23250 ( \23593 , \23592 , \9513 );
nor \U$23251 ( \23594 , \23591 , \23593 );
and \U$23252 ( \23595 , \23587 , \23594 );
and \U$23253 ( \23596 , \23579 , \23586 );
or \U$23254 ( \23597 , \23595 , \23596 );
and \U$23255 ( \23598 , \23572 , \23597 );
and \U$23256 ( \23599 , \23545 , \23571 );
or \U$23257 ( \23600 , \23598 , \23599 );
xor \U$23258 ( \23601 , \23520 , \23600 );
and \U$23259 ( \23602 , \2274 , RI98706f0_91);
and \U$23260 ( \23603 , RI9870600_89, \2272 );
nor \U$23261 ( \23604 , \23602 , \23603 );
and \U$23262 ( \23605 , \23604 , \2030 );
not \U$23263 ( \23606 , \23604 );
and \U$23264 ( \23607 , \23606 , \2031 );
nor \U$23265 ( \23608 , \23605 , \23607 );
and \U$23266 ( \23609 , \2464 , RI98708d0_95);
and \U$23267 ( \23610 , RI98707e0_93, \2462 );
nor \U$23268 ( \23611 , \23609 , \23610 );
and \U$23269 ( \23612 , \23611 , \2468 );
not \U$23270 ( \23613 , \23611 );
and \U$23271 ( \23614 , \23613 , \2263 );
nor \U$23272 ( \23615 , \23612 , \23614 );
xor \U$23273 ( \23616 , \23608 , \23615 );
not \U$23274 ( \23617 , \3406 );
and \U$23275 ( \23618 , \3254 , RI986fac0_65);
and \U$23276 ( \23619 , RI986fbb0_67, \3252 );
nor \U$23277 ( \23620 , \23618 , \23619 );
not \U$23278 ( \23621 , \23620 );
or \U$23279 ( \23622 , \23617 , \23621 );
or \U$23280 ( \23623 , \23620 , \3406 );
nand \U$23281 ( \23624 , \23622 , \23623 );
and \U$23282 ( \23625 , \23616 , \23624 );
and \U$23283 ( \23626 , \23608 , \23615 );
or \U$23284 ( \23627 , \23625 , \23626 );
nand \U$23285 ( \23628 , RI9870420_85, \1327 );
and \U$23286 ( \23629 , \23628 , \1336 );
not \U$23287 ( \23630 , \23628 );
and \U$23288 ( \23631 , \23630 , \1337 );
nor \U$23289 ( \23632 , \23629 , \23631 );
xor \U$23290 ( \23633 , \23627 , \23632 );
xor \U$23291 ( \23634 , \23117 , \23125 );
xor \U$23292 ( \23635 , \23634 , \23133 );
and \U$23293 ( \23636 , \23633 , \23635 );
and \U$23294 ( \23637 , \23627 , \23632 );
or \U$23295 ( \23638 , \23636 , \23637 );
and \U$23296 ( \23639 , \23601 , \23638 );
and \U$23297 ( \23640 , \23520 , \23600 );
or \U$23298 ( \23641 , \23639 , \23640 );
xor \U$23299 ( \23642 , \23439 , \23641 );
xor \U$23300 ( \23643 , \23110 , \23136 );
xor \U$23301 ( \23644 , \23643 , \23139 );
xor \U$23302 ( \23645 , \23067 , \23069 );
xor \U$23303 ( \23646 , \23645 , \23072 );
and \U$23304 ( \23647 , \23644 , \23646 );
xor \U$23305 ( \23648 , \22811 , \22818 );
xor \U$23306 ( \23649 , \23648 , \22827 );
xor \U$23307 ( \23650 , \23055 , \23060 );
xor \U$23308 ( \23651 , \23649 , \23650 );
xor \U$23309 ( \23652 , \23067 , \23069 );
xor \U$23310 ( \23653 , \23652 , \23072 );
and \U$23311 ( \23654 , \23651 , \23653 );
and \U$23312 ( \23655 , \23644 , \23651 );
or \U$23313 ( \23656 , \23647 , \23654 , \23655 );
and \U$23314 ( \23657 , \23642 , \23656 );
and \U$23315 ( \23658 , \23439 , \23641 );
or \U$23316 ( \23659 , \23657 , \23658 );
not \U$23317 ( \23660 , \23659 );
nor \U$23318 ( \23661 , \23411 , \23660 );
nor \U$23319 ( \23662 , \23410 , \23661 );
nor \U$23320 ( \23663 , \23380 , \23662 );
nor \U$23321 ( \23664 , \23377 , \23663 );
not \U$23322 ( \23665 , \22969 );
not \U$23323 ( \23666 , \23005 );
or \U$23324 ( \23667 , \23665 , \23666 );
or \U$23325 ( \23668 , \23005 , \22969 );
nand \U$23326 ( \23669 , \23667 , \23668 );
not \U$23327 ( \23670 , \23669 );
not \U$23328 ( \23671 , \22979 );
and \U$23329 ( \23672 , \23670 , \23671 );
and \U$23330 ( \23673 , \23669 , \22979 );
nor \U$23331 ( \23674 , \23672 , \23673 );
or \U$23332 ( \23675 , \23664 , \23674 );
not \U$23333 ( \23676 , \23674 );
not \U$23334 ( \23677 , \23664 );
or \U$23335 ( \23678 , \23676 , \23677 );
xor \U$23336 ( \23679 , \23053 , \23345 );
xor \U$23337 ( \23680 , \23679 , \23350 );
nand \U$23338 ( \23681 , \23678 , \23680 );
nand \U$23339 ( \23682 , \23675 , \23681 );
and \U$23340 ( \23683 , \23360 , \23682 );
xor \U$23341 ( \23684 , \23682 , \23360 );
not \U$23342 ( \23685 , \23362 );
not \U$23343 ( \23686 , \23376 );
not \U$23344 ( \23687 , \23662 );
and \U$23345 ( \23688 , \23686 , \23687 );
and \U$23346 ( \23689 , \23376 , \23662 );
nor \U$23347 ( \23690 , \23688 , \23689 );
not \U$23348 ( \23691 , \23690 );
or \U$23349 ( \23692 , \23685 , \23691 );
or \U$23350 ( \23693 , \23690 , \23362 );
nand \U$23351 ( \23694 , \23692 , \23693 );
xor \U$23352 ( \23695 , \23323 , \23325 );
xor \U$23353 ( \23696 , \23695 , \23342 );
xor \U$23354 ( \23697 , \23694 , \23696 );
not \U$23355 ( \23698 , \23404 );
not \U$23356 ( \23699 , \23407 );
or \U$23357 ( \23700 , \23698 , \23699 );
or \U$23358 ( \23701 , \23407 , \23404 );
nand \U$23359 ( \23702 , \23700 , \23701 );
xor \U$23360 ( \23703 , \23382 , \23384 );
xor \U$23361 ( \23704 , \23703 , \23389 );
and \U$23362 ( \23705 , \23702 , \23704 );
xor \U$23363 ( \23706 , \23439 , \23641 );
xor \U$23364 ( \23707 , \23706 , \23656 );
xor \U$23365 ( \23708 , \23382 , \23384 );
xor \U$23366 ( \23709 , \23708 , \23389 );
and \U$23367 ( \23710 , \23707 , \23709 );
and \U$23368 ( \23711 , \23702 , \23707 );
or \U$23369 ( \23712 , \23705 , \23710 , \23711 );
xor \U$23370 ( \23713 , \23608 , \23615 );
xor \U$23371 ( \23714 , \23713 , \23624 );
and \U$23372 ( \23715 , \1311 , RI9870420_85);
and \U$23373 ( \23716 , RI9870510_87, \1309 );
nor \U$23374 ( \23717 , \23715 , \23716 );
and \U$23375 ( \23718 , \23717 , \1319 );
not \U$23376 ( \23719 , \23717 );
and \U$23377 ( \23720 , \23719 , \1315 );
nor \U$23378 ( \23721 , \23718 , \23720 );
xor \U$23379 ( \23722 , \23714 , \23721 );
xor \U$23380 ( \23723 , \23472 , \23479 );
xor \U$23381 ( \23724 , \23723 , \23488 );
and \U$23382 ( \23725 , \23722 , \23724 );
and \U$23383 ( \23726 , \23714 , \23721 );
or \U$23384 ( \23727 , \23725 , \23726 );
not \U$23385 ( \23728 , \1336 );
not \U$23386 ( \23729 , \23204 );
not \U$23387 ( \23730 , \23215 );
or \U$23388 ( \23731 , \23729 , \23730 );
or \U$23389 ( \23732 , \23215 , \23204 );
nand \U$23390 ( \23733 , \23731 , \23732 );
not \U$23391 ( \23734 , \23733 );
or \U$23392 ( \23735 , \23728 , \23734 );
or \U$23393 ( \23736 , \23733 , \1336 );
nand \U$23394 ( \23737 , \23735 , \23736 );
xor \U$23395 ( \23738 , \23727 , \23737 );
xor \U$23396 ( \23739 , \23499 , \23506 );
xor \U$23397 ( \23740 , \23739 , \23514 );
xor \U$23398 ( \23741 , \23446 , \23453 );
xor \U$23399 ( \23742 , \23741 , \23461 );
and \U$23400 ( \23743 , \23740 , \23742 );
xor \U$23401 ( \23744 , \23579 , \23586 );
xor \U$23402 ( \23745 , \23744 , \23594 );
xor \U$23403 ( \23746 , \23446 , \23453 );
xor \U$23404 ( \23747 , \23746 , \23461 );
and \U$23405 ( \23748 , \23745 , \23747 );
and \U$23406 ( \23749 , \23740 , \23745 );
or \U$23407 ( \23750 , \23743 , \23748 , \23749 );
and \U$23408 ( \23751 , \23738 , \23750 );
and \U$23409 ( \23752 , \23727 , \23737 );
or \U$23410 ( \23753 , \23751 , \23752 );
and \U$23411 ( \23754 , \10424 , RI98715f0_123);
and \U$23412 ( \23755 , RI986ead0_31, \10422 );
nor \U$23413 ( \23756 , \23754 , \23755 );
and \U$23414 ( \23757 , \23756 , \9840 );
not \U$23415 ( \23758 , \23756 );
and \U$23416 ( \23759 , \23758 , \10428 );
nor \U$23417 ( \23760 , \23757 , \23759 );
and \U$23418 ( \23761 , \9505 , RI98717d0_127);
and \U$23419 ( \23762 , RI9871500_121, \9503 );
nor \U$23420 ( \23763 , \23761 , \23762 );
and \U$23421 ( \23764 , \23763 , \9510 );
not \U$23422 ( \23765 , \23763 );
and \U$23423 ( \23766 , \23765 , \9513 );
nor \U$23424 ( \23767 , \23764 , \23766 );
xor \U$23425 ( \23768 , \23760 , \23767 );
and \U$23426 ( \23769 , \11696 , RI986e9e0_29);
and \U$23427 ( \23770 , RI986e8f0_27, \11694 );
nor \U$23428 ( \23771 , \23769 , \23770 );
and \U$23429 ( \23772 , \23771 , \10965 );
not \U$23430 ( \23773 , \23771 );
and \U$23431 ( \23774 , \23773 , \11702 );
nor \U$23432 ( \23775 , \23772 , \23774 );
and \U$23433 ( \23776 , \23768 , \23775 );
and \U$23434 ( \23777 , \23760 , \23767 );
or \U$23435 ( \23778 , \23776 , \23777 );
not \U$23436 ( \23779 , RI9873558_190);
and \U$23437 ( \23780 , \15780 , RI986f160_45);
and \U$23438 ( \23781 , RI9873648_192, RI986e530_19);
nor \U$23439 ( \23782 , \23780 , \23781 );
not \U$23440 ( \23783 , \23782 );
or \U$23441 ( \23784 , \23779 , \23783 );
or \U$23442 ( \23785 , \23782 , RI9873558_190);
nand \U$23443 ( \23786 , \23784 , \23785 );
xor \U$23444 ( \23787 , \23786 , \1315 );
and \U$23445 ( \23788 , \14937 , RI986ef80_41);
and \U$23446 ( \23789 , RI986f250_47, \14935 );
nor \U$23447 ( \23790 , \23788 , \23789 );
and \U$23448 ( \23791 , \23790 , \14539 );
not \U$23449 ( \23792 , \23790 );
and \U$23450 ( \23793 , \23792 , \14538 );
nor \U$23451 ( \23794 , \23791 , \23793 );
and \U$23452 ( \23795 , \23787 , \23794 );
and \U$23453 ( \23796 , \23786 , \1315 );
or \U$23454 ( \23797 , \23795 , \23796 );
xor \U$23455 ( \23798 , \23778 , \23797 );
and \U$23456 ( \23799 , \12293 , RI986e800_25);
and \U$23457 ( \23800 , RI986ee90_39, \12291 );
nor \U$23458 ( \23801 , \23799 , \23800 );
and \U$23459 ( \23802 , \23801 , \11687 );
not \U$23460 ( \23803 , \23801 );
and \U$23461 ( \23804 , \23803 , \11686 );
nor \U$23462 ( \23805 , \23802 , \23804 );
and \U$23463 ( \23806 , \13045 , RI986eda0_37);
and \U$23464 ( \23807 , RI986ebc0_33, \13043 );
nor \U$23465 ( \23808 , \23806 , \23807 );
and \U$23466 ( \23809 , \23808 , \13047 );
not \U$23467 ( \23810 , \23808 );
and \U$23468 ( \23811 , \23810 , \12619 );
nor \U$23469 ( \23812 , \23809 , \23811 );
xor \U$23470 ( \23813 , \23805 , \23812 );
and \U$23471 ( \23814 , \13882 , RI986ecb0_35);
and \U$23472 ( \23815 , RI986f070_43, \13880 );
nor \U$23473 ( \23816 , \23814 , \23815 );
and \U$23474 ( \23817 , \23816 , \13358 );
not \U$23475 ( \23818 , \23816 );
and \U$23476 ( \23819 , \23818 , \13359 );
nor \U$23477 ( \23820 , \23817 , \23819 );
and \U$23478 ( \23821 , \23813 , \23820 );
and \U$23479 ( \23822 , \23805 , \23812 );
or \U$23480 ( \23823 , \23821 , \23822 );
and \U$23481 ( \23824 , \23798 , \23823 );
and \U$23482 ( \23825 , \23778 , \23797 );
or \U$23483 ( \23826 , \23824 , \23825 );
and \U$23484 ( \23827 , \2274 , RI9870240_81);
and \U$23485 ( \23828 , RI98706f0_91, \2272 );
nor \U$23486 ( \23829 , \23827 , \23828 );
and \U$23487 ( \23830 , \23829 , \2030 );
not \U$23488 ( \23831 , \23829 );
and \U$23489 ( \23832 , \23831 , \2031 );
nor \U$23490 ( \23833 , \23830 , \23832 );
nand \U$23491 ( \23834 , RI9870420_85, \1309 );
and \U$23492 ( \23835 , \23834 , \1458 );
not \U$23493 ( \23836 , \23834 );
and \U$23494 ( \23837 , \23836 , \1315 );
nor \U$23495 ( \23838 , \23835 , \23837 );
xor \U$23496 ( \23839 , \23833 , \23838 );
not \U$23497 ( \23840 , \1462 );
and \U$23498 ( \23841 , \2042 , RI9870510_87);
and \U$23499 ( \23842 , RI9870330_83, \2040 );
nor \U$23500 ( \23843 , \23841 , \23842 );
not \U$23501 ( \23844 , \23843 );
or \U$23502 ( \23845 , \23840 , \23844 );
or \U$23503 ( \23846 , \23843 , \1462 );
nand \U$23504 ( \23847 , \23845 , \23846 );
and \U$23505 ( \23848 , \23839 , \23847 );
and \U$23506 ( \23849 , \23833 , \23838 );
or \U$23507 ( \23850 , \23848 , \23849 );
not \U$23508 ( \23851 , \1462 );
and \U$23509 ( \23852 , \2042 , RI9870330_83);
and \U$23510 ( \23853 , RI9870240_81, \2040 );
nor \U$23511 ( \23854 , \23852 , \23853 );
not \U$23512 ( \23855 , \23854 );
or \U$23513 ( \23856 , \23851 , \23855 );
or \U$23514 ( \23857 , \23854 , \2034 );
nand \U$23515 ( \23858 , \23856 , \23857 );
xor \U$23516 ( \23859 , \23850 , \23858 );
and \U$23517 ( \23860 , \2464 , RI9870600_89);
and \U$23518 ( \23861 , RI98708d0_95, \2462 );
nor \U$23519 ( \23862 , \23860 , \23861 );
and \U$23520 ( \23863 , \23862 , \2468 );
not \U$23521 ( \23864 , \23862 );
and \U$23522 ( \23865 , \23864 , \2263 );
nor \U$23523 ( \23866 , \23863 , \23865 );
not \U$23524 ( \23867 , \3406 );
and \U$23525 ( \23868 , \3254 , RI98707e0_93);
and \U$23526 ( \23869 , RI986fac0_65, \3252 );
nor \U$23527 ( \23870 , \23868 , \23869 );
not \U$23528 ( \23871 , \23870 );
or \U$23529 ( \23872 , \23867 , \23871 );
or \U$23530 ( \23873 , \23870 , \2935 );
nand \U$23531 ( \23874 , \23872 , \23873 );
xor \U$23532 ( \23875 , \23866 , \23874 );
not \U$23533 ( \23876 , \3412 );
and \U$23534 ( \23877 , \3683 , RI986fbb0_67);
and \U$23535 ( \23878 , RI986fd90_71, \3681 );
nor \U$23536 ( \23879 , \23877 , \23878 );
not \U$23537 ( \23880 , \23879 );
or \U$23538 ( \23881 , \23876 , \23880 );
or \U$23539 ( \23882 , \23879 , \3412 );
nand \U$23540 ( \23883 , \23881 , \23882 );
and \U$23541 ( \23884 , \23875 , \23883 );
and \U$23542 ( \23885 , \23866 , \23874 );
or \U$23543 ( \23886 , \23884 , \23885 );
and \U$23544 ( \23887 , \23859 , \23886 );
and \U$23545 ( \23888 , \23850 , \23858 );
or \U$23546 ( \23889 , \23887 , \23888 );
xor \U$23547 ( \23890 , \23826 , \23889 );
and \U$23548 ( \23891 , \7729 , RI9870c90_103);
and \U$23549 ( \23892 , RI9871230_115, \7727 );
nor \U$23550 ( \23893 , \23891 , \23892 );
and \U$23551 ( \23894 , \23893 , \7480 );
not \U$23552 ( \23895 , \23893 );
and \U$23553 ( \23896 , \23895 , \7733 );
nor \U$23554 ( \23897 , \23894 , \23896 );
and \U$23555 ( \23898 , \8486 , RI9871140_113);
and \U$23556 ( \23899 , RI9871320_117, \8484 );
nor \U$23557 ( \23900 , \23898 , \23899 );
and \U$23558 ( \23901 , \23900 , \8050 );
not \U$23559 ( \23902 , \23900 );
and \U$23560 ( \23903 , \23902 , \8051 );
nor \U$23561 ( \23904 , \23901 , \23903 );
xor \U$23562 ( \23905 , \23897 , \23904 );
and \U$23563 ( \23906 , \9237 , RI9871410_119);
and \U$23564 ( \23907 , RI98716e0_125, \9235 );
nor \U$23565 ( \23908 , \23906 , \23907 );
and \U$23566 ( \23909 , \23908 , \9241 );
not \U$23567 ( \23910 , \23908 );
and \U$23568 ( \23911 , \23910 , \8836 );
nor \U$23569 ( \23912 , \23909 , \23911 );
and \U$23570 ( \23913 , \23905 , \23912 );
and \U$23571 ( \23914 , \23897 , \23904 );
or \U$23572 ( \23915 , \23913 , \23914 );
and \U$23573 ( \23916 , \7079 , RI9870ba0_101);
and \U$23574 ( \23917 , RI9871050_111, \7077 );
nor \U$23575 ( \23918 , \23916 , \23917 );
and \U$23576 ( \23919 , \23918 , \6710 );
not \U$23577 ( \23920 , \23918 );
and \U$23578 ( \23921 , \23920 , \6709 );
nor \U$23579 ( \23922 , \23919 , \23921 );
and \U$23580 ( \23923 , \5881 , RI9870ab0_99);
and \U$23581 ( \23924 , RI9870d80_105, \5879 );
nor \U$23582 ( \23925 , \23923 , \23924 );
and \U$23583 ( \23926 , \23925 , \5594 );
not \U$23584 ( \23927 , \23925 );
and \U$23585 ( \23928 , \23927 , \5885 );
nor \U$23586 ( \23929 , \23926 , \23928 );
xor \U$23587 ( \23930 , \23922 , \23929 );
and \U$23588 ( \23931 , \6453 , RI98709c0_97);
and \U$23589 ( \23932 , RI9870e70_107, \6451 );
nor \U$23590 ( \23933 , \23931 , \23932 );
and \U$23591 ( \23934 , \23933 , \6190 );
not \U$23592 ( \23935 , \23933 );
and \U$23593 ( \23936 , \23935 , \6705 );
nor \U$23594 ( \23937 , \23934 , \23936 );
and \U$23595 ( \23938 , \23930 , \23937 );
and \U$23596 ( \23939 , \23922 , \23929 );
or \U$23597 ( \23940 , \23938 , \23939 );
xor \U$23598 ( \23941 , \23915 , \23940 );
and \U$23599 ( \23942 , \4203 , RI986fca0_69);
and \U$23600 ( \23943 , RI986ff70_75, \4201 );
nor \U$23601 ( \23944 , \23942 , \23943 );
and \U$23602 ( \23945 , \23944 , \4207 );
not \U$23603 ( \23946 , \23944 );
and \U$23604 ( \23947 , \23946 , \3922 );
nor \U$23605 ( \23948 , \23945 , \23947 );
not \U$23606 ( \23949 , \4521 );
and \U$23607 ( \23950 , \4710 , RI986fe80_73);
and \U$23608 ( \23951 , RI9870060_77, \4708 );
nor \U$23609 ( \23952 , \23950 , \23951 );
not \U$23610 ( \23953 , \23952 );
or \U$23611 ( \23954 , \23949 , \23953 );
or \U$23612 ( \23955 , \23952 , \4519 );
nand \U$23613 ( \23956 , \23954 , \23955 );
xor \U$23614 ( \23957 , \23948 , \23956 );
and \U$23615 ( \23958 , \5318 , RI9870150_79);
and \U$23616 ( \23959 , RI9870f60_109, \5316 );
nor \U$23617 ( \23960 , \23958 , \23959 );
and \U$23618 ( \23961 , \23960 , \5052 );
not \U$23619 ( \23962 , \23960 );
and \U$23620 ( \23963 , \23962 , \5322 );
nor \U$23621 ( \23964 , \23961 , \23963 );
and \U$23622 ( \23965 , \23957 , \23964 );
and \U$23623 ( \23966 , \23948 , \23956 );
or \U$23624 ( \23967 , \23965 , \23966 );
and \U$23625 ( \23968 , \23941 , \23967 );
and \U$23626 ( \23969 , \23915 , \23940 );
or \U$23627 ( \23970 , \23968 , \23969 );
and \U$23628 ( \23971 , \23890 , \23970 );
and \U$23629 ( \23972 , \23826 , \23889 );
or \U$23630 ( \23973 , \23971 , \23972 );
xor \U$23631 ( \23974 , \23753 , \23973 );
xor \U$23632 ( \23975 , \23627 , \23632 );
xor \U$23633 ( \23976 , \23975 , \23635 );
xor \U$23634 ( \23977 , \23413 , \23415 );
xor \U$23635 ( \23978 , \23977 , \23418 );
and \U$23636 ( \23979 , \23976 , \23978 );
xor \U$23637 ( \23980 , \23282 , \23289 );
xor \U$23638 ( \23981 , \23980 , \23297 );
xor \U$23639 ( \23982 , \23426 , \23431 );
xor \U$23640 ( \23983 , \23981 , \23982 );
xor \U$23641 ( \23984 , \23413 , \23415 );
xor \U$23642 ( \23985 , \23984 , \23418 );
and \U$23643 ( \23986 , \23983 , \23985 );
and \U$23644 ( \23987 , \23976 , \23983 );
or \U$23645 ( \23988 , \23979 , \23986 , \23987 );
and \U$23646 ( \23989 , \23974 , \23988 );
and \U$23647 ( \23990 , \23753 , \23973 );
or \U$23648 ( \23991 , \23989 , \23990 );
xor \U$23649 ( \23992 , \23520 , \23600 );
xor \U$23650 ( \23993 , \23992 , \23638 );
xor \U$23651 ( \23994 , \23421 , \23423 );
xor \U$23652 ( \23995 , \23994 , \23436 );
and \U$23653 ( \23996 , \23993 , \23995 );
xor \U$23654 ( \23997 , \23991 , \23996 );
xor \U$23655 ( \23998 , \23248 , \23274 );
xor \U$23656 ( \23999 , \23998 , \23300 );
not \U$23657 ( \24000 , \23167 );
xor \U$23658 ( \24001 , \23217 , \23193 );
not \U$23659 ( \24002 , \24001 );
or \U$23660 ( \24003 , \24000 , \24002 );
or \U$23661 ( \24004 , \24001 , \23167 );
nand \U$23662 ( \24005 , \24003 , \24004 );
xor \U$23663 ( \24006 , \23999 , \24005 );
xor \U$23664 ( \24007 , \23067 , \23069 );
xor \U$23665 ( \24008 , \24007 , \23072 );
xor \U$23666 ( \24009 , \23644 , \23651 );
xor \U$23667 ( \24010 , \24008 , \24009 );
and \U$23668 ( \24011 , \24006 , \24010 );
and \U$23669 ( \24012 , \23999 , \24005 );
or \U$23670 ( \24013 , \24011 , \24012 );
and \U$23671 ( \24014 , \23997 , \24013 );
and \U$23672 ( \24015 , \23991 , \23996 );
or \U$23673 ( \24016 , \24014 , \24015 );
xor \U$23674 ( \24017 , \23712 , \24016 );
xor \U$23675 ( \24018 , \23083 , \23305 );
xor \U$23676 ( \24019 , \24018 , \23320 );
xor \U$23677 ( \24020 , \23364 , \23371 );
xor \U$23678 ( \24021 , \24019 , \24020 );
and \U$23679 ( \24022 , \24017 , \24021 );
and \U$23680 ( \24023 , \23712 , \24016 );
or \U$23681 ( \24024 , \24022 , \24023 );
xor \U$23682 ( \24025 , \23697 , \24024 );
not \U$23683 ( \24026 , \23408 );
not \U$23684 ( \24027 , \23659 );
not \U$23685 ( \24028 , \23393 );
or \U$23686 ( \24029 , \24027 , \24028 );
or \U$23687 ( \24030 , \23393 , \23659 );
nand \U$23688 ( \24031 , \24029 , \24030 );
not \U$23689 ( \24032 , \24031 );
or \U$23690 ( \24033 , \24026 , \24032 );
or \U$23691 ( \24034 , \24031 , \23408 );
nand \U$23692 ( \24035 , \24033 , \24034 );
not \U$23693 ( \24036 , \24035 );
xor \U$23694 ( \24037 , \23712 , \24016 );
xor \U$23695 ( \24038 , \24037 , \24021 );
not \U$23696 ( \24039 , \24038 );
or \U$23697 ( \24040 , \24036 , \24039 );
or \U$23698 ( \24041 , \24038 , \24035 );
xor \U$23699 ( \24042 , \23786 , \1315 );
xor \U$23700 ( \24043 , \24042 , \23794 );
xor \U$23701 ( \24044 , \23760 , \23767 );
xor \U$23702 ( \24045 , \24044 , \23775 );
and \U$23703 ( \24046 , \24043 , \24045 );
xor \U$23704 ( \24047 , \23805 , \23812 );
xor \U$23705 ( \24048 , \24047 , \23820 );
xor \U$23706 ( \24049 , \23760 , \23767 );
xor \U$23707 ( \24050 , \24049 , \23775 );
and \U$23708 ( \24051 , \24048 , \24050 );
and \U$23709 ( \24052 , \24043 , \24048 );
or \U$23710 ( \24053 , \24046 , \24051 , \24052 );
xor \U$23711 ( \24054 , \23527 , \23534 );
xor \U$23712 ( \24055 , \24054 , \23542 );
xor \U$23713 ( \24056 , \24053 , \24055 );
xor \U$23714 ( \24057 , \23948 , \23956 );
xor \U$23715 ( \24058 , \24057 , \23964 );
xor \U$23716 ( \24059 , \23922 , \23929 );
xor \U$23717 ( \24060 , \24059 , \23937 );
xor \U$23718 ( \24061 , \24058 , \24060 );
xor \U$23719 ( \24062 , \23897 , \23904 );
xor \U$23720 ( \24063 , \24062 , \23912 );
and \U$23721 ( \24064 , \24061 , \24063 );
and \U$23722 ( \24065 , \24058 , \24060 );
or \U$23723 ( \24066 , \24064 , \24065 );
and \U$23724 ( \24067 , \24056 , \24066 );
and \U$23725 ( \24068 , \24053 , \24055 );
or \U$23726 ( \24069 , \24067 , \24068 );
and \U$23727 ( \24070 , \5318 , RI9870060_77);
and \U$23728 ( \24071 , RI9870150_79, \5316 );
nor \U$23729 ( \24072 , \24070 , \24071 );
and \U$23730 ( \24073 , \24072 , \5052 );
not \U$23731 ( \24074 , \24072 );
and \U$23732 ( \24075 , \24074 , \5322 );
nor \U$23733 ( \24076 , \24073 , \24075 );
and \U$23734 ( \24077 , \5881 , RI9870f60_109);
and \U$23735 ( \24078 , RI9870ab0_99, \5879 );
nor \U$23736 ( \24079 , \24077 , \24078 );
and \U$23737 ( \24080 , \24079 , \5594 );
not \U$23738 ( \24081 , \24079 );
and \U$23739 ( \24082 , \24081 , \5885 );
nor \U$23740 ( \24083 , \24080 , \24082 );
xor \U$23741 ( \24084 , \24076 , \24083 );
and \U$23742 ( \24085 , \6453 , RI9870d80_105);
and \U$23743 ( \24086 , RI98709c0_97, \6451 );
nor \U$23744 ( \24087 , \24085 , \24086 );
and \U$23745 ( \24088 , \24087 , \6190 );
not \U$23746 ( \24089 , \24087 );
and \U$23747 ( \24090 , \24089 , \6180 );
nor \U$23748 ( \24091 , \24088 , \24090 );
and \U$23749 ( \24092 , \24084 , \24091 );
and \U$23750 ( \24093 , \24076 , \24083 );
or \U$23751 ( \24094 , \24092 , \24093 );
not \U$23752 ( \24095 , \3412 );
and \U$23753 ( \24096 , \3683 , RI986fac0_65);
and \U$23754 ( \24097 , RI986fbb0_67, \3681 );
nor \U$23755 ( \24098 , \24096 , \24097 );
not \U$23756 ( \24099 , \24098 );
or \U$23757 ( \24100 , \24095 , \24099 );
or \U$23758 ( \24101 , \24098 , \3918 );
nand \U$23759 ( \24102 , \24100 , \24101 );
and \U$23760 ( \24103 , \4203 , RI986fd90_71);
and \U$23761 ( \24104 , RI986fca0_69, \4201 );
nor \U$23762 ( \24105 , \24103 , \24104 );
and \U$23763 ( \24106 , \24105 , \4207 );
not \U$23764 ( \24107 , \24105 );
and \U$23765 ( \24108 , \24107 , \3922 );
nor \U$23766 ( \24109 , \24106 , \24108 );
xor \U$23767 ( \24110 , \24102 , \24109 );
not \U$23768 ( \24111 , \4519 );
and \U$23769 ( \24112 , \4710 , RI986ff70_75);
and \U$23770 ( \24113 , RI986fe80_73, \4708 );
nor \U$23771 ( \24114 , \24112 , \24113 );
not \U$23772 ( \24115 , \24114 );
or \U$23773 ( \24116 , \24111 , \24115 );
or \U$23774 ( \24117 , \24114 , \4521 );
nand \U$23775 ( \24118 , \24116 , \24117 );
and \U$23776 ( \24119 , \24110 , \24118 );
and \U$23777 ( \24120 , \24102 , \24109 );
or \U$23778 ( \24121 , \24119 , \24120 );
xor \U$23779 ( \24122 , \24094 , \24121 );
and \U$23780 ( \24123 , \7079 , RI9870e70_107);
and \U$23781 ( \24124 , RI9870ba0_101, \7077 );
nor \U$23782 ( \24125 , \24123 , \24124 );
and \U$23783 ( \24126 , \24125 , \6710 );
not \U$23784 ( \24127 , \24125 );
and \U$23785 ( \24128 , \24127 , \6709 );
nor \U$23786 ( \24129 , \24126 , \24128 );
and \U$23787 ( \24130 , \7729 , RI9871050_111);
and \U$23788 ( \24131 , RI9870c90_103, \7727 );
nor \U$23789 ( \24132 , \24130 , \24131 );
and \U$23790 ( \24133 , \24132 , \7480 );
not \U$23791 ( \24134 , \24132 );
and \U$23792 ( \24135 , \24134 , \7733 );
nor \U$23793 ( \24136 , \24133 , \24135 );
xor \U$23794 ( \24137 , \24129 , \24136 );
and \U$23795 ( \24138 , \8486 , RI9871230_115);
and \U$23796 ( \24139 , RI9871140_113, \8484 );
nor \U$23797 ( \24140 , \24138 , \24139 );
and \U$23798 ( \24141 , \24140 , \8050 );
not \U$23799 ( \24142 , \24140 );
and \U$23800 ( \24143 , \24142 , \8051 );
nor \U$23801 ( \24144 , \24141 , \24143 );
and \U$23802 ( \24145 , \24137 , \24144 );
and \U$23803 ( \24146 , \24129 , \24136 );
or \U$23804 ( \24147 , \24145 , \24146 );
and \U$23805 ( \24148 , \24122 , \24147 );
and \U$23806 ( \24149 , \24094 , \24121 );
or \U$23807 ( \24150 , \24148 , \24149 );
and \U$23808 ( \24151 , \11696 , RI986ead0_31);
and \U$23809 ( \24152 , RI986e9e0_29, \11694 );
nor \U$23810 ( \24153 , \24151 , \24152 );
and \U$23811 ( \24154 , \24153 , \10965 );
not \U$23812 ( \24155 , \24153 );
and \U$23813 ( \24156 , \24155 , \11702 );
nor \U$23814 ( \24157 , \24154 , \24156 );
and \U$23815 ( \24158 , \12293 , RI986e8f0_27);
and \U$23816 ( \24159 , RI986e800_25, \12291 );
nor \U$23817 ( \24160 , \24158 , \24159 );
and \U$23818 ( \24161 , \24160 , \11687 );
not \U$23819 ( \24162 , \24160 );
and \U$23820 ( \24163 , \24162 , \11686 );
nor \U$23821 ( \24164 , \24161 , \24163 );
xor \U$23822 ( \24165 , \24157 , \24164 );
and \U$23823 ( \24166 , \13045 , RI986ee90_39);
and \U$23824 ( \24167 , RI986eda0_37, \13043 );
nor \U$23825 ( \24168 , \24166 , \24167 );
and \U$23826 ( \24169 , \24168 , \13047 );
not \U$23827 ( \24170 , \24168 );
and \U$23828 ( \24171 , \24170 , \12619 );
nor \U$23829 ( \24172 , \24169 , \24171 );
and \U$23830 ( \24173 , \24165 , \24172 );
and \U$23831 ( \24174 , \24157 , \24164 );
or \U$23832 ( \24175 , \24173 , \24174 );
and \U$23833 ( \24176 , \13882 , RI986ebc0_33);
and \U$23834 ( \24177 , RI986ecb0_35, \13880 );
nor \U$23835 ( \24178 , \24176 , \24177 );
and \U$23836 ( \24179 , \24178 , \13358 );
not \U$23837 ( \24180 , \24178 );
and \U$23838 ( \24181 , \24180 , \13359 );
nor \U$23839 ( \24182 , \24179 , \24181 );
not \U$23840 ( \24183 , RI9873558_190);
and \U$23841 ( \24184 , \15780 , RI986f250_47);
and \U$23842 ( \24185 , RI9873648_192, RI986f160_45);
nor \U$23843 ( \24186 , \24184 , \24185 );
not \U$23844 ( \24187 , \24186 );
or \U$23845 ( \24188 , \24183 , \24187 );
or \U$23846 ( \24189 , \24186 , RI9873558_190);
nand \U$23847 ( \24190 , \24188 , \24189 );
xor \U$23848 ( \24191 , \24182 , \24190 );
and \U$23849 ( \24192 , \14937 , RI986f070_43);
and \U$23850 ( \24193 , RI986ef80_41, \14935 );
nor \U$23851 ( \24194 , \24192 , \24193 );
and \U$23852 ( \24195 , \24194 , \14539 );
not \U$23853 ( \24196 , \24194 );
and \U$23854 ( \24197 , \24196 , \14538 );
nor \U$23855 ( \24198 , \24195 , \24197 );
and \U$23856 ( \24199 , \24191 , \24198 );
and \U$23857 ( \24200 , \24182 , \24190 );
or \U$23858 ( \24201 , \24199 , \24200 );
xor \U$23859 ( \24202 , \24175 , \24201 );
and \U$23860 ( \24203 , \10424 , RI9871500_121);
and \U$23861 ( \24204 , RI98715f0_123, \10422 );
nor \U$23862 ( \24205 , \24203 , \24204 );
and \U$23863 ( \24206 , \24205 , \9840 );
not \U$23864 ( \24207 , \24205 );
and \U$23865 ( \24208 , \24207 , \10428 );
nor \U$23866 ( \24209 , \24206 , \24208 );
and \U$23867 ( \24210 , \9237 , RI9871320_117);
and \U$23868 ( \24211 , RI9871410_119, \9235 );
nor \U$23869 ( \24212 , \24210 , \24211 );
and \U$23870 ( \24213 , \24212 , \9241 );
not \U$23871 ( \24214 , \24212 );
and \U$23872 ( \24215 , \24214 , \8836 );
nor \U$23873 ( \24216 , \24213 , \24215 );
xor \U$23874 ( \24217 , \24209 , \24216 );
and \U$23875 ( \24218 , \9505 , RI98716e0_125);
and \U$23876 ( \24219 , RI98717d0_127, \9503 );
nor \U$23877 ( \24220 , \24218 , \24219 );
and \U$23878 ( \24221 , \24220 , \9510 );
not \U$23879 ( \24222 , \24220 );
and \U$23880 ( \24223 , \24222 , \9513 );
nor \U$23881 ( \24224 , \24221 , \24223 );
and \U$23882 ( \24225 , \24217 , \24224 );
and \U$23883 ( \24226 , \24209 , \24216 );
or \U$23884 ( \24227 , \24225 , \24226 );
and \U$23885 ( \24228 , \24202 , \24227 );
and \U$23886 ( \24229 , \24175 , \24201 );
or \U$23887 ( \24230 , \24228 , \24229 );
xor \U$23888 ( \24231 , \24150 , \24230 );
and \U$23889 ( \24232 , \2274 , RI9870330_83);
and \U$23890 ( \24233 , RI9870240_81, \2272 );
nor \U$23891 ( \24234 , \24232 , \24233 );
and \U$23892 ( \24235 , \24234 , \2030 );
not \U$23893 ( \24236 , \24234 );
and \U$23894 ( \24237 , \24236 , \2031 );
nor \U$23895 ( \24238 , \24235 , \24237 );
and \U$23896 ( \24239 , \2464 , RI98706f0_91);
and \U$23897 ( \24240 , RI9870600_89, \2462 );
nor \U$23898 ( \24241 , \24239 , \24240 );
and \U$23899 ( \24242 , \24241 , \2468 );
not \U$23900 ( \24243 , \24241 );
and \U$23901 ( \24244 , \24243 , \2263 );
nor \U$23902 ( \24245 , \24242 , \24244 );
xor \U$23903 ( \24246 , \24238 , \24245 );
not \U$23904 ( \24247 , \3406 );
and \U$23905 ( \24248 , \3254 , RI98708d0_95);
and \U$23906 ( \24249 , RI98707e0_93, \3252 );
nor \U$23907 ( \24250 , \24248 , \24249 );
not \U$23908 ( \24251 , \24250 );
or \U$23909 ( \24252 , \24247 , \24251 );
or \U$23910 ( \24253 , \24250 , \2935 );
nand \U$23911 ( \24254 , \24252 , \24253 );
and \U$23912 ( \24255 , \24246 , \24254 );
and \U$23913 ( \24256 , \24238 , \24245 );
or \U$23914 ( \24257 , \24255 , \24256 );
xor \U$23915 ( \24258 , \23833 , \23838 );
xor \U$23916 ( \24259 , \24258 , \23847 );
and \U$23917 ( \24260 , \24257 , \24259 );
xor \U$23918 ( \24261 , \23866 , \23874 );
xor \U$23919 ( \24262 , \24261 , \23883 );
xor \U$23920 ( \24263 , \23833 , \23838 );
xor \U$23921 ( \24264 , \24263 , \23847 );
and \U$23922 ( \24265 , \24262 , \24264 );
and \U$23923 ( \24266 , \24257 , \24262 );
or \U$23924 ( \24267 , \24260 , \24265 , \24266 );
and \U$23925 ( \24268 , \24231 , \24267 );
and \U$23926 ( \24269 , \24150 , \24230 );
or \U$23927 ( \24270 , \24268 , \24269 );
xor \U$23928 ( \24271 , \24069 , \24270 );
xor \U$23929 ( \24272 , \23552 , \23560 );
xor \U$23930 ( \24273 , \24272 , \23568 );
xor \U$23931 ( \24274 , \23714 , \23721 );
xor \U$23932 ( \24275 , \24274 , \23724 );
and \U$23933 ( \24276 , \24273 , \24275 );
xor \U$23934 ( \24277 , \23446 , \23453 );
xor \U$23935 ( \24278 , \24277 , \23461 );
xor \U$23936 ( \24279 , \23740 , \23745 );
xor \U$23937 ( \24280 , \24278 , \24279 );
xor \U$23938 ( \24281 , \23714 , \23721 );
xor \U$23939 ( \24282 , \24281 , \23724 );
and \U$23940 ( \24283 , \24280 , \24282 );
and \U$23941 ( \24284 , \24273 , \24280 );
or \U$23942 ( \24285 , \24276 , \24283 , \24284 );
and \U$23943 ( \24286 , \24271 , \24285 );
and \U$23944 ( \24287 , \24069 , \24270 );
or \U$23945 ( \24288 , \24286 , \24287 );
xor \U$23946 ( \24289 , \23545 , \23571 );
xor \U$23947 ( \24290 , \24289 , \23597 );
xor \U$23948 ( \24291 , \23464 , \23491 );
xor \U$23949 ( \24292 , \24291 , \23517 );
and \U$23950 ( \24293 , \24290 , \24292 );
xor \U$23951 ( \24294 , \23915 , \23940 );
xor \U$23952 ( \24295 , \24294 , \23967 );
xor \U$23953 ( \24296 , \23778 , \23797 );
xor \U$23954 ( \24297 , \24296 , \23823 );
xor \U$23955 ( \24298 , \24295 , \24297 );
xor \U$23956 ( \24299 , \23850 , \23858 );
xor \U$23957 ( \24300 , \24299 , \23886 );
and \U$23958 ( \24301 , \24298 , \24300 );
and \U$23959 ( \24302 , \24295 , \24297 );
or \U$23960 ( \24303 , \24301 , \24302 );
xor \U$23961 ( \24304 , \23464 , \23491 );
xor \U$23962 ( \24305 , \24304 , \23517 );
and \U$23963 ( \24306 , \24303 , \24305 );
and \U$23964 ( \24307 , \24290 , \24303 );
or \U$23965 ( \24308 , \24293 , \24306 , \24307 );
xor \U$23966 ( \24309 , \24288 , \24308 );
xor \U$23967 ( \24310 , \23826 , \23889 );
xor \U$23968 ( \24311 , \24310 , \23970 );
xor \U$23969 ( \24312 , \23727 , \23737 );
xor \U$23970 ( \24313 , \24312 , \23750 );
and \U$23971 ( \24314 , \24311 , \24313 );
xor \U$23972 ( \24315 , \23413 , \23415 );
xor \U$23973 ( \24316 , \24315 , \23418 );
xor \U$23974 ( \24317 , \23976 , \23983 );
xor \U$23975 ( \24318 , \24316 , \24317 );
xor \U$23976 ( \24319 , \23727 , \23737 );
xor \U$23977 ( \24320 , \24319 , \23750 );
and \U$23978 ( \24321 , \24318 , \24320 );
and \U$23979 ( \24322 , \24311 , \24318 );
or \U$23980 ( \24323 , \24314 , \24321 , \24322 );
and \U$23981 ( \24324 , \24309 , \24323 );
and \U$23982 ( \24325 , \24288 , \24308 );
or \U$23983 ( \24326 , \24324 , \24325 );
xor \U$23984 ( \24327 , \23993 , \23995 );
xor \U$23985 ( \24328 , \23999 , \24005 );
xor \U$23986 ( \24329 , \24328 , \24010 );
and \U$23987 ( \24330 , \24327 , \24329 );
xor \U$23988 ( \24331 , \23753 , \23973 );
xor \U$23989 ( \24332 , \24331 , \23988 );
xor \U$23990 ( \24333 , \23999 , \24005 );
xor \U$23991 ( \24334 , \24333 , \24010 );
and \U$23992 ( \24335 , \24332 , \24334 );
and \U$23993 ( \24336 , \24327 , \24332 );
or \U$23994 ( \24337 , \24330 , \24335 , \24336 );
xor \U$23995 ( \24338 , \24326 , \24337 );
xor \U$23996 ( \24339 , \23382 , \23384 );
xor \U$23997 ( \24340 , \24339 , \23389 );
xor \U$23998 ( \24341 , \23702 , \23707 );
xor \U$23999 ( \24342 , \24340 , \24341 );
and \U$24000 ( \24343 , \24338 , \24342 );
and \U$24001 ( \24344 , \24326 , \24337 );
or \U$24002 ( \24345 , \24343 , \24344 );
nand \U$24003 ( \24346 , \24041 , \24345 );
nand \U$24004 ( \24347 , \24040 , \24346 );
and \U$24005 ( \24348 , \24025 , \24347 );
xor \U$24006 ( \24349 , \24347 , \24025 );
xor \U$24007 ( \24350 , \24069 , \24270 );
xor \U$24008 ( \24351 , \24350 , \24285 );
xor \U$24009 ( \24352 , \24053 , \24055 );
xor \U$24010 ( \24353 , \24352 , \24066 );
xor \U$24011 ( \24354 , \24295 , \24297 );
xor \U$24012 ( \24355 , \24354 , \24300 );
and \U$24013 ( \24356 , \24353 , \24355 );
xor \U$24014 ( \24357 , \23714 , \23721 );
xor \U$24015 ( \24358 , \24357 , \23724 );
xor \U$24016 ( \24359 , \24273 , \24280 );
xor \U$24017 ( \24360 , \24358 , \24359 );
xor \U$24018 ( \24361 , \24295 , \24297 );
xor \U$24019 ( \24362 , \24361 , \24300 );
and \U$24020 ( \24363 , \24360 , \24362 );
and \U$24021 ( \24364 , \24353 , \24360 );
or \U$24022 ( \24365 , \24356 , \24363 , \24364 );
xor \U$24023 ( \24366 , \24094 , \24121 );
xor \U$24024 ( \24367 , \24366 , \24147 );
xor \U$24025 ( \24368 , \24058 , \24060 );
xor \U$24026 ( \24369 , \24368 , \24063 );
and \U$24027 ( \24370 , \24367 , \24369 );
xor \U$24028 ( \24371 , \23833 , \23838 );
xor \U$24029 ( \24372 , \24371 , \23847 );
xor \U$24030 ( \24373 , \24257 , \24262 );
xor \U$24031 ( \24374 , \24372 , \24373 );
xor \U$24032 ( \24375 , \24058 , \24060 );
xor \U$24033 ( \24376 , \24375 , \24063 );
and \U$24034 ( \24377 , \24374 , \24376 );
and \U$24035 ( \24378 , \24367 , \24374 );
or \U$24036 ( \24379 , \24370 , \24377 , \24378 );
and \U$24037 ( \24380 , \12293 , RI986e9e0_29);
and \U$24038 ( \24381 , RI986e8f0_27, \12291 );
nor \U$24039 ( \24382 , \24380 , \24381 );
and \U$24040 ( \24383 , \24382 , \11687 );
not \U$24041 ( \24384 , \24382 );
and \U$24042 ( \24385 , \24384 , \11686 );
nor \U$24043 ( \24386 , \24383 , \24385 );
and \U$24044 ( \24387 , \13045 , RI986e800_25);
and \U$24045 ( \24388 , RI986ee90_39, \13043 );
nor \U$24046 ( \24389 , \24387 , \24388 );
and \U$24047 ( \24390 , \24389 , \13047 );
not \U$24048 ( \24391 , \24389 );
and \U$24049 ( \24392 , \24391 , \12619 );
nor \U$24050 ( \24393 , \24390 , \24392 );
xor \U$24051 ( \24394 , \24386 , \24393 );
and \U$24052 ( \24395 , \13882 , RI986eda0_37);
and \U$24053 ( \24396 , RI986ebc0_33, \13880 );
nor \U$24054 ( \24397 , \24395 , \24396 );
and \U$24055 ( \24398 , \24397 , \13358 );
not \U$24056 ( \24399 , \24397 );
and \U$24057 ( \24400 , \24399 , \13359 );
nor \U$24058 ( \24401 , \24398 , \24400 );
and \U$24059 ( \24402 , \24394 , \24401 );
and \U$24060 ( \24403 , \24386 , \24393 );
or \U$24061 ( \24404 , \24402 , \24403 );
not \U$24062 ( \24405 , RI9873558_190);
and \U$24063 ( \24406 , \15780 , RI986ef80_41);
and \U$24064 ( \24407 , RI9873648_192, RI986f250_47);
nor \U$24065 ( \24408 , \24406 , \24407 );
not \U$24066 ( \24409 , \24408 );
or \U$24067 ( \24410 , \24405 , \24409 );
or \U$24068 ( \24411 , \24408 , RI9873558_190);
nand \U$24069 ( \24412 , \24410 , \24411 );
xor \U$24070 ( \24413 , \24412 , \2034 );
and \U$24071 ( \24414 , \14937 , RI986ecb0_35);
and \U$24072 ( \24415 , RI986f070_43, \14935 );
nor \U$24073 ( \24416 , \24414 , \24415 );
and \U$24074 ( \24417 , \24416 , \14539 );
not \U$24075 ( \24418 , \24416 );
and \U$24076 ( \24419 , \24418 , \14538 );
nor \U$24077 ( \24420 , \24417 , \24419 );
and \U$24078 ( \24421 , \24413 , \24420 );
and \U$24079 ( \24422 , \24412 , \2034 );
or \U$24080 ( \24423 , \24421 , \24422 );
xor \U$24081 ( \24424 , \24404 , \24423 );
and \U$24082 ( \24425 , \9505 , RI9871410_119);
and \U$24083 ( \24426 , RI98716e0_125, \9503 );
nor \U$24084 ( \24427 , \24425 , \24426 );
and \U$24085 ( \24428 , \24427 , \9510 );
not \U$24086 ( \24429 , \24427 );
and \U$24087 ( \24430 , \24429 , \9513 );
nor \U$24088 ( \24431 , \24428 , \24430 );
and \U$24089 ( \24432 , \10424 , RI98717d0_127);
and \U$24090 ( \24433 , RI9871500_121, \10422 );
nor \U$24091 ( \24434 , \24432 , \24433 );
and \U$24092 ( \24435 , \24434 , \9840 );
not \U$24093 ( \24436 , \24434 );
and \U$24094 ( \24437 , \24436 , \10428 );
nor \U$24095 ( \24438 , \24435 , \24437 );
xor \U$24096 ( \24439 , \24431 , \24438 );
and \U$24097 ( \24440 , \11696 , RI98715f0_123);
and \U$24098 ( \24441 , RI986ead0_31, \11694 );
nor \U$24099 ( \24442 , \24440 , \24441 );
and \U$24100 ( \24443 , \24442 , \10965 );
not \U$24101 ( \24444 , \24442 );
and \U$24102 ( \24445 , \24444 , \11702 );
nor \U$24103 ( \24446 , \24443 , \24445 );
and \U$24104 ( \24447 , \24439 , \24446 );
and \U$24105 ( \24448 , \24431 , \24438 );
or \U$24106 ( \24449 , \24447 , \24448 );
and \U$24107 ( \24450 , \24424 , \24449 );
and \U$24108 ( \24451 , \24404 , \24423 );
or \U$24109 ( \24452 , \24450 , \24451 );
nand \U$24110 ( \24453 , RI9870420_85, \2040 );
not \U$24111 ( \24454 , \24453 );
not \U$24112 ( \24455 , \2034 );
or \U$24113 ( \24456 , \24454 , \24455 );
or \U$24114 ( \24457 , \1462 , \24453 );
nand \U$24115 ( \24458 , \24456 , \24457 );
and \U$24116 ( \24459 , \2274 , RI9870510_87);
and \U$24117 ( \24460 , RI9870330_83, \2272 );
nor \U$24118 ( \24461 , \24459 , \24460 );
and \U$24119 ( \24462 , \24461 , \2030 );
not \U$24120 ( \24463 , \24461 );
and \U$24121 ( \24464 , \24463 , \2031 );
nor \U$24122 ( \24465 , \24462 , \24464 );
and \U$24123 ( \24466 , \24458 , \24465 );
not \U$24124 ( \24467 , \1462 );
and \U$24125 ( \24468 , \2042 , RI9870420_85);
and \U$24126 ( \24469 , RI9870510_87, \2040 );
nor \U$24127 ( \24470 , \24468 , \24469 );
not \U$24128 ( \24471 , \24470 );
or \U$24129 ( \24472 , \24467 , \24471 );
or \U$24130 ( \24473 , \24470 , \2034 );
nand \U$24131 ( \24474 , \24472 , \24473 );
xor \U$24132 ( \24475 , \24466 , \24474 );
and \U$24133 ( \24476 , \2464 , RI9870240_81);
and \U$24134 ( \24477 , RI98706f0_91, \2462 );
nor \U$24135 ( \24478 , \24476 , \24477 );
and \U$24136 ( \24479 , \24478 , \2468 );
not \U$24137 ( \24480 , \24478 );
and \U$24138 ( \24481 , \24480 , \2263 );
nor \U$24139 ( \24482 , \24479 , \24481 );
not \U$24140 ( \24483 , \2935 );
and \U$24141 ( \24484 , \3254 , RI9870600_89);
and \U$24142 ( \24485 , RI98708d0_95, \3252 );
nor \U$24143 ( \24486 , \24484 , \24485 );
not \U$24144 ( \24487 , \24486 );
or \U$24145 ( \24488 , \24483 , \24487 );
or \U$24146 ( \24489 , \24486 , \2935 );
nand \U$24147 ( \24490 , \24488 , \24489 );
xor \U$24148 ( \24491 , \24482 , \24490 );
not \U$24149 ( \24492 , \3412 );
and \U$24150 ( \24493 , \3683 , RI98707e0_93);
and \U$24151 ( \24494 , RI986fac0_65, \3681 );
nor \U$24152 ( \24495 , \24493 , \24494 );
not \U$24153 ( \24496 , \24495 );
or \U$24154 ( \24497 , \24492 , \24496 );
or \U$24155 ( \24498 , \24495 , \3918 );
nand \U$24156 ( \24499 , \24497 , \24498 );
and \U$24157 ( \24500 , \24491 , \24499 );
and \U$24158 ( \24501 , \24482 , \24490 );
or \U$24159 ( \24502 , \24500 , \24501 );
and \U$24160 ( \24503 , \24475 , \24502 );
and \U$24161 ( \24504 , \24466 , \24474 );
or \U$24162 ( \24505 , \24503 , \24504 );
xor \U$24163 ( \24506 , \24452 , \24505 );
and \U$24164 ( \24507 , \7729 , RI9870ba0_101);
and \U$24165 ( \24508 , RI9871050_111, \7727 );
nor \U$24166 ( \24509 , \24507 , \24508 );
and \U$24167 ( \24510 , \24509 , \7480 );
not \U$24168 ( \24511 , \24509 );
and \U$24169 ( \24512 , \24511 , \7733 );
nor \U$24170 ( \24513 , \24510 , \24512 );
and \U$24171 ( \24514 , \8486 , RI9870c90_103);
and \U$24172 ( \24515 , RI9871230_115, \8484 );
nor \U$24173 ( \24516 , \24514 , \24515 );
and \U$24174 ( \24517 , \24516 , \8050 );
not \U$24175 ( \24518 , \24516 );
and \U$24176 ( \24519 , \24518 , \8051 );
nor \U$24177 ( \24520 , \24517 , \24519 );
xor \U$24178 ( \24521 , \24513 , \24520 );
and \U$24179 ( \24522 , \9237 , RI9871140_113);
and \U$24180 ( \24523 , RI9871320_117, \9235 );
nor \U$24181 ( \24524 , \24522 , \24523 );
and \U$24182 ( \24525 , \24524 , \9241 );
not \U$24183 ( \24526 , \24524 );
and \U$24184 ( \24527 , \24526 , \8836 );
nor \U$24185 ( \24528 , \24525 , \24527 );
and \U$24186 ( \24529 , \24521 , \24528 );
and \U$24187 ( \24530 , \24513 , \24520 );
or \U$24188 ( \24531 , \24529 , \24530 );
and \U$24189 ( \24532 , \5318 , RI986fe80_73);
and \U$24190 ( \24533 , RI9870060_77, \5316 );
nor \U$24191 ( \24534 , \24532 , \24533 );
and \U$24192 ( \24535 , \24534 , \5052 );
not \U$24193 ( \24536 , \24534 );
and \U$24194 ( \24537 , \24536 , \5322 );
nor \U$24195 ( \24538 , \24535 , \24537 );
and \U$24196 ( \24539 , \4203 , RI986fbb0_67);
and \U$24197 ( \24540 , RI986fd90_71, \4201 );
nor \U$24198 ( \24541 , \24539 , \24540 );
and \U$24199 ( \24542 , \24541 , \4207 );
not \U$24200 ( \24543 , \24541 );
and \U$24201 ( \24544 , \24543 , \3922 );
nor \U$24202 ( \24545 , \24542 , \24544 );
xor \U$24203 ( \24546 , \24538 , \24545 );
not \U$24204 ( \24547 , \4519 );
and \U$24205 ( \24548 , \4710 , RI986fca0_69);
and \U$24206 ( \24549 , RI986ff70_75, \4708 );
nor \U$24207 ( \24550 , \24548 , \24549 );
not \U$24208 ( \24551 , \24550 );
or \U$24209 ( \24552 , \24547 , \24551 );
or \U$24210 ( \24553 , \24550 , \4519 );
nand \U$24211 ( \24554 , \24552 , \24553 );
and \U$24212 ( \24555 , \24546 , \24554 );
and \U$24213 ( \24556 , \24538 , \24545 );
or \U$24214 ( \24557 , \24555 , \24556 );
xor \U$24215 ( \24558 , \24531 , \24557 );
and \U$24216 ( \24559 , \5881 , RI9870150_79);
and \U$24217 ( \24560 , RI9870f60_109, \5879 );
nor \U$24218 ( \24561 , \24559 , \24560 );
and \U$24219 ( \24562 , \24561 , \5594 );
not \U$24220 ( \24563 , \24561 );
and \U$24221 ( \24564 , \24563 , \5885 );
nor \U$24222 ( \24565 , \24562 , \24564 );
and \U$24223 ( \24566 , \6453 , RI9870ab0_99);
and \U$24224 ( \24567 , RI9870d80_105, \6451 );
nor \U$24225 ( \24568 , \24566 , \24567 );
and \U$24226 ( \24569 , \24568 , \6190 );
not \U$24227 ( \24570 , \24568 );
and \U$24228 ( \24571 , \24570 , \6705 );
nor \U$24229 ( \24572 , \24569 , \24571 );
xor \U$24230 ( \24573 , \24565 , \24572 );
and \U$24231 ( \24574 , \7079 , RI98709c0_97);
and \U$24232 ( \24575 , RI9870e70_107, \7077 );
nor \U$24233 ( \24576 , \24574 , \24575 );
and \U$24234 ( \24577 , \24576 , \6710 );
not \U$24235 ( \24578 , \24576 );
and \U$24236 ( \24579 , \24578 , \6709 );
nor \U$24237 ( \24580 , \24577 , \24579 );
and \U$24238 ( \24581 , \24573 , \24580 );
and \U$24239 ( \24582 , \24565 , \24572 );
or \U$24240 ( \24583 , \24581 , \24582 );
and \U$24241 ( \24584 , \24558 , \24583 );
and \U$24242 ( \24585 , \24531 , \24557 );
or \U$24243 ( \24586 , \24584 , \24585 );
and \U$24244 ( \24587 , \24506 , \24586 );
and \U$24245 ( \24588 , \24452 , \24505 );
or \U$24246 ( \24589 , \24587 , \24588 );
xor \U$24247 ( \24590 , \24379 , \24589 );
xor \U$24248 ( \24591 , \24209 , \24216 );
xor \U$24249 ( \24592 , \24591 , \24224 );
xor \U$24250 ( \24593 , \24129 , \24136 );
xor \U$24251 ( \24594 , \24593 , \24144 );
and \U$24252 ( \24595 , \24592 , \24594 );
xor \U$24253 ( \24596 , \24157 , \24164 );
xor \U$24254 ( \24597 , \24596 , \24172 );
xor \U$24255 ( \24598 , \24129 , \24136 );
xor \U$24256 ( \24599 , \24598 , \24144 );
and \U$24257 ( \24600 , \24597 , \24599 );
and \U$24258 ( \24601 , \24592 , \24597 );
or \U$24259 ( \24602 , \24595 , \24600 , \24601 );
xor \U$24260 ( \24603 , \24238 , \24245 );
xor \U$24261 ( \24604 , \24603 , \24254 );
xor \U$24262 ( \24605 , \24102 , \24109 );
xor \U$24263 ( \24606 , \24605 , \24118 );
xor \U$24264 ( \24607 , \24604 , \24606 );
xor \U$24265 ( \24608 , \24076 , \24083 );
xor \U$24266 ( \24609 , \24608 , \24091 );
and \U$24267 ( \24610 , \24607 , \24609 );
and \U$24268 ( \24611 , \24604 , \24606 );
or \U$24269 ( \24612 , \24610 , \24611 );
xor \U$24270 ( \24613 , \24602 , \24612 );
xor \U$24271 ( \24614 , \23760 , \23767 );
xor \U$24272 ( \24615 , \24614 , \23775 );
xor \U$24273 ( \24616 , \24043 , \24048 );
xor \U$24274 ( \24617 , \24615 , \24616 );
and \U$24275 ( \24618 , \24613 , \24617 );
and \U$24276 ( \24619 , \24602 , \24612 );
or \U$24277 ( \24620 , \24618 , \24619 );
and \U$24278 ( \24621 , \24590 , \24620 );
and \U$24279 ( \24622 , \24379 , \24589 );
or \U$24280 ( \24623 , \24621 , \24622 );
xor \U$24281 ( \24624 , \24365 , \24623 );
xor \U$24282 ( \24625 , \23727 , \23737 );
xor \U$24283 ( \24626 , \24625 , \23750 );
xor \U$24284 ( \24627 , \24311 , \24318 );
xor \U$24285 ( \24628 , \24626 , \24627 );
xor \U$24286 ( \24629 , \24624 , \24628 );
and \U$24287 ( \24630 , \24351 , \24629 );
not \U$24288 ( \24631 , \24630 );
xor \U$24289 ( \24632 , \24365 , \24623 );
and \U$24290 ( \24633 , \24632 , \24628 );
and \U$24291 ( \24634 , \24365 , \24623 );
or \U$24292 ( \24635 , \24633 , \24634 );
xor \U$24293 ( \24636 , \24288 , \24308 );
xor \U$24294 ( \24637 , \24636 , \24323 );
xor \U$24295 ( \24638 , \24635 , \24637 );
xor \U$24296 ( \24639 , \23999 , \24005 );
xor \U$24297 ( \24640 , \24639 , \24010 );
xor \U$24298 ( \24641 , \24327 , \24332 );
xor \U$24299 ( \24642 , \24640 , \24641 );
xor \U$24300 ( \24643 , \24638 , \24642 );
not \U$24301 ( \24644 , \24643 );
or \U$24302 ( \24645 , \24631 , \24644 );
or \U$24303 ( \24646 , \24643 , \24630 );
xor \U$24304 ( \24647 , \24379 , \24589 );
xor \U$24305 ( \24648 , \24647 , \24620 );
xor \U$24306 ( \24649 , \24295 , \24297 );
xor \U$24307 ( \24650 , \24649 , \24300 );
xor \U$24308 ( \24651 , \24353 , \24360 );
xor \U$24309 ( \24652 , \24650 , \24651 );
and \U$24310 ( \24653 , \24648 , \24652 );
xor \U$24311 ( \24654 , \23464 , \23491 );
xor \U$24312 ( \24655 , \24654 , \23517 );
xor \U$24313 ( \24656 , \24290 , \24303 );
xor \U$24314 ( \24657 , \24655 , \24656 );
xor \U$24315 ( \24658 , \24653 , \24657 );
xor \U$24316 ( \24659 , \24412 , \2034 );
xor \U$24317 ( \24660 , \24659 , \24420 );
xor \U$24318 ( \24661 , \24431 , \24438 );
xor \U$24319 ( \24662 , \24661 , \24446 );
and \U$24320 ( \24663 , \24660 , \24662 );
xor \U$24321 ( \24664 , \24386 , \24393 );
xor \U$24322 ( \24665 , \24664 , \24401 );
xor \U$24323 ( \24666 , \24431 , \24438 );
xor \U$24324 ( \24667 , \24666 , \24446 );
and \U$24325 ( \24668 , \24665 , \24667 );
and \U$24326 ( \24669 , \24660 , \24665 );
or \U$24327 ( \24670 , \24663 , \24668 , \24669 );
xor \U$24328 ( \24671 , \24182 , \24190 );
xor \U$24329 ( \24672 , \24671 , \24198 );
xor \U$24330 ( \24673 , \24670 , \24672 );
xor \U$24331 ( \24674 , \24538 , \24545 );
xor \U$24332 ( \24675 , \24674 , \24554 );
xor \U$24333 ( \24676 , \24565 , \24572 );
xor \U$24334 ( \24677 , \24676 , \24580 );
and \U$24335 ( \24678 , \24675 , \24677 );
xor \U$24336 ( \24679 , \24513 , \24520 );
xor \U$24337 ( \24680 , \24679 , \24528 );
xor \U$24338 ( \24681 , \24565 , \24572 );
xor \U$24339 ( \24682 , \24681 , \24580 );
and \U$24340 ( \24683 , \24680 , \24682 );
and \U$24341 ( \24684 , \24675 , \24680 );
or \U$24342 ( \24685 , \24678 , \24683 , \24684 );
and \U$24343 ( \24686 , \24673 , \24685 );
and \U$24344 ( \24687 , \24670 , \24672 );
or \U$24345 ( \24688 , \24686 , \24687 );
and \U$24346 ( \24689 , \5318 , RI986ff70_75);
and \U$24347 ( \24690 , RI986fe80_73, \5316 );
nor \U$24348 ( \24691 , \24689 , \24690 );
and \U$24349 ( \24692 , \24691 , \5052 );
not \U$24350 ( \24693 , \24691 );
and \U$24351 ( \24694 , \24693 , \5322 );
nor \U$24352 ( \24695 , \24692 , \24694 );
and \U$24353 ( \24696 , \5881 , RI9870060_77);
and \U$24354 ( \24697 , RI9870150_79, \5879 );
nor \U$24355 ( \24698 , \24696 , \24697 );
and \U$24356 ( \24699 , \24698 , \5594 );
not \U$24357 ( \24700 , \24698 );
and \U$24358 ( \24701 , \24700 , \5885 );
nor \U$24359 ( \24702 , \24699 , \24701 );
xor \U$24360 ( \24703 , \24695 , \24702 );
and \U$24361 ( \24704 , \6453 , RI9870f60_109);
and \U$24362 ( \24705 , RI9870ab0_99, \6451 );
nor \U$24363 ( \24706 , \24704 , \24705 );
and \U$24364 ( \24707 , \24706 , \6190 );
not \U$24365 ( \24708 , \24706 );
and \U$24366 ( \24709 , \24708 , \6705 );
nor \U$24367 ( \24710 , \24707 , \24709 );
and \U$24368 ( \24711 , \24703 , \24710 );
and \U$24369 ( \24712 , \24695 , \24702 );
or \U$24370 ( \24713 , \24711 , \24712 );
not \U$24371 ( \24714 , \3412 );
and \U$24372 ( \24715 , \3683 , RI98708d0_95);
and \U$24373 ( \24716 , RI98707e0_93, \3681 );
nor \U$24374 ( \24717 , \24715 , \24716 );
not \U$24375 ( \24718 , \24717 );
or \U$24376 ( \24719 , \24714 , \24718 );
or \U$24377 ( \24720 , \24717 , \3918 );
nand \U$24378 ( \24721 , \24719 , \24720 );
and \U$24379 ( \24722 , \4203 , RI986fac0_65);
and \U$24380 ( \24723 , RI986fbb0_67, \4201 );
nor \U$24381 ( \24724 , \24722 , \24723 );
and \U$24382 ( \24725 , \24724 , \4207 );
not \U$24383 ( \24726 , \24724 );
and \U$24384 ( \24727 , \24726 , \3923 );
nor \U$24385 ( \24728 , \24725 , \24727 );
xor \U$24386 ( \24729 , \24721 , \24728 );
not \U$24387 ( \24730 , \4519 );
and \U$24388 ( \24731 , \4710 , RI986fd90_71);
and \U$24389 ( \24732 , RI986fca0_69, \4708 );
nor \U$24390 ( \24733 , \24731 , \24732 );
not \U$24391 ( \24734 , \24733 );
or \U$24392 ( \24735 , \24730 , \24734 );
or \U$24393 ( \24736 , \24733 , \4519 );
nand \U$24394 ( \24737 , \24735 , \24736 );
and \U$24395 ( \24738 , \24729 , \24737 );
and \U$24396 ( \24739 , \24721 , \24728 );
or \U$24397 ( \24740 , \24738 , \24739 );
xor \U$24398 ( \24741 , \24713 , \24740 );
and \U$24399 ( \24742 , \7079 , RI9870d80_105);
and \U$24400 ( \24743 , RI98709c0_97, \7077 );
nor \U$24401 ( \24744 , \24742 , \24743 );
and \U$24402 ( \24745 , \24744 , \6710 );
not \U$24403 ( \24746 , \24744 );
and \U$24404 ( \24747 , \24746 , \6709 );
nor \U$24405 ( \24748 , \24745 , \24747 );
and \U$24406 ( \24749 , \7729 , RI9870e70_107);
and \U$24407 ( \24750 , RI9870ba0_101, \7727 );
nor \U$24408 ( \24751 , \24749 , \24750 );
and \U$24409 ( \24752 , \24751 , \7480 );
not \U$24410 ( \24753 , \24751 );
and \U$24411 ( \24754 , \24753 , \7733 );
nor \U$24412 ( \24755 , \24752 , \24754 );
xor \U$24413 ( \24756 , \24748 , \24755 );
and \U$24414 ( \24757 , \8486 , RI9871050_111);
and \U$24415 ( \24758 , RI9870c90_103, \8484 );
nor \U$24416 ( \24759 , \24757 , \24758 );
and \U$24417 ( \24760 , \24759 , \8050 );
not \U$24418 ( \24761 , \24759 );
and \U$24419 ( \24762 , \24761 , \8051 );
nor \U$24420 ( \24763 , \24760 , \24762 );
and \U$24421 ( \24764 , \24756 , \24763 );
and \U$24422 ( \24765 , \24748 , \24755 );
or \U$24423 ( \24766 , \24764 , \24765 );
and \U$24424 ( \24767 , \24741 , \24766 );
and \U$24425 ( \24768 , \24713 , \24740 );
or \U$24426 ( \24769 , \24767 , \24768 );
and \U$24427 ( \24770 , \9237 , RI9871230_115);
and \U$24428 ( \24771 , RI9871140_113, \9235 );
nor \U$24429 ( \24772 , \24770 , \24771 );
and \U$24430 ( \24773 , \24772 , \9241 );
not \U$24431 ( \24774 , \24772 );
and \U$24432 ( \24775 , \24774 , \8836 );
nor \U$24433 ( \24776 , \24773 , \24775 );
and \U$24434 ( \24777 , \9505 , RI9871320_117);
and \U$24435 ( \24778 , RI9871410_119, \9503 );
nor \U$24436 ( \24779 , \24777 , \24778 );
and \U$24437 ( \24780 , \24779 , \9510 );
not \U$24438 ( \24781 , \24779 );
and \U$24439 ( \24782 , \24781 , \9513 );
nor \U$24440 ( \24783 , \24780 , \24782 );
xor \U$24441 ( \24784 , \24776 , \24783 );
and \U$24442 ( \24785 , \10424 , RI98716e0_125);
and \U$24443 ( \24786 , RI98717d0_127, \10422 );
nor \U$24444 ( \24787 , \24785 , \24786 );
and \U$24445 ( \24788 , \24787 , \9840 );
not \U$24446 ( \24789 , \24787 );
and \U$24447 ( \24790 , \24789 , \10428 );
nor \U$24448 ( \24791 , \24788 , \24790 );
and \U$24449 ( \24792 , \24784 , \24791 );
and \U$24450 ( \24793 , \24776 , \24783 );
or \U$24451 ( \24794 , \24792 , \24793 );
and \U$24452 ( \24795 , \13882 , RI986ee90_39);
and \U$24453 ( \24796 , RI986eda0_37, \13880 );
nor \U$24454 ( \24797 , \24795 , \24796 );
and \U$24455 ( \24798 , \24797 , \13358 );
not \U$24456 ( \24799 , \24797 );
and \U$24457 ( \24800 , \24799 , \13359 );
nor \U$24458 ( \24801 , \24798 , \24800 );
not \U$24459 ( \24802 , RI9873558_190);
and \U$24460 ( \24803 , \15780 , RI986f070_43);
and \U$24461 ( \24804 , RI9873648_192, RI986ef80_41);
nor \U$24462 ( \24805 , \24803 , \24804 );
not \U$24463 ( \24806 , \24805 );
or \U$24464 ( \24807 , \24802 , \24806 );
or \U$24465 ( \24808 , \24805 , RI9873558_190);
nand \U$24466 ( \24809 , \24807 , \24808 );
xor \U$24467 ( \24810 , \24801 , \24809 );
and \U$24468 ( \24811 , \14937 , RI986ebc0_33);
and \U$24469 ( \24812 , RI986ecb0_35, \14935 );
nor \U$24470 ( \24813 , \24811 , \24812 );
and \U$24471 ( \24814 , \24813 , \14539 );
not \U$24472 ( \24815 , \24813 );
and \U$24473 ( \24816 , \24815 , \14538 );
nor \U$24474 ( \24817 , \24814 , \24816 );
and \U$24475 ( \24818 , \24810 , \24817 );
and \U$24476 ( \24819 , \24801 , \24809 );
or \U$24477 ( \24820 , \24818 , \24819 );
xor \U$24478 ( \24821 , \24794 , \24820 );
and \U$24479 ( \24822 , \13045 , RI986e8f0_27);
and \U$24480 ( \24823 , RI986e800_25, \13043 );
nor \U$24481 ( \24824 , \24822 , \24823 );
and \U$24482 ( \24825 , \24824 , \13047 );
not \U$24483 ( \24826 , \24824 );
and \U$24484 ( \24827 , \24826 , \12619 );
nor \U$24485 ( \24828 , \24825 , \24827 );
and \U$24486 ( \24829 , \11696 , RI9871500_121);
and \U$24487 ( \24830 , RI98715f0_123, \11694 );
nor \U$24488 ( \24831 , \24829 , \24830 );
and \U$24489 ( \24832 , \24831 , \10965 );
not \U$24490 ( \24833 , \24831 );
and \U$24491 ( \24834 , \24833 , \11702 );
nor \U$24492 ( \24835 , \24832 , \24834 );
xor \U$24493 ( \24836 , \24828 , \24835 );
and \U$24494 ( \24837 , \12293 , RI986ead0_31);
and \U$24495 ( \24838 , RI986e9e0_29, \12291 );
nor \U$24496 ( \24839 , \24837 , \24838 );
and \U$24497 ( \24840 , \24839 , \11687 );
not \U$24498 ( \24841 , \24839 );
and \U$24499 ( \24842 , \24841 , \11686 );
nor \U$24500 ( \24843 , \24840 , \24842 );
and \U$24501 ( \24844 , \24836 , \24843 );
and \U$24502 ( \24845 , \24828 , \24835 );
or \U$24503 ( \24846 , \24844 , \24845 );
and \U$24504 ( \24847 , \24821 , \24846 );
and \U$24505 ( \24848 , \24794 , \24820 );
or \U$24506 ( \24849 , \24847 , \24848 );
xor \U$24507 ( \24850 , \24769 , \24849 );
and \U$24508 ( \24851 , \2274 , RI9870420_85);
and \U$24509 ( \24852 , RI9870510_87, \2272 );
nor \U$24510 ( \24853 , \24851 , \24852 );
and \U$24511 ( \24854 , \24853 , \2030 );
not \U$24512 ( \24855 , \24853 );
and \U$24513 ( \24856 , \24855 , \2031 );
nor \U$24514 ( \24857 , \24854 , \24856 );
and \U$24515 ( \24858 , \2464 , RI9870330_83);
and \U$24516 ( \24859 , RI9870240_81, \2462 );
nor \U$24517 ( \24860 , \24858 , \24859 );
and \U$24518 ( \24861 , \24860 , \2468 );
not \U$24519 ( \24862 , \24860 );
and \U$24520 ( \24863 , \24862 , \2263 );
nor \U$24521 ( \24864 , \24861 , \24863 );
xor \U$24522 ( \24865 , \24857 , \24864 );
not \U$24523 ( \24866 , \2935 );
and \U$24524 ( \24867 , \3254 , RI98706f0_91);
and \U$24525 ( \24868 , RI9870600_89, \3252 );
nor \U$24526 ( \24869 , \24867 , \24868 );
not \U$24527 ( \24870 , \24869 );
or \U$24528 ( \24871 , \24866 , \24870 );
or \U$24529 ( \24872 , \24869 , \3406 );
nand \U$24530 ( \24873 , \24871 , \24872 );
and \U$24531 ( \24874 , \24865 , \24873 );
and \U$24532 ( \24875 , \24857 , \24864 );
or \U$24533 ( \24876 , \24874 , \24875 );
xor \U$24534 ( \24877 , \24458 , \24465 );
xor \U$24535 ( \24878 , \24876 , \24877 );
xor \U$24536 ( \24879 , \24482 , \24490 );
xor \U$24537 ( \24880 , \24879 , \24499 );
and \U$24538 ( \24881 , \24878 , \24880 );
and \U$24539 ( \24882 , \24876 , \24877 );
or \U$24540 ( \24883 , \24881 , \24882 );
and \U$24541 ( \24884 , \24850 , \24883 );
and \U$24542 ( \24885 , \24769 , \24849 );
or \U$24543 ( \24886 , \24884 , \24885 );
xor \U$24544 ( \24887 , \24688 , \24886 );
xor \U$24545 ( \24888 , \24466 , \24474 );
xor \U$24546 ( \24889 , \24888 , \24502 );
xor \U$24547 ( \24890 , \24604 , \24606 );
xor \U$24548 ( \24891 , \24890 , \24609 );
and \U$24549 ( \24892 , \24889 , \24891 );
xor \U$24550 ( \24893 , \24129 , \24136 );
xor \U$24551 ( \24894 , \24893 , \24144 );
xor \U$24552 ( \24895 , \24592 , \24597 );
xor \U$24553 ( \24896 , \24894 , \24895 );
xor \U$24554 ( \24897 , \24604 , \24606 );
xor \U$24555 ( \24898 , \24897 , \24609 );
and \U$24556 ( \24899 , \24896 , \24898 );
and \U$24557 ( \24900 , \24889 , \24896 );
or \U$24558 ( \24901 , \24892 , \24899 , \24900 );
and \U$24559 ( \24902 , \24887 , \24901 );
and \U$24560 ( \24903 , \24688 , \24886 );
or \U$24561 ( \24904 , \24902 , \24903 );
xor \U$24562 ( \24905 , \24150 , \24230 );
xor \U$24563 ( \24906 , \24905 , \24267 );
xor \U$24564 ( \24907 , \24904 , \24906 );
xor \U$24565 ( \24908 , \24175 , \24201 );
xor \U$24566 ( \24909 , \24908 , \24227 );
xor \U$24567 ( \24910 , \24602 , \24612 );
xor \U$24568 ( \24911 , \24910 , \24617 );
and \U$24569 ( \24912 , \24909 , \24911 );
xor \U$24570 ( \24913 , \24058 , \24060 );
xor \U$24571 ( \24914 , \24913 , \24063 );
xor \U$24572 ( \24915 , \24367 , \24374 );
xor \U$24573 ( \24916 , \24914 , \24915 );
xor \U$24574 ( \24917 , \24602 , \24612 );
xor \U$24575 ( \24918 , \24917 , \24617 );
and \U$24576 ( \24919 , \24916 , \24918 );
and \U$24577 ( \24920 , \24909 , \24916 );
or \U$24578 ( \24921 , \24912 , \24919 , \24920 );
and \U$24579 ( \24922 , \24907 , \24921 );
and \U$24580 ( \24923 , \24904 , \24906 );
or \U$24581 ( \24924 , \24922 , \24923 );
and \U$24582 ( \24925 , \24658 , \24924 );
and \U$24583 ( \24926 , \24653 , \24657 );
or \U$24584 ( \24927 , \24925 , \24926 );
nand \U$24585 ( \24928 , \24646 , \24927 );
nand \U$24586 ( \24929 , \24645 , \24928 );
xor \U$24587 ( \24930 , \24326 , \24337 );
xor \U$24588 ( \24931 , \24930 , \24342 );
xor \U$24589 ( \24932 , \23991 , \23996 );
xor \U$24590 ( \24933 , \24932 , \24013 );
xor \U$24591 ( \24934 , \24931 , \24933 );
xor \U$24592 ( \24935 , \24635 , \24637 );
and \U$24593 ( \24936 , \24935 , \24642 );
and \U$24594 ( \24937 , \24635 , \24637 );
or \U$24595 ( \24938 , \24936 , \24937 );
xor \U$24596 ( \24939 , \24934 , \24938 );
and \U$24597 ( \24940 , \24929 , \24939 );
xor \U$24598 ( \24941 , \24939 , \24929 );
xor \U$24599 ( \24942 , \24351 , \24629 );
xor \U$24600 ( \24943 , \24648 , \24652 );
xor \U$24601 ( \24944 , \24531 , \24557 );
xor \U$24602 ( \24945 , \24944 , \24583 );
xor \U$24603 ( \24946 , \24404 , \24423 );
xor \U$24604 ( \24947 , \24946 , \24449 );
xor \U$24605 ( \24948 , \24945 , \24947 );
xor \U$24606 ( \24949 , \24604 , \24606 );
xor \U$24607 ( \24950 , \24949 , \24609 );
xor \U$24608 ( \24951 , \24889 , \24896 );
xor \U$24609 ( \24952 , \24950 , \24951 );
and \U$24610 ( \24953 , \24948 , \24952 );
and \U$24611 ( \24954 , \24945 , \24947 );
or \U$24612 ( \24955 , \24953 , \24954 );
xor \U$24613 ( \24956 , \24452 , \24505 );
xor \U$24614 ( \24957 , \24956 , \24586 );
xor \U$24615 ( \24958 , \24955 , \24957 );
xor \U$24616 ( \24959 , \24713 , \24740 );
xor \U$24617 ( \24960 , \24959 , \24766 );
xor \U$24618 ( \24961 , \24876 , \24877 );
xor \U$24619 ( \24962 , \24961 , \24880 );
and \U$24620 ( \24963 , \24960 , \24962 );
xor \U$24621 ( \24964 , \24565 , \24572 );
xor \U$24622 ( \24965 , \24964 , \24580 );
xor \U$24623 ( \24966 , \24675 , \24680 );
xor \U$24624 ( \24967 , \24965 , \24966 );
xor \U$24625 ( \24968 , \24876 , \24877 );
xor \U$24626 ( \24969 , \24968 , \24880 );
and \U$24627 ( \24970 , \24967 , \24969 );
and \U$24628 ( \24971 , \24960 , \24967 );
or \U$24629 ( \24972 , \24963 , \24970 , \24971 );
and \U$24630 ( \24973 , \7729 , RI98709c0_97);
and \U$24631 ( \24974 , RI9870e70_107, \7727 );
nor \U$24632 ( \24975 , \24973 , \24974 );
and \U$24633 ( \24976 , \24975 , \7480 );
not \U$24634 ( \24977 , \24975 );
and \U$24635 ( \24978 , \24977 , \7733 );
nor \U$24636 ( \24979 , \24976 , \24978 );
and \U$24637 ( \24980 , \8486 , RI9870ba0_101);
and \U$24638 ( \24981 , RI9871050_111, \8484 );
nor \U$24639 ( \24982 , \24980 , \24981 );
and \U$24640 ( \24983 , \24982 , \8050 );
not \U$24641 ( \24984 , \24982 );
and \U$24642 ( \24985 , \24984 , \8051 );
nor \U$24643 ( \24986 , \24983 , \24985 );
xor \U$24644 ( \24987 , \24979 , \24986 );
and \U$24645 ( \24988 , \9237 , RI9870c90_103);
and \U$24646 ( \24989 , RI9871230_115, \9235 );
nor \U$24647 ( \24990 , \24988 , \24989 );
and \U$24648 ( \24991 , \24990 , \9241 );
not \U$24649 ( \24992 , \24990 );
and \U$24650 ( \24993 , \24992 , \8836 );
nor \U$24651 ( \24994 , \24991 , \24993 );
and \U$24652 ( \24995 , \24987 , \24994 );
and \U$24653 ( \24996 , \24979 , \24986 );
or \U$24654 ( \24997 , \24995 , \24996 );
and \U$24655 ( \24998 , \4203 , RI98707e0_93);
and \U$24656 ( \24999 , RI986fac0_65, \4201 );
nor \U$24657 ( \25000 , \24998 , \24999 );
and \U$24658 ( \25001 , \25000 , \4207 );
not \U$24659 ( \25002 , \25000 );
and \U$24660 ( \25003 , \25002 , \3922 );
nor \U$24661 ( \25004 , \25001 , \25003 );
not \U$24662 ( \25005 , \4519 );
and \U$24663 ( \25006 , \4710 , RI986fbb0_67);
and \U$24664 ( \25007 , RI986fd90_71, \4708 );
nor \U$24665 ( \25008 , \25006 , \25007 );
not \U$24666 ( \25009 , \25008 );
or \U$24667 ( \25010 , \25005 , \25009 );
or \U$24668 ( \25011 , \25008 , \4519 );
nand \U$24669 ( \25012 , \25010 , \25011 );
xor \U$24670 ( \25013 , \25004 , \25012 );
and \U$24671 ( \25014 , \5318 , RI986fca0_69);
and \U$24672 ( \25015 , RI986ff70_75, \5316 );
nor \U$24673 ( \25016 , \25014 , \25015 );
and \U$24674 ( \25017 , \25016 , \5052 );
not \U$24675 ( \25018 , \25016 );
and \U$24676 ( \25019 , \25018 , \5322 );
nor \U$24677 ( \25020 , \25017 , \25019 );
and \U$24678 ( \25021 , \25013 , \25020 );
and \U$24679 ( \25022 , \25004 , \25012 );
or \U$24680 ( \25023 , \25021 , \25022 );
xor \U$24681 ( \25024 , \24997 , \25023 );
and \U$24682 ( \25025 , \5881 , RI986fe80_73);
and \U$24683 ( \25026 , RI9870060_77, \5879 );
nor \U$24684 ( \25027 , \25025 , \25026 );
and \U$24685 ( \25028 , \25027 , \5594 );
not \U$24686 ( \25029 , \25027 );
and \U$24687 ( \25030 , \25029 , \5885 );
nor \U$24688 ( \25031 , \25028 , \25030 );
and \U$24689 ( \25032 , \6453 , RI9870150_79);
and \U$24690 ( \25033 , RI9870f60_109, \6451 );
nor \U$24691 ( \25034 , \25032 , \25033 );
and \U$24692 ( \25035 , \25034 , \6190 );
not \U$24693 ( \25036 , \25034 );
and \U$24694 ( \25037 , \25036 , \6180 );
nor \U$24695 ( \25038 , \25035 , \25037 );
xor \U$24696 ( \25039 , \25031 , \25038 );
and \U$24697 ( \25040 , \7079 , RI9870ab0_99);
and \U$24698 ( \25041 , RI9870d80_105, \7077 );
nor \U$24699 ( \25042 , \25040 , \25041 );
and \U$24700 ( \25043 , \25042 , \6710 );
not \U$24701 ( \25044 , \25042 );
and \U$24702 ( \25045 , \25044 , \6709 );
nor \U$24703 ( \25046 , \25043 , \25045 );
and \U$24704 ( \25047 , \25039 , \25046 );
and \U$24705 ( \25048 , \25031 , \25038 );
or \U$24706 ( \25049 , \25047 , \25048 );
and \U$24707 ( \25050 , \25024 , \25049 );
and \U$24708 ( \25051 , \24997 , \25023 );
or \U$24709 ( \25052 , \25050 , \25051 );
and \U$24710 ( \25053 , \9505 , RI9871140_113);
and \U$24711 ( \25054 , RI9871320_117, \9503 );
nor \U$24712 ( \25055 , \25053 , \25054 );
and \U$24713 ( \25056 , \25055 , \9510 );
not \U$24714 ( \25057 , \25055 );
and \U$24715 ( \25058 , \25057 , \9513 );
nor \U$24716 ( \25059 , \25056 , \25058 );
and \U$24717 ( \25060 , \10424 , RI9871410_119);
and \U$24718 ( \25061 , RI98716e0_125, \10422 );
nor \U$24719 ( \25062 , \25060 , \25061 );
and \U$24720 ( \25063 , \25062 , \9840 );
not \U$24721 ( \25064 , \25062 );
and \U$24722 ( \25065 , \25064 , \10428 );
nor \U$24723 ( \25066 , \25063 , \25065 );
xor \U$24724 ( \25067 , \25059 , \25066 );
and \U$24725 ( \25068 , \11696 , RI98717d0_127);
and \U$24726 ( \25069 , RI9871500_121, \11694 );
nor \U$24727 ( \25070 , \25068 , \25069 );
and \U$24728 ( \25071 , \25070 , \10965 );
not \U$24729 ( \25072 , \25070 );
and \U$24730 ( \25073 , \25072 , \11702 );
nor \U$24731 ( \25074 , \25071 , \25073 );
and \U$24732 ( \25075 , \25067 , \25074 );
and \U$24733 ( \25076 , \25059 , \25066 );
or \U$24734 ( \25077 , \25075 , \25076 );
not \U$24735 ( \25078 , RI9873558_190);
and \U$24736 ( \25079 , \15780 , RI986ecb0_35);
and \U$24737 ( \25080 , RI9873648_192, RI986f070_43);
nor \U$24738 ( \25081 , \25079 , \25080 );
not \U$24739 ( \25082 , \25081 );
or \U$24740 ( \25083 , \25078 , \25082 );
or \U$24741 ( \25084 , \25081 , RI9873558_190);
nand \U$24742 ( \25085 , \25083 , \25084 );
xor \U$24743 ( \25086 , \25085 , \2031 );
and \U$24744 ( \25087 , \14937 , RI986eda0_37);
and \U$24745 ( \25088 , RI986ebc0_33, \14935 );
nor \U$24746 ( \25089 , \25087 , \25088 );
and \U$24747 ( \25090 , \25089 , \14539 );
not \U$24748 ( \25091 , \25089 );
and \U$24749 ( \25092 , \25091 , \14538 );
nor \U$24750 ( \25093 , \25090 , \25092 );
and \U$24751 ( \25094 , \25086 , \25093 );
and \U$24752 ( \25095 , \25085 , \2031 );
or \U$24753 ( \25096 , \25094 , \25095 );
xor \U$24754 ( \25097 , \25077 , \25096 );
and \U$24755 ( \25098 , \13882 , RI986e800_25);
and \U$24756 ( \25099 , RI986ee90_39, \13880 );
nor \U$24757 ( \25100 , \25098 , \25099 );
and \U$24758 ( \25101 , \25100 , \13358 );
not \U$24759 ( \25102 , \25100 );
and \U$24760 ( \25103 , \25102 , \13359 );
nor \U$24761 ( \25104 , \25101 , \25103 );
and \U$24762 ( \25105 , \12293 , RI98715f0_123);
and \U$24763 ( \25106 , RI986ead0_31, \12291 );
nor \U$24764 ( \25107 , \25105 , \25106 );
and \U$24765 ( \25108 , \25107 , \11687 );
not \U$24766 ( \25109 , \25107 );
and \U$24767 ( \25110 , \25109 , \11686 );
nor \U$24768 ( \25111 , \25108 , \25110 );
xor \U$24769 ( \25112 , \25104 , \25111 );
and \U$24770 ( \25113 , \13045 , RI986e9e0_29);
and \U$24771 ( \25114 , RI986e8f0_27, \13043 );
nor \U$24772 ( \25115 , \25113 , \25114 );
and \U$24773 ( \25116 , \25115 , \13047 );
not \U$24774 ( \25117 , \25115 );
and \U$24775 ( \25118 , \25117 , \12619 );
nor \U$24776 ( \25119 , \25116 , \25118 );
and \U$24777 ( \25120 , \25112 , \25119 );
and \U$24778 ( \25121 , \25104 , \25111 );
or \U$24779 ( \25122 , \25120 , \25121 );
and \U$24780 ( \25123 , \25097 , \25122 );
and \U$24781 ( \25124 , \25077 , \25096 );
or \U$24782 ( \25125 , \25123 , \25124 );
xor \U$24783 ( \25126 , \25052 , \25125 );
and \U$24784 ( \25127 , \2464 , RI9870510_87);
and \U$24785 ( \25128 , RI9870330_83, \2462 );
nor \U$24786 ( \25129 , \25127 , \25128 );
and \U$24787 ( \25130 , \25129 , \2468 );
not \U$24788 ( \25131 , \25129 );
and \U$24789 ( \25132 , \25131 , \2263 );
nor \U$24790 ( \25133 , \25130 , \25132 );
not \U$24791 ( \25134 , \2935 );
and \U$24792 ( \25135 , \3254 , RI9870240_81);
and \U$24793 ( \25136 , RI98706f0_91, \3252 );
nor \U$24794 ( \25137 , \25135 , \25136 );
not \U$24795 ( \25138 , \25137 );
or \U$24796 ( \25139 , \25134 , \25138 );
or \U$24797 ( \25140 , \25137 , \3406 );
nand \U$24798 ( \25141 , \25139 , \25140 );
xor \U$24799 ( \25142 , \25133 , \25141 );
not \U$24800 ( \25143 , \3918 );
and \U$24801 ( \25144 , \3683 , RI9870600_89);
and \U$24802 ( \25145 , RI98708d0_95, \3681 );
nor \U$24803 ( \25146 , \25144 , \25145 );
not \U$24804 ( \25147 , \25146 );
or \U$24805 ( \25148 , \25143 , \25147 );
or \U$24806 ( \25149 , \25146 , \3918 );
nand \U$24807 ( \25150 , \25148 , \25149 );
and \U$24808 ( \25151 , \25142 , \25150 );
and \U$24809 ( \25152 , \25133 , \25141 );
or \U$24810 ( \25153 , \25151 , \25152 );
xor \U$24811 ( \25154 , \24857 , \24864 );
xor \U$24812 ( \25155 , \25154 , \24873 );
and \U$24813 ( \25156 , \25153 , \25155 );
xor \U$24814 ( \25157 , \24721 , \24728 );
xor \U$24815 ( \25158 , \25157 , \24737 );
xor \U$24816 ( \25159 , \24857 , \24864 );
xor \U$24817 ( \25160 , \25159 , \24873 );
and \U$24818 ( \25161 , \25158 , \25160 );
and \U$24819 ( \25162 , \25153 , \25158 );
or \U$24820 ( \25163 , \25156 , \25161 , \25162 );
and \U$24821 ( \25164 , \25126 , \25163 );
and \U$24822 ( \25165 , \25052 , \25125 );
or \U$24823 ( \25166 , \25164 , \25165 );
xor \U$24824 ( \25167 , \24972 , \25166 );
xor \U$24825 ( \25168 , \24695 , \24702 );
xor \U$24826 ( \25169 , \25168 , \24710 );
xor \U$24827 ( \25170 , \24776 , \24783 );
xor \U$24828 ( \25171 , \25170 , \24791 );
and \U$24829 ( \25172 , \25169 , \25171 );
xor \U$24830 ( \25173 , \24748 , \24755 );
xor \U$24831 ( \25174 , \25173 , \24763 );
xor \U$24832 ( \25175 , \24776 , \24783 );
xor \U$24833 ( \25176 , \25175 , \24791 );
and \U$24834 ( \25177 , \25174 , \25176 );
and \U$24835 ( \25178 , \25169 , \25174 );
or \U$24836 ( \25179 , \25172 , \25177 , \25178 );
xor \U$24837 ( \25180 , \24828 , \24835 );
xor \U$24838 ( \25181 , \25180 , \24843 );
xor \U$24839 ( \25182 , \24801 , \24809 );
xor \U$24840 ( \25183 , \25182 , \24817 );
and \U$24841 ( \25184 , \25181 , \25183 );
xor \U$24842 ( \25185 , \25179 , \25184 );
xor \U$24843 ( \25186 , \24431 , \24438 );
xor \U$24844 ( \25187 , \25186 , \24446 );
xor \U$24845 ( \25188 , \24660 , \24665 );
xor \U$24846 ( \25189 , \25187 , \25188 );
and \U$24847 ( \25190 , \25185 , \25189 );
and \U$24848 ( \25191 , \25179 , \25184 );
or \U$24849 ( \25192 , \25190 , \25191 );
and \U$24850 ( \25193 , \25167 , \25192 );
and \U$24851 ( \25194 , \24972 , \25166 );
or \U$24852 ( \25195 , \25193 , \25194 );
and \U$24853 ( \25196 , \24958 , \25195 );
and \U$24854 ( \25197 , \24955 , \24957 );
or \U$24855 ( \25198 , \25196 , \25197 );
xor \U$24856 ( \25199 , \24943 , \25198 );
xor \U$24857 ( \25200 , \24904 , \24906 );
xor \U$24858 ( \25201 , \25200 , \24921 );
and \U$24859 ( \25202 , \25199 , \25201 );
and \U$24860 ( \25203 , \24943 , \25198 );
or \U$24861 ( \25204 , \25202 , \25203 );
xor \U$24862 ( \25205 , \24942 , \25204 );
xor \U$24863 ( \25206 , \24653 , \24657 );
xor \U$24864 ( \25207 , \25206 , \24924 );
xor \U$24865 ( \25208 , \25205 , \25207 );
xor \U$24866 ( \25209 , \24688 , \24886 );
xor \U$24867 ( \25210 , \25209 , \24901 );
xor \U$24868 ( \25211 , \24955 , \24957 );
xor \U$24869 ( \25212 , \25211 , \25195 );
and \U$24870 ( \25213 , \25210 , \25212 );
not \U$24871 ( \25214 , \25213 );
xor \U$24872 ( \25215 , \24943 , \25198 );
xor \U$24873 ( \25216 , \25215 , \25201 );
not \U$24874 ( \25217 , \25216 );
or \U$24875 ( \25218 , \25214 , \25217 );
or \U$24876 ( \25219 , \25216 , \25213 );
xor \U$24877 ( \25220 , \24769 , \24849 );
xor \U$24878 ( \25221 , \25220 , \24883 );
xor \U$24879 ( \25222 , \24945 , \24947 );
xor \U$24880 ( \25223 , \25222 , \24952 );
and \U$24881 ( \25224 , \25221 , \25223 );
xor \U$24882 ( \25225 , \24972 , \25166 );
xor \U$24883 ( \25226 , \25225 , \25192 );
xor \U$24884 ( \25227 , \24945 , \24947 );
xor \U$24885 ( \25228 , \25227 , \24952 );
and \U$24886 ( \25229 , \25226 , \25228 );
and \U$24887 ( \25230 , \25221 , \25226 );
or \U$24888 ( \25231 , \25224 , \25229 , \25230 );
xor \U$24889 ( \25232 , \24602 , \24612 );
xor \U$24890 ( \25233 , \25232 , \24617 );
xor \U$24891 ( \25234 , \24909 , \24916 );
xor \U$24892 ( \25235 , \25233 , \25234 );
xor \U$24893 ( \25236 , \25231 , \25235 );
xor \U$24894 ( \25237 , \24997 , \25023 );
xor \U$24895 ( \25238 , \25237 , \25049 );
xor \U$24896 ( \25239 , \25077 , \25096 );
xor \U$24897 ( \25240 , \25239 , \25122 );
xor \U$24898 ( \25241 , \25238 , \25240 );
xor \U$24899 ( \25242 , \24857 , \24864 );
xor \U$24900 ( \25243 , \25242 , \24873 );
xor \U$24901 ( \25244 , \25153 , \25158 );
xor \U$24902 ( \25245 , \25243 , \25244 );
and \U$24903 ( \25246 , \25241 , \25245 );
and \U$24904 ( \25247 , \25238 , \25240 );
or \U$24905 ( \25248 , \25246 , \25247 );
and \U$24906 ( \25249 , \7729 , RI9870d80_105);
and \U$24907 ( \25250 , RI98709c0_97, \7727 );
nor \U$24908 ( \25251 , \25249 , \25250 );
and \U$24909 ( \25252 , \25251 , \7733 );
not \U$24910 ( \25253 , \25251 );
and \U$24911 ( \25254 , \25253 , \7480 );
nor \U$24912 ( \25255 , \25252 , \25254 );
and \U$24913 ( \25256 , \8486 , RI9870e70_107);
and \U$24914 ( \25257 , RI9870ba0_101, \8484 );
nor \U$24915 ( \25258 , \25256 , \25257 );
and \U$24916 ( \25259 , \25258 , \8051 );
not \U$24917 ( \25260 , \25258 );
and \U$24918 ( \25261 , \25260 , \8050 );
nor \U$24919 ( \25262 , \25259 , \25261 );
xor \U$24920 ( \25263 , \25255 , \25262 );
and \U$24921 ( \25264 , \7079 , RI9870f60_109);
and \U$24922 ( \25265 , RI9870ab0_99, \7077 );
nor \U$24923 ( \25266 , \25264 , \25265 );
and \U$24924 ( \25267 , \25266 , \6709 );
not \U$24925 ( \25268 , \25266 );
and \U$24926 ( \25269 , \25268 , \6710 );
nor \U$24927 ( \25270 , \25267 , \25269 );
and \U$24928 ( \25271 , \25263 , \25270 );
and \U$24929 ( \25272 , \25255 , \25262 );
nor \U$24930 ( \25273 , \25271 , \25272 );
and \U$24931 ( \25274 , \5318 , RI986fd90_71);
and \U$24932 ( \25275 , RI986fca0_69, \5316 );
nor \U$24933 ( \25276 , \25274 , \25275 );
and \U$24934 ( \25277 , \25276 , \5052 );
not \U$24935 ( \25278 , \25276 );
and \U$24936 ( \25279 , \25278 , \5322 );
nor \U$24937 ( \25280 , \25277 , \25279 );
and \U$24938 ( \25281 , \5881 , RI986ff70_75);
and \U$24939 ( \25282 , RI986fe80_73, \5879 );
nor \U$24940 ( \25283 , \25281 , \25282 );
and \U$24941 ( \25284 , \25283 , \5594 );
not \U$24942 ( \25285 , \25283 );
and \U$24943 ( \25286 , \25285 , \5885 );
nor \U$24944 ( \25287 , \25284 , \25286 );
xor \U$24945 ( \25288 , \25280 , \25287 );
and \U$24946 ( \25289 , \6453 , RI9870060_77);
and \U$24947 ( \25290 , RI9870150_79, \6451 );
nor \U$24948 ( \25291 , \25289 , \25290 );
and \U$24949 ( \25292 , \25291 , \6190 );
not \U$24950 ( \25293 , \25291 );
and \U$24951 ( \25294 , \25293 , \6705 );
nor \U$24952 ( \25295 , \25292 , \25294 );
and \U$24953 ( \25296 , \25288 , \25295 );
and \U$24954 ( \25297 , \25280 , \25287 );
or \U$24955 ( \25298 , \25296 , \25297 );
xor \U$24956 ( \25299 , \25273 , \25298 );
and \U$24957 ( \25300 , \4203 , RI98708d0_95);
and \U$24958 ( \25301 , RI98707e0_93, \4201 );
nor \U$24959 ( \25302 , \25300 , \25301 );
and \U$24960 ( \25303 , \25302 , \3922 );
not \U$24961 ( \25304 , \25302 );
and \U$24962 ( \25305 , \25304 , \4207 );
nor \U$24963 ( \25306 , \25303 , \25305 );
and \U$24964 ( \25307 , \4710 , RI986fac0_65);
and \U$24965 ( \25308 , RI986fbb0_67, \4708 );
nor \U$24966 ( \25309 , \25307 , \25308 );
not \U$24967 ( \25310 , \25309 );
not \U$24968 ( \25311 , \4521 );
and \U$24969 ( \25312 , \25310 , \25311 );
and \U$24970 ( \25313 , \25309 , \4519 );
nor \U$24971 ( \25314 , \25312 , \25313 );
xor \U$24972 ( \25315 , \25306 , \25314 );
and \U$24973 ( \25316 , \3683 , RI98706f0_91);
and \U$24974 ( \25317 , RI9870600_89, \3681 );
nor \U$24975 ( \25318 , \25316 , \25317 );
not \U$24976 ( \25319 , \25318 );
not \U$24977 ( \25320 , \3918 );
and \U$24978 ( \25321 , \25319 , \25320 );
and \U$24979 ( \25322 , \25318 , \3918 );
nor \U$24980 ( \25323 , \25321 , \25322 );
and \U$24981 ( \25324 , \25315 , \25323 );
and \U$24982 ( \25325 , \25306 , \25314 );
nor \U$24983 ( \25326 , \25324 , \25325 );
and \U$24984 ( \25327 , \25299 , \25326 );
and \U$24985 ( \25328 , \25273 , \25298 );
or \U$24986 ( \25329 , \25327 , \25328 );
and \U$24987 ( \25330 , \9237 , RI9871050_111);
and \U$24988 ( \25331 , RI9870c90_103, \9235 );
nor \U$24989 ( \25332 , \25330 , \25331 );
and \U$24990 ( \25333 , \25332 , \8836 );
not \U$24991 ( \25334 , \25332 );
and \U$24992 ( \25335 , \25334 , \9241 );
nor \U$24993 ( \25336 , \25333 , \25335 );
and \U$24994 ( \25337 , \10424 , RI9871320_117);
and \U$24995 ( \25338 , RI9871410_119, \10422 );
nor \U$24996 ( \25339 , \25337 , \25338 );
and \U$24997 ( \25340 , \25339 , \10428 );
not \U$24998 ( \25341 , \25339 );
and \U$24999 ( \25342 , \25341 , \9840 );
nor \U$25000 ( \25343 , \25340 , \25342 );
or \U$25001 ( \25344 , \25336 , \25343 );
not \U$25002 ( \25345 , \25343 );
not \U$25003 ( \25346 , \25336 );
or \U$25004 ( \25347 , \25345 , \25346 );
and \U$25005 ( \25348 , \9505 , RI9871230_115);
and \U$25006 ( \25349 , RI9871140_113, \9503 );
nor \U$25007 ( \25350 , \25348 , \25349 );
and \U$25008 ( \25351 , \25350 , \9510 );
not \U$25009 ( \25352 , \25350 );
and \U$25010 ( \25353 , \25352 , \9513 );
nor \U$25011 ( \25354 , \25351 , \25353 );
nand \U$25012 ( \25355 , \25347 , \25354 );
nand \U$25013 ( \25356 , \25344 , \25355 );
and \U$25014 ( \25357 , \15780 , RI986ebc0_33);
and \U$25015 ( \25358 , RI9873648_192, RI986ecb0_35);
nor \U$25016 ( \25359 , \25357 , \25358 );
not \U$25017 ( \25360 , \25359 );
not \U$25018 ( \25361 , RI9873558_190);
and \U$25019 ( \25362 , \25360 , \25361 );
and \U$25020 ( \25363 , \25359 , RI9873558_190);
nor \U$25021 ( \25364 , \25362 , \25363 );
and \U$25022 ( \25365 , \14937 , RI986ee90_39);
and \U$25023 ( \25366 , RI986eda0_37, \14935 );
nor \U$25024 ( \25367 , \25365 , \25366 );
and \U$25025 ( \25368 , \25367 , \14538 );
not \U$25026 ( \25369 , \25367 );
and \U$25027 ( \25370 , \25369 , \14539 );
nor \U$25028 ( \25371 , \25368 , \25370 );
xor \U$25029 ( \25372 , \25364 , \25371 );
and \U$25030 ( \25373 , \13882 , RI986e8f0_27);
and \U$25031 ( \25374 , RI986e800_25, \13880 );
nor \U$25032 ( \25375 , \25373 , \25374 );
and \U$25033 ( \25376 , \25375 , \13359 );
not \U$25034 ( \25377 , \25375 );
and \U$25035 ( \25378 , \25377 , \13358 );
nor \U$25036 ( \25379 , \25376 , \25378 );
and \U$25037 ( \25380 , \25372 , \25379 );
and \U$25038 ( \25381 , \25364 , \25371 );
nor \U$25039 ( \25382 , \25380 , \25381 );
xor \U$25040 ( \25383 , \25356 , \25382 );
and \U$25041 ( \25384 , \12293 , RI9871500_121);
and \U$25042 ( \25385 , RI98715f0_123, \12291 );
nor \U$25043 ( \25386 , \25384 , \25385 );
and \U$25044 ( \25387 , \25386 , \11687 );
not \U$25045 ( \25388 , \25386 );
and \U$25046 ( \25389 , \25388 , \11686 );
nor \U$25047 ( \25390 , \25387 , \25389 );
and \U$25048 ( \25391 , \11696 , RI98716e0_125);
and \U$25049 ( \25392 , RI98717d0_127, \11694 );
nor \U$25050 ( \25393 , \25391 , \25392 );
and \U$25051 ( \25394 , \25393 , \10965 );
not \U$25052 ( \25395 , \25393 );
and \U$25053 ( \25396 , \25395 , \11702 );
nor \U$25054 ( \25397 , \25394 , \25396 );
xor \U$25055 ( \25398 , \25390 , \25397 );
and \U$25056 ( \25399 , \13045 , RI986ead0_31);
and \U$25057 ( \25400 , RI986e9e0_29, \13043 );
nor \U$25058 ( \25401 , \25399 , \25400 );
and \U$25059 ( \25402 , \25401 , \13047 );
not \U$25060 ( \25403 , \25401 );
and \U$25061 ( \25404 , \25403 , \12619 );
nor \U$25062 ( \25405 , \25402 , \25404 );
and \U$25063 ( \25406 , \25398 , \25405 );
and \U$25064 ( \25407 , \25390 , \25397 );
or \U$25065 ( \25408 , \25406 , \25407 );
and \U$25066 ( \25409 , \25383 , \25408 );
and \U$25067 ( \25410 , \25356 , \25382 );
or \U$25068 ( \25411 , \25409 , \25410 );
xor \U$25069 ( \25412 , \25329 , \25411 );
xor \U$25070 ( \25413 , \25133 , \25141 );
xor \U$25071 ( \25414 , \25413 , \25150 );
nand \U$25072 ( \25415 , RI9870420_85, \2272 );
and \U$25073 ( \25416 , \25415 , \2030 );
not \U$25074 ( \25417 , \25415 );
and \U$25075 ( \25418 , \25417 , \2031 );
nor \U$25076 ( \25419 , \25416 , \25418 );
xor \U$25077 ( \25420 , \25414 , \25419 );
xor \U$25078 ( \25421 , \25004 , \25012 );
xor \U$25079 ( \25422 , \25421 , \25020 );
and \U$25080 ( \25423 , \25420 , \25422 );
and \U$25081 ( \25424 , \25414 , \25419 );
or \U$25082 ( \25425 , \25423 , \25424 );
and \U$25083 ( \25426 , \25412 , \25425 );
and \U$25084 ( \25427 , \25329 , \25411 );
or \U$25085 ( \25428 , \25426 , \25427 );
xor \U$25086 ( \25429 , \25248 , \25428 );
xor \U$25087 ( \25430 , \25031 , \25038 );
xor \U$25088 ( \25431 , \25430 , \25046 );
xor \U$25089 ( \25432 , \24979 , \24986 );
xor \U$25090 ( \25433 , \25432 , \24994 );
and \U$25091 ( \25434 , \25431 , \25433 );
xor \U$25092 ( \25435 , \25059 , \25066 );
xor \U$25093 ( \25436 , \25435 , \25074 );
xor \U$25094 ( \25437 , \24979 , \24986 );
xor \U$25095 ( \25438 , \25437 , \24994 );
and \U$25096 ( \25439 , \25436 , \25438 );
and \U$25097 ( \25440 , \25431 , \25436 );
or \U$25098 ( \25441 , \25434 , \25439 , \25440 );
xor \U$25099 ( \25442 , \25181 , \25183 );
xor \U$25100 ( \25443 , \25441 , \25442 );
xor \U$25101 ( \25444 , \24776 , \24783 );
xor \U$25102 ( \25445 , \25444 , \24791 );
xor \U$25103 ( \25446 , \25169 , \25174 );
xor \U$25104 ( \25447 , \25445 , \25446 );
and \U$25105 ( \25448 , \25443 , \25447 );
and \U$25106 ( \25449 , \25441 , \25442 );
or \U$25107 ( \25450 , \25448 , \25449 );
and \U$25108 ( \25451 , \25429 , \25450 );
and \U$25109 ( \25452 , \25248 , \25428 );
or \U$25110 ( \25453 , \25451 , \25452 );
xor \U$25111 ( \25454 , \24670 , \24672 );
xor \U$25112 ( \25455 , \25454 , \24685 );
xor \U$25113 ( \25456 , \25453 , \25455 );
xor \U$25114 ( \25457 , \24794 , \24820 );
xor \U$25115 ( \25458 , \25457 , \24846 );
xor \U$25116 ( \25459 , \25179 , \25184 );
xor \U$25117 ( \25460 , \25459 , \25189 );
and \U$25118 ( \25461 , \25458 , \25460 );
xor \U$25119 ( \25462 , \24876 , \24877 );
xor \U$25120 ( \25463 , \25462 , \24880 );
xor \U$25121 ( \25464 , \24960 , \24967 );
xor \U$25122 ( \25465 , \25463 , \25464 );
xor \U$25123 ( \25466 , \25179 , \25184 );
xor \U$25124 ( \25467 , \25466 , \25189 );
and \U$25125 ( \25468 , \25465 , \25467 );
and \U$25126 ( \25469 , \25458 , \25465 );
or \U$25127 ( \25470 , \25461 , \25468 , \25469 );
and \U$25128 ( \25471 , \25456 , \25470 );
and \U$25129 ( \25472 , \25453 , \25455 );
or \U$25130 ( \25473 , \25471 , \25472 );
and \U$25131 ( \25474 , \25236 , \25473 );
and \U$25132 ( \25475 , \25231 , \25235 );
or \U$25133 ( \25476 , \25474 , \25475 );
nand \U$25134 ( \25477 , \25219 , \25476 );
nand \U$25135 ( \25478 , \25218 , \25477 );
and \U$25136 ( \25479 , \25208 , \25478 );
xor \U$25137 ( \25480 , \25478 , \25208 );
xor \U$25138 ( \25481 , \25210 , \25212 );
xor \U$25139 ( \25482 , \25231 , \25235 );
xor \U$25140 ( \25483 , \25482 , \25473 );
xor \U$25141 ( \25484 , \25481 , \25483 );
xor \U$25142 ( \25485 , \25364 , \25371 );
xor \U$25143 ( \25486 , \25485 , \25379 );
not \U$25144 ( \25487 , \25343 );
not \U$25145 ( \25488 , \25354 );
or \U$25146 ( \25489 , \25487 , \25488 );
or \U$25147 ( \25490 , \25343 , \25354 );
nand \U$25148 ( \25491 , \25489 , \25490 );
not \U$25149 ( \25492 , \25491 );
not \U$25150 ( \25493 , \25336 );
and \U$25151 ( \25494 , \25492 , \25493 );
and \U$25152 ( \25495 , \25491 , \25336 );
nor \U$25153 ( \25496 , \25494 , \25495 );
or \U$25154 ( \25497 , \25486 , \25496 );
not \U$25155 ( \25498 , \25496 );
not \U$25156 ( \25499 , \25486 );
or \U$25157 ( \25500 , \25498 , \25499 );
xor \U$25158 ( \25501 , \25390 , \25397 );
xor \U$25159 ( \25502 , \25501 , \25405 );
nand \U$25160 ( \25503 , \25500 , \25502 );
nand \U$25161 ( \25504 , \25497 , \25503 );
xor \U$25162 ( \25505 , \25104 , \25111 );
xor \U$25163 ( \25506 , \25505 , \25119 );
xor \U$25164 ( \25507 , \25504 , \25506 );
xor \U$25165 ( \25508 , \25306 , \25314 );
xor \U$25166 ( \25509 , \25508 , \25323 );
xor \U$25167 ( \25510 , \25255 , \25262 );
xor \U$25168 ( \25511 , \25510 , \25270 );
or \U$25169 ( \25512 , \25509 , \25511 );
not \U$25170 ( \25513 , \25511 );
not \U$25171 ( \25514 , \25509 );
or \U$25172 ( \25515 , \25513 , \25514 );
xor \U$25173 ( \25516 , \25280 , \25287 );
xor \U$25174 ( \25517 , \25516 , \25295 );
nand \U$25175 ( \25518 , \25515 , \25517 );
nand \U$25176 ( \25519 , \25512 , \25518 );
and \U$25177 ( \25520 , \25507 , \25519 );
and \U$25178 ( \25521 , \25504 , \25506 );
or \U$25179 ( \25522 , \25520 , \25521 );
and \U$25180 ( \25523 , \5881 , RI986fca0_69);
and \U$25181 ( \25524 , RI986ff70_75, \5879 );
nor \U$25182 ( \25525 , \25523 , \25524 );
and \U$25183 ( \25526 , \25525 , \5885 );
not \U$25184 ( \25527 , \25525 );
and \U$25185 ( \25528 , \25527 , \5594 );
nor \U$25186 ( \25529 , \25526 , \25528 );
not \U$25187 ( \25530 , \25529 );
and \U$25188 ( \25531 , \6453 , RI986fe80_73);
and \U$25189 ( \25532 , RI9870060_77, \6451 );
nor \U$25190 ( \25533 , \25531 , \25532 );
and \U$25191 ( \25534 , \25533 , \6180 );
not \U$25192 ( \25535 , \25533 );
and \U$25193 ( \25536 , \25535 , \6190 );
nor \U$25194 ( \25537 , \25534 , \25536 );
not \U$25195 ( \25538 , \25537 );
and \U$25196 ( \25539 , \25530 , \25538 );
and \U$25197 ( \25540 , \25537 , \25529 );
and \U$25198 ( \25541 , \7079 , RI9870150_79);
and \U$25199 ( \25542 , RI9870f60_109, \7077 );
nor \U$25200 ( \25543 , \25541 , \25542 );
and \U$25201 ( \25544 , \25543 , \6709 );
not \U$25202 ( \25545 , \25543 );
and \U$25203 ( \25546 , \25545 , \6710 );
nor \U$25204 ( \25547 , \25544 , \25546 );
nor \U$25205 ( \25548 , \25540 , \25547 );
nor \U$25206 ( \25549 , \25539 , \25548 );
and \U$25207 ( \25550 , \4203 , RI9870600_89);
and \U$25208 ( \25551 , RI98708d0_95, \4201 );
nor \U$25209 ( \25552 , \25550 , \25551 );
and \U$25210 ( \25553 , \25552 , \3923 );
not \U$25211 ( \25554 , \25552 );
and \U$25212 ( \25555 , \25554 , \4207 );
nor \U$25213 ( \25556 , \25553 , \25555 );
not \U$25214 ( \25557 , \25556 );
and \U$25215 ( \25558 , \4710 , RI98707e0_93);
and \U$25216 ( \25559 , RI986fac0_65, \4708 );
nor \U$25217 ( \25560 , \25558 , \25559 );
not \U$25218 ( \25561 , \25560 );
not \U$25219 ( \25562 , \4521 );
and \U$25220 ( \25563 , \25561 , \25562 );
and \U$25221 ( \25564 , \25560 , \4521 );
nor \U$25222 ( \25565 , \25563 , \25564 );
not \U$25223 ( \25566 , \25565 );
and \U$25224 ( \25567 , \25557 , \25566 );
and \U$25225 ( \25568 , \25565 , \25556 );
and \U$25226 ( \25569 , \5318 , RI986fbb0_67);
and \U$25227 ( \25570 , RI986fd90_71, \5316 );
nor \U$25228 ( \25571 , \25569 , \25570 );
and \U$25229 ( \25572 , \25571 , \5322 );
not \U$25230 ( \25573 , \25571 );
and \U$25231 ( \25574 , \25573 , \5052 );
nor \U$25232 ( \25575 , \25572 , \25574 );
nor \U$25233 ( \25576 , \25568 , \25575 );
nor \U$25234 ( \25577 , \25567 , \25576 );
xor \U$25235 ( \25578 , \25549 , \25577 );
and \U$25236 ( \25579 , \7729 , RI9870ab0_99);
and \U$25237 ( \25580 , RI9870d80_105, \7727 );
nor \U$25238 ( \25581 , \25579 , \25580 );
and \U$25239 ( \25582 , \25581 , \7733 );
not \U$25240 ( \25583 , \25581 );
and \U$25241 ( \25584 , \25583 , \7480 );
nor \U$25242 ( \25585 , \25582 , \25584 );
not \U$25243 ( \25586 , \25585 );
and \U$25244 ( \25587 , \8486 , RI98709c0_97);
and \U$25245 ( \25588 , RI9870e70_107, \8484 );
nor \U$25246 ( \25589 , \25587 , \25588 );
and \U$25247 ( \25590 , \25589 , \8051 );
not \U$25248 ( \25591 , \25589 );
and \U$25249 ( \25592 , \25591 , \8050 );
nor \U$25250 ( \25593 , \25590 , \25592 );
not \U$25251 ( \25594 , \25593 );
and \U$25252 ( \25595 , \25586 , \25594 );
and \U$25253 ( \25596 , \25593 , \25585 );
and \U$25254 ( \25597 , \9237 , RI9870ba0_101);
and \U$25255 ( \25598 , RI9871050_111, \9235 );
nor \U$25256 ( \25599 , \25597 , \25598 );
and \U$25257 ( \25600 , \25599 , \8836 );
not \U$25258 ( \25601 , \25599 );
and \U$25259 ( \25602 , \25601 , \9241 );
nor \U$25260 ( \25603 , \25600 , \25602 );
nor \U$25261 ( \25604 , \25596 , \25603 );
nor \U$25262 ( \25605 , \25595 , \25604 );
and \U$25263 ( \25606 , \25578 , \25605 );
and \U$25264 ( \25607 , \25549 , \25577 );
or \U$25265 ( \25608 , \25606 , \25607 );
and \U$25266 ( \25609 , \3254 , RI9870330_83);
and \U$25267 ( \25610 , RI9870240_81, \3252 );
nor \U$25268 ( \25611 , \25609 , \25610 );
not \U$25269 ( \25612 , \25611 );
not \U$25270 ( \25613 , \3406 );
and \U$25271 ( \25614 , \25612 , \25613 );
and \U$25272 ( \25615 , \25611 , \3406 );
nor \U$25273 ( \25616 , \25614 , \25615 );
and \U$25274 ( \25617 , \2464 , RI9870420_85);
and \U$25275 ( \25618 , RI9870510_87, \2462 );
nor \U$25276 ( \25619 , \25617 , \25618 );
and \U$25277 ( \25620 , \25619 , \2263 );
not \U$25278 ( \25621 , \25619 );
and \U$25279 ( \25622 , \25621 , \2468 );
nor \U$25280 ( \25623 , \25620 , \25622 );
xor \U$25281 ( \25624 , \25616 , \25623 );
and \U$25282 ( \25625 , \3683 , RI9870240_81);
and \U$25283 ( \25626 , RI98706f0_91, \3681 );
nor \U$25284 ( \25627 , \25625 , \25626 );
not \U$25285 ( \25628 , \25627 );
not \U$25286 ( \25629 , \3412 );
and \U$25287 ( \25630 , \25628 , \25629 );
and \U$25288 ( \25631 , \25627 , \3412 );
nor \U$25289 ( \25632 , \25630 , \25631 );
not \U$25290 ( \25633 , \25632 );
nand \U$25291 ( \25634 , RI9870420_85, \2462 );
and \U$25292 ( \25635 , \25634 , \2263 );
not \U$25293 ( \25636 , \25634 );
and \U$25294 ( \25637 , \25636 , \2468 );
nor \U$25295 ( \25638 , \25635 , \25637 );
not \U$25296 ( \25639 , \25638 );
and \U$25297 ( \25640 , \25633 , \25639 );
and \U$25298 ( \25641 , \25632 , \25638 );
and \U$25299 ( \25642 , \3254 , RI9870510_87);
and \U$25300 ( \25643 , RI9870330_83, \3252 );
nor \U$25301 ( \25644 , \25642 , \25643 );
not \U$25302 ( \25645 , \25644 );
not \U$25303 ( \25646 , \3406 );
and \U$25304 ( \25647 , \25645 , \25646 );
and \U$25305 ( \25648 , \25644 , \2935 );
nor \U$25306 ( \25649 , \25647 , \25648 );
nor \U$25307 ( \25650 , \25641 , \25649 );
nor \U$25308 ( \25651 , \25640 , \25650 );
and \U$25309 ( \25652 , \25624 , \25651 );
and \U$25310 ( \25653 , \25616 , \25623 );
or \U$25311 ( \25654 , \25652 , \25653 );
or \U$25312 ( \25655 , \25608 , \25654 );
not \U$25313 ( \25656 , \25654 );
not \U$25314 ( \25657 , \25608 );
or \U$25315 ( \25658 , \25656 , \25657 );
and \U$25316 ( \25659 , \9505 , RI9870c90_103);
and \U$25317 ( \25660 , RI9871230_115, \9503 );
nor \U$25318 ( \25661 , \25659 , \25660 );
and \U$25319 ( \25662 , \25661 , \9513 );
not \U$25320 ( \25663 , \25661 );
and \U$25321 ( \25664 , \25663 , \9510 );
nor \U$25322 ( \25665 , \25662 , \25664 );
not \U$25323 ( \25666 , \25665 );
and \U$25324 ( \25667 , \10424 , RI9871140_113);
and \U$25325 ( \25668 , RI9871320_117, \10422 );
nor \U$25326 ( \25669 , \25667 , \25668 );
and \U$25327 ( \25670 , \25669 , \10428 );
not \U$25328 ( \25671 , \25669 );
and \U$25329 ( \25672 , \25671 , \9840 );
nor \U$25330 ( \25673 , \25670 , \25672 );
not \U$25331 ( \25674 , \25673 );
and \U$25332 ( \25675 , \25666 , \25674 );
and \U$25333 ( \25676 , \25673 , \25665 );
and \U$25334 ( \25677 , \11696 , RI9871410_119);
and \U$25335 ( \25678 , RI98716e0_125, \11694 );
nor \U$25336 ( \25679 , \25677 , \25678 );
and \U$25337 ( \25680 , \25679 , \11702 );
not \U$25338 ( \25681 , \25679 );
and \U$25339 ( \25682 , \25681 , \10965 );
nor \U$25340 ( \25683 , \25680 , \25682 );
nor \U$25341 ( \25684 , \25676 , \25683 );
nor \U$25342 ( \25685 , \25675 , \25684 );
and \U$25343 ( \25686 , \12293 , RI98717d0_127);
and \U$25344 ( \25687 , RI9871500_121, \12291 );
nor \U$25345 ( \25688 , \25686 , \25687 );
and \U$25346 ( \25689 , \25688 , \11686 );
not \U$25347 ( \25690 , \25688 );
and \U$25348 ( \25691 , \25690 , \11687 );
nor \U$25349 ( \25692 , \25689 , \25691 );
not \U$25350 ( \25693 , \25692 );
and \U$25351 ( \25694 , \13882 , RI986e9e0_29);
and \U$25352 ( \25695 , RI986e8f0_27, \13880 );
nor \U$25353 ( \25696 , \25694 , \25695 );
and \U$25354 ( \25697 , \25696 , \13359 );
not \U$25355 ( \25698 , \25696 );
and \U$25356 ( \25699 , \25698 , \13358 );
nor \U$25357 ( \25700 , \25697 , \25699 );
not \U$25358 ( \25701 , \25700 );
and \U$25359 ( \25702 , \25693 , \25701 );
and \U$25360 ( \25703 , \25700 , \25692 );
and \U$25361 ( \25704 , \13045 , RI98715f0_123);
and \U$25362 ( \25705 , RI986ead0_31, \13043 );
nor \U$25363 ( \25706 , \25704 , \25705 );
and \U$25364 ( \25707 , \25706 , \12619 );
not \U$25365 ( \25708 , \25706 );
and \U$25366 ( \25709 , \25708 , \13047 );
nor \U$25367 ( \25710 , \25707 , \25709 );
nor \U$25368 ( \25711 , \25703 , \25710 );
nor \U$25369 ( \25712 , \25702 , \25711 );
or \U$25370 ( \25713 , \25685 , \25712 );
not \U$25371 ( \25714 , \25685 );
not \U$25372 ( \25715 , \25712 );
or \U$25373 ( \25716 , \25714 , \25715 );
not \U$25374 ( \25717 , RI9873558_190);
and \U$25375 ( \25718 , \15780 , RI986eda0_37);
and \U$25376 ( \25719 , RI9873648_192, RI986ebc0_33);
nor \U$25377 ( \25720 , \25718 , \25719 );
not \U$25378 ( \25721 , \25720 );
or \U$25379 ( \25722 , \25717 , \25721 );
or \U$25380 ( \25723 , \25720 , RI9873558_190);
nand \U$25381 ( \25724 , \25722 , \25723 );
xor \U$25382 ( \25725 , \25724 , \2263 );
and \U$25383 ( \25726 , \14937 , RI986e800_25);
and \U$25384 ( \25727 , RI986ee90_39, \14935 );
nor \U$25385 ( \25728 , \25726 , \25727 );
and \U$25386 ( \25729 , \25728 , \14539 );
not \U$25387 ( \25730 , \25728 );
and \U$25388 ( \25731 , \25730 , \14538 );
nor \U$25389 ( \25732 , \25729 , \25731 );
and \U$25390 ( \25733 , \25725 , \25732 );
and \U$25391 ( \25734 , \25724 , \2263 );
or \U$25392 ( \25735 , \25733 , \25734 );
nand \U$25393 ( \25736 , \25716 , \25735 );
nand \U$25394 ( \25737 , \25713 , \25736 );
nand \U$25395 ( \25738 , \25658 , \25737 );
nand \U$25396 ( \25739 , \25655 , \25738 );
xor \U$25397 ( \25740 , \25522 , \25739 );
xor \U$25398 ( \25741 , \25085 , \2031 );
xor \U$25399 ( \25742 , \25741 , \25093 );
xor \U$25400 ( \25743 , \25414 , \25419 );
xor \U$25401 ( \25744 , \25743 , \25422 );
and \U$25402 ( \25745 , \25742 , \25744 );
xor \U$25403 ( \25746 , \24979 , \24986 );
xor \U$25404 ( \25747 , \25746 , \24994 );
xor \U$25405 ( \25748 , \25431 , \25436 );
xor \U$25406 ( \25749 , \25747 , \25748 );
xor \U$25407 ( \25750 , \25414 , \25419 );
xor \U$25408 ( \25751 , \25750 , \25422 );
and \U$25409 ( \25752 , \25749 , \25751 );
and \U$25410 ( \25753 , \25742 , \25749 );
or \U$25411 ( \25754 , \25745 , \25752 , \25753 );
and \U$25412 ( \25755 , \25740 , \25754 );
and \U$25413 ( \25756 , \25522 , \25739 );
or \U$25414 ( \25757 , \25755 , \25756 );
xor \U$25415 ( \25758 , \25052 , \25125 );
xor \U$25416 ( \25759 , \25758 , \25163 );
xor \U$25417 ( \25760 , \25757 , \25759 );
xor \U$25418 ( \25761 , \25329 , \25411 );
xor \U$25419 ( \25762 , \25761 , \25425 );
xor \U$25420 ( \25763 , \25238 , \25240 );
xor \U$25421 ( \25764 , \25763 , \25245 );
and \U$25422 ( \25765 , \25762 , \25764 );
xor \U$25423 ( \25766 , \25441 , \25442 );
xor \U$25424 ( \25767 , \25766 , \25447 );
xor \U$25425 ( \25768 , \25238 , \25240 );
xor \U$25426 ( \25769 , \25768 , \25245 );
and \U$25427 ( \25770 , \25767 , \25769 );
and \U$25428 ( \25771 , \25762 , \25767 );
or \U$25429 ( \25772 , \25765 , \25770 , \25771 );
and \U$25430 ( \25773 , \25760 , \25772 );
and \U$25431 ( \25774 , \25757 , \25759 );
or \U$25432 ( \25775 , \25773 , \25774 );
xor \U$25433 ( \25776 , \25248 , \25428 );
xor \U$25434 ( \25777 , \25776 , \25450 );
xor \U$25435 ( \25778 , \25179 , \25184 );
xor \U$25436 ( \25779 , \25778 , \25189 );
xor \U$25437 ( \25780 , \25458 , \25465 );
xor \U$25438 ( \25781 , \25779 , \25780 );
and \U$25439 ( \25782 , \25777 , \25781 );
xor \U$25440 ( \25783 , \25775 , \25782 );
xor \U$25441 ( \25784 , \24945 , \24947 );
xor \U$25442 ( \25785 , \25784 , \24952 );
xor \U$25443 ( \25786 , \25221 , \25226 );
xor \U$25444 ( \25787 , \25785 , \25786 );
and \U$25445 ( \25788 , \25783 , \25787 );
and \U$25446 ( \25789 , \25775 , \25782 );
or \U$25447 ( \25790 , \25788 , \25789 );
xor \U$25448 ( \25791 , \25484 , \25790 );
xor \U$25449 ( \25792 , \25453 , \25455 );
xor \U$25450 ( \25793 , \25792 , \25470 );
not \U$25451 ( \25794 , \25793 );
xor \U$25452 ( \25795 , \25775 , \25782 );
xor \U$25453 ( \25796 , \25795 , \25787 );
not \U$25454 ( \25797 , \25796 );
or \U$25455 ( \25798 , \25794 , \25797 );
or \U$25456 ( \25799 , \25796 , \25793 );
xor \U$25457 ( \25800 , \25777 , \25781 );
not \U$25458 ( \25801 , \25800 );
xor \U$25459 ( \25802 , \25757 , \25759 );
xor \U$25460 ( \25803 , \25802 , \25772 );
not \U$25461 ( \25804 , \25803 );
or \U$25462 ( \25805 , \25801 , \25804 );
or \U$25463 ( \25806 , \25803 , \25800 );
and \U$25464 ( \25807 , \7079 , RI9870060_77);
and \U$25465 ( \25808 , RI9870150_79, \7077 );
nor \U$25466 ( \25809 , \25807 , \25808 );
and \U$25467 ( \25810 , \25809 , \6709 );
not \U$25468 ( \25811 , \25809 );
and \U$25469 ( \25812 , \25811 , \6710 );
nor \U$25470 ( \25813 , \25810 , \25812 );
and \U$25471 ( \25814 , \8486 , RI9870d80_105);
and \U$25472 ( \25815 , RI98709c0_97, \8484 );
nor \U$25473 ( \25816 , \25814 , \25815 );
and \U$25474 ( \25817 , \25816 , \8051 );
not \U$25475 ( \25818 , \25816 );
and \U$25476 ( \25819 , \25818 , \8050 );
nor \U$25477 ( \25820 , \25817 , \25819 );
or \U$25478 ( \25821 , \25813 , \25820 );
not \U$25479 ( \25822 , \25820 );
not \U$25480 ( \25823 , \25813 );
or \U$25481 ( \25824 , \25822 , \25823 );
and \U$25482 ( \25825 , \7729 , RI9870f60_109);
and \U$25483 ( \25826 , RI9870ab0_99, \7727 );
nor \U$25484 ( \25827 , \25825 , \25826 );
and \U$25485 ( \25828 , \25827 , \7480 );
not \U$25486 ( \25829 , \25827 );
and \U$25487 ( \25830 , \25829 , \7733 );
nor \U$25488 ( \25831 , \25828 , \25830 );
nand \U$25489 ( \25832 , \25824 , \25831 );
nand \U$25490 ( \25833 , \25821 , \25832 );
not \U$25491 ( \25834 , \4521 );
and \U$25492 ( \25835 , \4710 , RI98708d0_95);
and \U$25493 ( \25836 , RI98707e0_93, \4708 );
nor \U$25494 ( \25837 , \25835 , \25836 );
not \U$25495 ( \25838 , \25837 );
or \U$25496 ( \25839 , \25834 , \25838 );
or \U$25497 ( \25840 , \25837 , \4521 );
nand \U$25498 ( \25841 , \25839 , \25840 );
not \U$25499 ( \25842 , \3412 );
and \U$25500 ( \25843 , \3683 , RI9870330_83);
and \U$25501 ( \25844 , RI9870240_81, \3681 );
nor \U$25502 ( \25845 , \25843 , \25844 );
not \U$25503 ( \25846 , \25845 );
or \U$25504 ( \25847 , \25842 , \25846 );
or \U$25505 ( \25848 , \25845 , \3918 );
nand \U$25506 ( \25849 , \25847 , \25848 );
xor \U$25507 ( \25850 , \25841 , \25849 );
and \U$25508 ( \25851 , \4203 , RI98706f0_91);
and \U$25509 ( \25852 , RI9870600_89, \4201 );
nor \U$25510 ( \25853 , \25851 , \25852 );
and \U$25511 ( \25854 , \25853 , \4207 );
not \U$25512 ( \25855 , \25853 );
and \U$25513 ( \25856 , \25855 , \3922 );
nor \U$25514 ( \25857 , \25854 , \25856 );
and \U$25515 ( \25858 , \25850 , \25857 );
and \U$25516 ( \25859 , \25841 , \25849 );
or \U$25517 ( \25860 , \25858 , \25859 );
xor \U$25518 ( \25861 , \25833 , \25860 );
and \U$25519 ( \25862 , \5318 , RI986fac0_65);
and \U$25520 ( \25863 , RI986fbb0_67, \5316 );
nor \U$25521 ( \25864 , \25862 , \25863 );
and \U$25522 ( \25865 , \25864 , \5322 );
not \U$25523 ( \25866 , \25864 );
and \U$25524 ( \25867 , \25866 , \5052 );
nor \U$25525 ( \25868 , \25865 , \25867 );
and \U$25526 ( \25869 , \6453 , RI986ff70_75);
and \U$25527 ( \25870 , RI986fe80_73, \6451 );
nor \U$25528 ( \25871 , \25869 , \25870 );
and \U$25529 ( \25872 , \25871 , \6180 );
not \U$25530 ( \25873 , \25871 );
and \U$25531 ( \25874 , \25873 , \6190 );
nor \U$25532 ( \25875 , \25872 , \25874 );
or \U$25533 ( \25876 , \25868 , \25875 );
not \U$25534 ( \25877 , \25875 );
not \U$25535 ( \25878 , \25868 );
or \U$25536 ( \25879 , \25877 , \25878 );
and \U$25537 ( \25880 , \5881 , RI986fd90_71);
and \U$25538 ( \25881 , RI986fca0_69, \5879 );
nor \U$25539 ( \25882 , \25880 , \25881 );
and \U$25540 ( \25883 , \25882 , \5594 );
not \U$25541 ( \25884 , \25882 );
and \U$25542 ( \25885 , \25884 , \5885 );
nor \U$25543 ( \25886 , \25883 , \25885 );
nand \U$25544 ( \25887 , \25879 , \25886 );
nand \U$25545 ( \25888 , \25876 , \25887 );
and \U$25546 ( \25889 , \25861 , \25888 );
and \U$25547 ( \25890 , \25833 , \25860 );
or \U$25548 ( \25891 , \25889 , \25890 );
and \U$25549 ( \25892 , \9505 , RI9871050_111);
and \U$25550 ( \25893 , RI9870c90_103, \9503 );
nor \U$25551 ( \25894 , \25892 , \25893 );
and \U$25552 ( \25895 , \25894 , \9513 );
not \U$25553 ( \25896 , \25894 );
and \U$25554 ( \25897 , \25896 , \9510 );
nor \U$25555 ( \25898 , \25895 , \25897 );
and \U$25556 ( \25899 , \10424 , RI9871230_115);
and \U$25557 ( \25900 , RI9871140_113, \10422 );
nor \U$25558 ( \25901 , \25899 , \25900 );
and \U$25559 ( \25902 , \25901 , \10428 );
not \U$25560 ( \25903 , \25901 );
and \U$25561 ( \25904 , \25903 , \9840 );
nor \U$25562 ( \25905 , \25902 , \25904 );
xor \U$25563 ( \25906 , \25898 , \25905 );
and \U$25564 ( \25907 , \9237 , RI9870e70_107);
and \U$25565 ( \25908 , RI9870ba0_101, \9235 );
nor \U$25566 ( \25909 , \25907 , \25908 );
and \U$25567 ( \25910 , \25909 , \8836 );
not \U$25568 ( \25911 , \25909 );
and \U$25569 ( \25912 , \25911 , \9241 );
nor \U$25570 ( \25913 , \25910 , \25912 );
and \U$25571 ( \25914 , \25906 , \25913 );
and \U$25572 ( \25915 , \25898 , \25905 );
nor \U$25573 ( \25916 , \25914 , \25915 );
and \U$25574 ( \25917 , \13882 , RI986ead0_31);
and \U$25575 ( \25918 , RI986e9e0_29, \13880 );
nor \U$25576 ( \25919 , \25917 , \25918 );
and \U$25577 ( \25920 , \25919 , \13359 );
not \U$25578 ( \25921 , \25919 );
and \U$25579 ( \25922 , \25921 , \13358 );
nor \U$25580 ( \25923 , \25920 , \25922 );
and \U$25581 ( \25924 , \15780 , RI986ee90_39);
and \U$25582 ( \25925 , RI9873648_192, RI986eda0_37);
nor \U$25583 ( \25926 , \25924 , \25925 );
not \U$25584 ( \25927 , \25926 );
not \U$25585 ( \25928 , RI9873558_190);
and \U$25586 ( \25929 , \25927 , \25928 );
and \U$25587 ( \25930 , \25926 , RI9873558_190);
nor \U$25588 ( \25931 , \25929 , \25930 );
or \U$25589 ( \25932 , \25923 , \25931 );
not \U$25590 ( \25933 , \25931 );
not \U$25591 ( \25934 , \25923 );
or \U$25592 ( \25935 , \25933 , \25934 );
and \U$25593 ( \25936 , \14937 , RI986e8f0_27);
and \U$25594 ( \25937 , RI986e800_25, \14935 );
nor \U$25595 ( \25938 , \25936 , \25937 );
and \U$25596 ( \25939 , \25938 , \14539 );
not \U$25597 ( \25940 , \25938 );
and \U$25598 ( \25941 , \25940 , \14538 );
nor \U$25599 ( \25942 , \25939 , \25941 );
nand \U$25600 ( \25943 , \25935 , \25942 );
nand \U$25601 ( \25944 , \25932 , \25943 );
xor \U$25602 ( \25945 , \25916 , \25944 );
and \U$25603 ( \25946 , \11696 , RI9871320_117);
and \U$25604 ( \25947 , RI9871410_119, \11694 );
nor \U$25605 ( \25948 , \25946 , \25947 );
and \U$25606 ( \25949 , \25948 , \11702 );
not \U$25607 ( \25950 , \25948 );
and \U$25608 ( \25951 , \25950 , \10965 );
nor \U$25609 ( \25952 , \25949 , \25951 );
and \U$25610 ( \25953 , \13045 , RI9871500_121);
and \U$25611 ( \25954 , RI98715f0_123, \13043 );
nor \U$25612 ( \25955 , \25953 , \25954 );
and \U$25613 ( \25956 , \25955 , \12619 );
not \U$25614 ( \25957 , \25955 );
and \U$25615 ( \25958 , \25957 , \13047 );
nor \U$25616 ( \25959 , \25956 , \25958 );
or \U$25617 ( \25960 , \25952 , \25959 );
not \U$25618 ( \25961 , \25959 );
not \U$25619 ( \25962 , \25952 );
or \U$25620 ( \25963 , \25961 , \25962 );
and \U$25621 ( \25964 , \12293 , RI98716e0_125);
and \U$25622 ( \25965 , RI98717d0_127, \12291 );
nor \U$25623 ( \25966 , \25964 , \25965 );
and \U$25624 ( \25967 , \25966 , \11687 );
not \U$25625 ( \25968 , \25966 );
and \U$25626 ( \25969 , \25968 , \11686 );
nor \U$25627 ( \25970 , \25967 , \25969 );
nand \U$25628 ( \25971 , \25963 , \25970 );
nand \U$25629 ( \25972 , \25960 , \25971 );
and \U$25630 ( \25973 , \25945 , \25972 );
and \U$25631 ( \25974 , \25916 , \25944 );
or \U$25632 ( \25975 , \25973 , \25974 );
xor \U$25633 ( \25976 , \25891 , \25975 );
not \U$25634 ( \25977 , \25638 );
xor \U$25635 ( \25978 , \25649 , \25632 );
not \U$25636 ( \25979 , \25978 );
or \U$25637 ( \25980 , \25977 , \25979 );
or \U$25638 ( \25981 , \25978 , \25638 );
nand \U$25639 ( \25982 , \25980 , \25981 );
not \U$25640 ( \25983 , \25556 );
xor \U$25641 ( \25984 , \25565 , \25575 );
not \U$25642 ( \25985 , \25984 );
or \U$25643 ( \25986 , \25983 , \25985 );
or \U$25644 ( \25987 , \25984 , \25556 );
nand \U$25645 ( \25988 , \25986 , \25987 );
xor \U$25646 ( \25989 , \25982 , \25988 );
not \U$25647 ( \25990 , \25529 );
xor \U$25648 ( \25991 , \25537 , \25547 );
not \U$25649 ( \25992 , \25991 );
or \U$25650 ( \25993 , \25990 , \25992 );
or \U$25651 ( \25994 , \25991 , \25529 );
nand \U$25652 ( \25995 , \25993 , \25994 );
and \U$25653 ( \25996 , \25989 , \25995 );
and \U$25654 ( \25997 , \25982 , \25988 );
or \U$25655 ( \25998 , \25996 , \25997 );
and \U$25656 ( \25999 , \25976 , \25998 );
and \U$25657 ( \26000 , \25891 , \25975 );
nor \U$25658 ( \26001 , \25999 , \26000 );
xor \U$25659 ( \26002 , \25549 , \25577 );
xor \U$25660 ( \26003 , \26002 , \25605 );
not \U$25661 ( \26004 , \26003 );
not \U$25662 ( \26005 , \25735 );
not \U$25663 ( \26006 , \25685 );
or \U$25664 ( \26007 , \26005 , \26006 );
or \U$25665 ( \26008 , \25685 , \25735 );
nand \U$25666 ( \26009 , \26007 , \26008 );
not \U$25667 ( \26010 , \26009 );
not \U$25668 ( \26011 , \25712 );
and \U$25669 ( \26012 , \26010 , \26011 );
and \U$25670 ( \26013 , \26009 , \25712 );
nor \U$25671 ( \26014 , \26012 , \26013 );
not \U$25672 ( \26015 , \26014 );
and \U$25673 ( \26016 , \26004 , \26015 );
and \U$25674 ( \26017 , \26003 , \26014 );
xor \U$25675 ( \26018 , \25616 , \25623 );
xor \U$25676 ( \26019 , \26018 , \25651 );
nor \U$25677 ( \26020 , \26017 , \26019 );
nor \U$25678 ( \26021 , \26016 , \26020 );
xor \U$25679 ( \26022 , \26001 , \26021 );
not \U$25680 ( \26023 , \25502 );
not \U$25681 ( \26024 , \25486 );
or \U$25682 ( \26025 , \26023 , \26024 );
or \U$25683 ( \26026 , \25486 , \25502 );
nand \U$25684 ( \26027 , \26025 , \26026 );
not \U$25685 ( \26028 , \26027 );
not \U$25686 ( \26029 , \25496 );
and \U$25687 ( \26030 , \26028 , \26029 );
and \U$25688 ( \26031 , \26027 , \25496 );
nor \U$25689 ( \26032 , \26030 , \26031 );
not \U$25690 ( \26033 , \26032 );
not \U$25691 ( \26034 , \25511 );
not \U$25692 ( \26035 , \25517 );
or \U$25693 ( \26036 , \26034 , \26035 );
or \U$25694 ( \26037 , \25511 , \25517 );
nand \U$25695 ( \26038 , \26036 , \26037 );
not \U$25696 ( \26039 , \26038 );
not \U$25697 ( \26040 , \25509 );
and \U$25698 ( \26041 , \26039 , \26040 );
and \U$25699 ( \26042 , \26038 , \25509 );
nor \U$25700 ( \26043 , \26041 , \26042 );
not \U$25701 ( \26044 , \26043 );
and \U$25702 ( \26045 , \26033 , \26044 );
and \U$25703 ( \26046 , \26032 , \26043 );
not \U$25704 ( \26047 , \25585 );
xor \U$25705 ( \26048 , \25593 , \25603 );
not \U$25706 ( \26049 , \26048 );
or \U$25707 ( \26050 , \26047 , \26049 );
or \U$25708 ( \26051 , \26048 , \25585 );
nand \U$25709 ( \26052 , \26050 , \26051 );
not \U$25710 ( \26053 , \25665 );
xor \U$25711 ( \26054 , \25673 , \25683 );
not \U$25712 ( \26055 , \26054 );
or \U$25713 ( \26056 , \26053 , \26055 );
or \U$25714 ( \26057 , \26054 , \25665 );
nand \U$25715 ( \26058 , \26056 , \26057 );
xor \U$25716 ( \26059 , \26052 , \26058 );
not \U$25717 ( \26060 , \25692 );
xor \U$25718 ( \26061 , \25710 , \25700 );
not \U$25719 ( \26062 , \26061 );
or \U$25720 ( \26063 , \26060 , \26062 );
or \U$25721 ( \26064 , \26061 , \25692 );
nand \U$25722 ( \26065 , \26063 , \26064 );
and \U$25723 ( \26066 , \26059 , \26065 );
and \U$25724 ( \26067 , \26052 , \26058 );
nor \U$25725 ( \26068 , \26066 , \26067 );
nor \U$25726 ( \26069 , \26046 , \26068 );
nor \U$25727 ( \26070 , \26045 , \26069 );
and \U$25728 ( \26071 , \26022 , \26070 );
and \U$25729 ( \26072 , \26001 , \26021 );
nor \U$25730 ( \26073 , \26071 , \26072 );
xor \U$25731 ( \26074 , \25356 , \25382 );
xor \U$25732 ( \26075 , \26074 , \25408 );
xor \U$25733 ( \26076 , \25273 , \25298 );
xor \U$25734 ( \26077 , \26076 , \25326 );
and \U$25735 ( \26078 , \26075 , \26077 );
xor \U$25736 ( \26079 , \25414 , \25419 );
xor \U$25737 ( \26080 , \26079 , \25422 );
xor \U$25738 ( \26081 , \25742 , \25749 );
xor \U$25739 ( \26082 , \26080 , \26081 );
xor \U$25740 ( \26083 , \25273 , \25298 );
xor \U$25741 ( \26084 , \26083 , \25326 );
and \U$25742 ( \26085 , \26082 , \26084 );
and \U$25743 ( \26086 , \26075 , \26082 );
or \U$25744 ( \26087 , \26078 , \26085 , \26086 );
xor \U$25745 ( \26088 , \26073 , \26087 );
xor \U$25746 ( \26089 , \25238 , \25240 );
xor \U$25747 ( \26090 , \26089 , \25245 );
xor \U$25748 ( \26091 , \25762 , \25767 );
xor \U$25749 ( \26092 , \26090 , \26091 );
and \U$25750 ( \26093 , \26088 , \26092 );
and \U$25751 ( \26094 , \26073 , \26087 );
or \U$25752 ( \26095 , \26093 , \26094 );
nand \U$25753 ( \26096 , \25806 , \26095 );
nand \U$25754 ( \26097 , \25805 , \26096 );
nand \U$25755 ( \26098 , \25799 , \26097 );
nand \U$25756 ( \26099 , \25798 , \26098 );
and \U$25757 ( \26100 , \25791 , \26099 );
xor \U$25758 ( \26101 , \26099 , \25791 );
and \U$25759 ( \26102 , \15780 , RI98715f0_123);
and \U$25760 ( \26103 , RI9873648_192, RI986ead0_31);
nor \U$25761 ( \26104 , \26102 , \26103 );
not \U$25762 ( \26105 , \26104 );
not \U$25763 ( \26106 , RI9873558_190);
and \U$25764 ( \26107 , \26105 , \26106 );
and \U$25765 ( \26108 , \26104 , RI9873558_190);
nor \U$25766 ( \26109 , \26107 , \26108 );
xor \U$25767 ( \26110 , \26109 , \4207 );
and \U$25768 ( \26111 , \14937 , RI98717d0_127);
and \U$25769 ( \26112 , RI9871500_121, \14935 );
nor \U$25770 ( \26113 , \26111 , \26112 );
and \U$25771 ( \26114 , \26113 , \14538 );
not \U$25772 ( \26115 , \26113 );
and \U$25773 ( \26116 , \26115 , \14539 );
nor \U$25774 ( \26117 , \26114 , \26116 );
xor \U$25775 ( \26118 , \26110 , \26117 );
and \U$25776 ( \26119 , \13882 , RI9871410_119);
and \U$25777 ( \26120 , RI98716e0_125, \13880 );
nor \U$25778 ( \26121 , \26119 , \26120 );
and \U$25779 ( \26122 , \26121 , \13359 );
not \U$25780 ( \26123 , \26121 );
and \U$25781 ( \26124 , \26123 , \13358 );
nor \U$25782 ( \26125 , \26122 , \26124 );
and \U$25783 ( \26126 , \12293 , RI9870c90_103);
and \U$25784 ( \26127 , RI9871230_115, \12291 );
nor \U$25785 ( \26128 , \26126 , \26127 );
and \U$25786 ( \26129 , \26128 , \11686 );
not \U$25787 ( \26130 , \26128 );
and \U$25788 ( \26131 , \26130 , \11687 );
nor \U$25789 ( \26132 , \26129 , \26131 );
xor \U$25790 ( \26133 , \26125 , \26132 );
and \U$25791 ( \26134 , \13045 , RI9871140_113);
and \U$25792 ( \26135 , RI9871320_117, \13043 );
nor \U$25793 ( \26136 , \26134 , \26135 );
and \U$25794 ( \26137 , \26136 , \12619 );
not \U$25795 ( \26138 , \26136 );
and \U$25796 ( \26139 , \26138 , \13047 );
nor \U$25797 ( \26140 , \26137 , \26139 );
xor \U$25798 ( \26141 , \26133 , \26140 );
or \U$25799 ( \26142 , \26118 , \26141 );
and \U$25800 ( \26143 , \26118 , \26141 );
and \U$25801 ( \26144 , \9237 , RI9870150_79);
and \U$25802 ( \26145 , RI9870f60_109, \9235 );
nor \U$25803 ( \26146 , \26144 , \26145 );
and \U$25804 ( \26147 , \26146 , \8836 );
not \U$25805 ( \26148 , \26146 );
and \U$25806 ( \26149 , \26148 , \9241 );
nor \U$25807 ( \26150 , \26147 , \26149 );
and \U$25808 ( \26151 , \7729 , RI986fca0_69);
and \U$25809 ( \26152 , RI986ff70_75, \7727 );
nor \U$25810 ( \26153 , \26151 , \26152 );
and \U$25811 ( \26154 , \26153 , \7733 );
not \U$25812 ( \26155 , \26153 );
and \U$25813 ( \26156 , \26155 , \7480 );
nor \U$25814 ( \26157 , \26154 , \26156 );
xor \U$25815 ( \26158 , \26150 , \26157 );
and \U$25816 ( \26159 , \8486 , RI986fe80_73);
and \U$25817 ( \26160 , RI9870060_77, \8484 );
nor \U$25818 ( \26161 , \26159 , \26160 );
and \U$25819 ( \26162 , \26161 , \8051 );
not \U$25820 ( \26163 , \26161 );
and \U$25821 ( \26164 , \26163 , \8050 );
nor \U$25822 ( \26165 , \26162 , \26164 );
xor \U$25823 ( \26166 , \26158 , \26165 );
and \U$25824 ( \26167 , \7079 , RI986fbb0_67);
and \U$25825 ( \26168 , RI986fd90_71, \7077 );
nor \U$25826 ( \26169 , \26167 , \26168 );
and \U$25827 ( \26170 , \26169 , \6709 );
not \U$25828 ( \26171 , \26169 );
and \U$25829 ( \26172 , \26171 , \6710 );
nor \U$25830 ( \26173 , \26170 , \26172 );
and \U$25831 ( \26174 , \5881 , RI9870600_89);
and \U$25832 ( \26175 , RI98708d0_95, \5879 );
nor \U$25833 ( \26176 , \26174 , \26175 );
and \U$25834 ( \26177 , \26176 , \5885 );
not \U$25835 ( \26178 , \26176 );
and \U$25836 ( \26179 , \26178 , \5594 );
nor \U$25837 ( \26180 , \26177 , \26179 );
xor \U$25838 ( \26181 , \26173 , \26180 );
and \U$25839 ( \26182 , \6453 , RI98707e0_93);
and \U$25840 ( \26183 , RI986fac0_65, \6451 );
nor \U$25841 ( \26184 , \26182 , \26183 );
and \U$25842 ( \26185 , \26184 , \6705 );
not \U$25843 ( \26186 , \26184 );
and \U$25844 ( \26187 , \26186 , \6190 );
nor \U$25845 ( \26188 , \26185 , \26187 );
xor \U$25846 ( \26189 , \26181 , \26188 );
and \U$25847 ( \26190 , \10424 , RI98709c0_97);
and \U$25848 ( \26191 , RI9870e70_107, \10422 );
nor \U$25849 ( \26192 , \26190 , \26191 );
and \U$25850 ( \26193 , \26192 , \10428 );
not \U$25851 ( \26194 , \26192 );
and \U$25852 ( \26195 , \26194 , \9840 );
nor \U$25853 ( \26196 , \26193 , \26195 );
and \U$25854 ( \26197 , \9505 , RI9870ab0_99);
and \U$25855 ( \26198 , RI9870d80_105, \9503 );
nor \U$25856 ( \26199 , \26197 , \26198 );
and \U$25857 ( \26200 , \26199 , \9513 );
not \U$25858 ( \26201 , \26199 );
and \U$25859 ( \26202 , \26201 , \9510 );
nor \U$25860 ( \26203 , \26200 , \26202 );
xor \U$25861 ( \26204 , \26196 , \26203 );
and \U$25862 ( \26205 , \11696 , RI9870ba0_101);
and \U$25863 ( \26206 , RI9871050_111, \11694 );
nor \U$25864 ( \26207 , \26205 , \26206 );
and \U$25865 ( \26208 , \26207 , \11702 );
not \U$25866 ( \26209 , \26207 );
and \U$25867 ( \26210 , \26209 , \10965 );
nor \U$25868 ( \26211 , \26208 , \26210 );
xor \U$25869 ( \26212 , \26204 , \26211 );
xor \U$25870 ( \26213 , \26189 , \26212 );
xor \U$25871 ( \26214 , \26166 , \26213 );
nor \U$25872 ( \26215 , \26143 , \26214 );
not \U$25873 ( \26216 , \26215 );
nand \U$25874 ( \26217 , \26142 , \26216 );
not \U$25875 ( \26218 , \26217 );
and \U$25876 ( \26219 , \13882 , RI9871140_113);
and \U$25877 ( \26220 , RI9871320_117, \13880 );
nor \U$25878 ( \26221 , \26219 , \26220 );
and \U$25879 ( \26222 , \26221 , \13358 );
not \U$25880 ( \26223 , \26221 );
and \U$25881 ( \26224 , \26223 , \13359 );
nor \U$25882 ( \26225 , \26222 , \26224 );
and \U$25883 ( \26226 , \12293 , RI9870ba0_101);
and \U$25884 ( \26227 , RI9871050_111, \12291 );
nor \U$25885 ( \26228 , \26226 , \26227 );
and \U$25886 ( \26229 , \26228 , \11687 );
not \U$25887 ( \26230 , \26228 );
and \U$25888 ( \26231 , \26230 , \11686 );
nor \U$25889 ( \26232 , \26229 , \26231 );
xor \U$25890 ( \26233 , \26225 , \26232 );
and \U$25891 ( \26234 , \13045 , RI9870c90_103);
and \U$25892 ( \26235 , RI9871230_115, \13043 );
nor \U$25893 ( \26236 , \26234 , \26235 );
and \U$25894 ( \26237 , \26236 , \13047 );
not \U$25895 ( \26238 , \26236 );
and \U$25896 ( \26239 , \26238 , \12619 );
nor \U$25897 ( \26240 , \26237 , \26239 );
and \U$25898 ( \26241 , \26233 , \26240 );
and \U$25899 ( \26242 , \26225 , \26232 );
or \U$25900 ( \26243 , \26241 , \26242 );
not \U$25901 ( \26244 , RI9873558_190);
and \U$25902 ( \26245 , \15780 , RI98717d0_127);
and \U$25903 ( \26246 , RI9873648_192, RI9871500_121);
nor \U$25904 ( \26247 , \26245 , \26246 );
not \U$25905 ( \26248 , \26247 );
or \U$25906 ( \26249 , \26244 , \26248 );
or \U$25907 ( \26250 , \26247 , RI9873558_190);
nand \U$25908 ( \26251 , \26249 , \26250 );
xor \U$25909 ( \26252 , \26251 , \4521 );
and \U$25910 ( \26253 , \14937 , RI9871410_119);
and \U$25911 ( \26254 , RI98716e0_125, \14935 );
nor \U$25912 ( \26255 , \26253 , \26254 );
and \U$25913 ( \26256 , \26255 , \14539 );
not \U$25914 ( \26257 , \26255 );
and \U$25915 ( \26258 , \26257 , \14538 );
nor \U$25916 ( \26259 , \26256 , \26258 );
and \U$25917 ( \26260 , \26252 , \26259 );
and \U$25918 ( \26261 , \26251 , \4521 );
or \U$25919 ( \26262 , \26260 , \26261 );
and \U$25920 ( \26263 , \26243 , \26262 );
not \U$25921 ( \26264 , \26243 );
not \U$25922 ( \26265 , \26262 );
and \U$25923 ( \26266 , \26264 , \26265 );
and \U$25924 ( \26267 , \10424 , RI9870ab0_99);
and \U$25925 ( \26268 , RI9870d80_105, \10422 );
nor \U$25926 ( \26269 , \26267 , \26268 );
and \U$25927 ( \26270 , \26269 , \9840 );
not \U$25928 ( \26271 , \26269 );
and \U$25929 ( \26272 , \26271 , \10428 );
nor \U$25930 ( \26273 , \26270 , \26272 );
and \U$25931 ( \26274 , \11696 , RI98709c0_97);
and \U$25932 ( \26275 , RI9870e70_107, \11694 );
nor \U$25933 ( \26276 , \26274 , \26275 );
and \U$25934 ( \26277 , \26276 , \10965 );
not \U$25935 ( \26278 , \26276 );
and \U$25936 ( \26279 , \26278 , \11702 );
nor \U$25937 ( \26280 , \26277 , \26279 );
xor \U$25938 ( \26281 , \26273 , \26280 );
and \U$25939 ( \26282 , \9505 , RI9870150_79);
and \U$25940 ( \26283 , RI9870f60_109, \9503 );
nor \U$25941 ( \26284 , \26282 , \26283 );
and \U$25942 ( \26285 , \26284 , \9510 );
not \U$25943 ( \26286 , \26284 );
and \U$25944 ( \26287 , \26286 , \9513 );
nor \U$25945 ( \26288 , \26285 , \26287 );
and \U$25946 ( \26289 , \26281 , \26288 );
and \U$25947 ( \26290 , \26273 , \26280 );
nor \U$25948 ( \26291 , \26289 , \26290 );
nor \U$25949 ( \26292 , \26266 , \26291 );
nor \U$25950 ( \26293 , \26263 , \26292 );
and \U$25951 ( \26294 , \6453 , RI9870600_89);
and \U$25952 ( \26295 , RI98708d0_95, \6451 );
nor \U$25953 ( \26296 , \26294 , \26295 );
and \U$25954 ( \26297 , \26296 , \6190 );
not \U$25955 ( \26298 , \26296 );
and \U$25956 ( \26299 , \26298 , \6180 );
nor \U$25957 ( \26300 , \26297 , \26299 );
and \U$25958 ( \26301 , \7079 , RI98707e0_93);
and \U$25959 ( \26302 , RI986fac0_65, \7077 );
nor \U$25960 ( \26303 , \26301 , \26302 );
and \U$25961 ( \26304 , \26303 , \6710 );
not \U$25962 ( \26305 , \26303 );
and \U$25963 ( \26306 , \26305 , \6709 );
nor \U$25964 ( \26307 , \26304 , \26306 );
xor \U$25965 ( \26308 , \26300 , \26307 );
and \U$25966 ( \26309 , \5881 , RI9870240_81);
and \U$25967 ( \26310 , RI98706f0_91, \5879 );
nor \U$25968 ( \26311 , \26309 , \26310 );
and \U$25969 ( \26312 , \26311 , \5594 );
not \U$25970 ( \26313 , \26311 );
and \U$25971 ( \26314 , \26313 , \5885 );
nor \U$25972 ( \26315 , \26312 , \26314 );
and \U$25973 ( \26316 , \26308 , \26315 );
and \U$25974 ( \26317 , \26300 , \26307 );
nor \U$25975 ( \26318 , \26316 , \26317 );
not \U$25976 ( \26319 , \26318 );
and \U$25977 ( \26320 , \4710 , RI9870420_85);
and \U$25978 ( \26321 , RI9870510_87, \4708 );
nor \U$25979 ( \26322 , \26320 , \26321 );
not \U$25980 ( \26323 , \26322 );
not \U$25981 ( \26324 , \4521 );
and \U$25982 ( \26325 , \26323 , \26324 );
and \U$25983 ( \26326 , \26322 , \4519 );
nor \U$25984 ( \26327 , \26325 , \26326 );
not \U$25985 ( \26328 , \26327 );
and \U$25986 ( \26329 , \26319 , \26328 );
and \U$25987 ( \26330 , \26318 , \26327 );
and \U$25988 ( \26331 , \8486 , RI986fca0_69);
and \U$25989 ( \26332 , RI986ff70_75, \8484 );
nor \U$25990 ( \26333 , \26331 , \26332 );
and \U$25991 ( \26334 , \26333 , \8050 );
not \U$25992 ( \26335 , \26333 );
and \U$25993 ( \26336 , \26335 , \8051 );
nor \U$25994 ( \26337 , \26334 , \26336 );
and \U$25995 ( \26338 , \9237 , RI986fe80_73);
and \U$25996 ( \26339 , RI9870060_77, \9235 );
nor \U$25997 ( \26340 , \26338 , \26339 );
and \U$25998 ( \26341 , \26340 , \9241 );
not \U$25999 ( \26342 , \26340 );
and \U$26000 ( \26343 , \26342 , \8836 );
nor \U$26001 ( \26344 , \26341 , \26343 );
xor \U$26002 ( \26345 , \26337 , \26344 );
and \U$26003 ( \26346 , \7729 , RI986fbb0_67);
and \U$26004 ( \26347 , RI986fd90_71, \7727 );
nor \U$26005 ( \26348 , \26346 , \26347 );
and \U$26006 ( \26349 , \26348 , \7480 );
not \U$26007 ( \26350 , \26348 );
and \U$26008 ( \26351 , \26350 , \7733 );
nor \U$26009 ( \26352 , \26349 , \26351 );
and \U$26010 ( \26353 , \26345 , \26352 );
and \U$26011 ( \26354 , \26337 , \26344 );
nor \U$26012 ( \26355 , \26353 , \26354 );
nor \U$26013 ( \26356 , \26330 , \26355 );
nor \U$26014 ( \26357 , \26329 , \26356 );
xor \U$26015 ( \26358 , \26293 , \26357 );
and \U$26016 ( \26359 , \5318 , RI9870330_83);
and \U$26017 ( \26360 , RI9870240_81, \5316 );
nor \U$26018 ( \26361 , \26359 , \26360 );
and \U$26019 ( \26362 , \26361 , \5322 );
not \U$26020 ( \26363 , \26361 );
and \U$26021 ( \26364 , \26363 , \5052 );
nor \U$26022 ( \26365 , \26362 , \26364 );
not \U$26023 ( \26366 , \26365 );
and \U$26024 ( \26367 , \5881 , RI98706f0_91);
and \U$26025 ( \26368 , RI9870600_89, \5879 );
nor \U$26026 ( \26369 , \26367 , \26368 );
and \U$26027 ( \26370 , \26369 , \5885 );
not \U$26028 ( \26371 , \26369 );
and \U$26029 ( \26372 , \26371 , \5594 );
nor \U$26030 ( \26373 , \26370 , \26372 );
and \U$26031 ( \26374 , \6453 , RI98708d0_95);
and \U$26032 ( \26375 , RI98707e0_93, \6451 );
nor \U$26033 ( \26376 , \26374 , \26375 );
and \U$26034 ( \26377 , \26376 , \6180 );
not \U$26035 ( \26378 , \26376 );
and \U$26036 ( \26379 , \26378 , \6190 );
nor \U$26037 ( \26380 , \26377 , \26379 );
xor \U$26038 ( \26381 , \26373 , \26380 );
not \U$26039 ( \26382 , \26381 );
or \U$26040 ( \26383 , \26366 , \26382 );
or \U$26041 ( \26384 , \26381 , \26365 );
nand \U$26042 ( \26385 , \26383 , \26384 );
and \U$26043 ( \26386 , \7079 , RI986fac0_65);
and \U$26044 ( \26387 , RI986fbb0_67, \7077 );
nor \U$26045 ( \26388 , \26386 , \26387 );
and \U$26046 ( \26389 , \26388 , \6709 );
not \U$26047 ( \26390 , \26388 );
and \U$26048 ( \26391 , \26390 , \6710 );
nor \U$26049 ( \26392 , \26389 , \26391 );
not \U$26050 ( \26393 , \26392 );
and \U$26051 ( \26394 , \7729 , RI986fd90_71);
and \U$26052 ( \26395 , RI986fca0_69, \7727 );
nor \U$26053 ( \26396 , \26394 , \26395 );
and \U$26054 ( \26397 , \26396 , \7733 );
not \U$26055 ( \26398 , \26396 );
and \U$26056 ( \26399 , \26398 , \7480 );
nor \U$26057 ( \26400 , \26397 , \26399 );
and \U$26058 ( \26401 , \8486 , RI986ff70_75);
and \U$26059 ( \26402 , RI986fe80_73, \8484 );
nor \U$26060 ( \26403 , \26401 , \26402 );
and \U$26061 ( \26404 , \26403 , \8051 );
not \U$26062 ( \26405 , \26403 );
and \U$26063 ( \26406 , \26405 , \8050 );
nor \U$26064 ( \26407 , \26404 , \26406 );
xor \U$26065 ( \26408 , \26400 , \26407 );
not \U$26066 ( \26409 , \26408 );
or \U$26067 ( \26410 , \26393 , \26409 );
or \U$26068 ( \26411 , \26408 , \26392 );
nand \U$26069 ( \26412 , \26410 , \26411 );
xor \U$26070 ( \26413 , \26385 , \26412 );
and \U$26071 ( \26414 , \9505 , RI9870f60_109);
and \U$26072 ( \26415 , RI9870ab0_99, \9503 );
nor \U$26073 ( \26416 , \26414 , \26415 );
and \U$26074 ( \26417 , \26416 , \9510 );
not \U$26075 ( \26418 , \26416 );
and \U$26076 ( \26419 , \26418 , \9513 );
nor \U$26077 ( \26420 , \26417 , \26419 );
and \U$26078 ( \26421 , \9237 , RI9870060_77);
and \U$26079 ( \26422 , RI9870150_79, \9235 );
nor \U$26080 ( \26423 , \26421 , \26422 );
and \U$26081 ( \26424 , \26423 , \9241 );
not \U$26082 ( \26425 , \26423 );
and \U$26083 ( \26426 , \26425 , \8836 );
nor \U$26084 ( \26427 , \26424 , \26426 );
xor \U$26085 ( \26428 , \26420 , \26427 );
and \U$26086 ( \26429 , \10424 , RI9870d80_105);
and \U$26087 ( \26430 , RI98709c0_97, \10422 );
nor \U$26088 ( \26431 , \26429 , \26430 );
and \U$26089 ( \26432 , \26431 , \9840 );
not \U$26090 ( \26433 , \26431 );
and \U$26091 ( \26434 , \26433 , \10428 );
nor \U$26092 ( \26435 , \26432 , \26434 );
xor \U$26093 ( \26436 , \26428 , \26435 );
and \U$26094 ( \26437 , \26413 , \26436 );
and \U$26095 ( \26438 , \26385 , \26412 );
nor \U$26096 ( \26439 , \26437 , \26438 );
and \U$26097 ( \26440 , \26358 , \26439 );
and \U$26098 ( \26441 , \26293 , \26357 );
or \U$26099 ( \26442 , \26440 , \26441 );
not \U$26100 ( \26443 , \26442 );
or \U$26101 ( \26444 , \26218 , \26443 );
or \U$26102 ( \26445 , \26442 , \26217 );
nand \U$26103 ( \26446 , \26444 , \26445 );
not \U$26104 ( \26447 , \26446 );
not \U$26105 ( \26448 , \26365 );
not \U$26106 ( \26449 , \26373 );
and \U$26107 ( \26450 , \26448 , \26449 );
and \U$26108 ( \26451 , \26373 , \26365 );
nor \U$26109 ( \26452 , \26451 , \26380 );
nor \U$26110 ( \26453 , \26450 , \26452 );
not \U$26111 ( \26454 , \26392 );
not \U$26112 ( \26455 , \26400 );
and \U$26113 ( \26456 , \26454 , \26455 );
and \U$26114 ( \26457 , \26400 , \26392 );
nor \U$26115 ( \26458 , \26457 , \26407 );
nor \U$26116 ( \26459 , \26456 , \26458 );
xor \U$26117 ( \26460 , \26453 , \26459 );
and \U$26118 ( \26461 , \5318 , RI9870240_81);
and \U$26119 ( \26462 , RI98706f0_91, \5316 );
nor \U$26120 ( \26463 , \26461 , \26462 );
and \U$26121 ( \26464 , \26463 , \5322 );
not \U$26122 ( \26465 , \26463 );
and \U$26123 ( \26466 , \26465 , \5052 );
nor \U$26124 ( \26467 , \26464 , \26466 );
nand \U$26125 ( \26468 , RI9870420_85, \4201 );
and \U$26126 ( \26469 , \26468 , \3923 );
not \U$26127 ( \26470 , \26468 );
and \U$26128 ( \26471 , \26470 , \4207 );
nor \U$26129 ( \26472 , \26469 , \26471 );
xor \U$26130 ( \26473 , \26467 , \26472 );
and \U$26131 ( \26474 , \4710 , RI9870510_87);
and \U$26132 ( \26475 , RI9870330_83, \4708 );
nor \U$26133 ( \26476 , \26474 , \26475 );
not \U$26134 ( \26477 , \26476 );
not \U$26135 ( \26478 , \4519 );
and \U$26136 ( \26479 , \26477 , \26478 );
and \U$26137 ( \26480 , \26476 , \4521 );
nor \U$26138 ( \26481 , \26479 , \26480 );
xor \U$26139 ( \26482 , \26473 , \26481 );
xor \U$26140 ( \26483 , \26460 , \26482 );
not \U$26141 ( \26484 , \26483 );
and \U$26142 ( \26485 , \11696 , RI9870e70_107);
and \U$26143 ( \26486 , RI9870ba0_101, \11694 );
nor \U$26144 ( \26487 , \26485 , \26486 );
and \U$26145 ( \26488 , \26487 , \10965 );
not \U$26146 ( \26489 , \26487 );
and \U$26147 ( \26490 , \26489 , \11702 );
nor \U$26148 ( \26491 , \26488 , \26490 );
and \U$26149 ( \26492 , \12293 , RI9871050_111);
and \U$26150 ( \26493 , RI9870c90_103, \12291 );
nor \U$26151 ( \26494 , \26492 , \26493 );
and \U$26152 ( \26495 , \26494 , \11687 );
not \U$26153 ( \26496 , \26494 );
and \U$26154 ( \26497 , \26496 , \11686 );
nor \U$26155 ( \26498 , \26495 , \26497 );
xor \U$26156 ( \26499 , \26491 , \26498 );
and \U$26157 ( \26500 , \13045 , RI9871230_115);
and \U$26158 ( \26501 , RI9871140_113, \13043 );
nor \U$26159 ( \26502 , \26500 , \26501 );
and \U$26160 ( \26503 , \26502 , \13047 );
not \U$26161 ( \26504 , \26502 );
and \U$26162 ( \26505 , \26504 , \12619 );
nor \U$26163 ( \26506 , \26503 , \26505 );
and \U$26164 ( \26507 , \26499 , \26506 );
and \U$26165 ( \26508 , \26491 , \26498 );
or \U$26166 ( \26509 , \26507 , \26508 );
and \U$26167 ( \26510 , \13882 , RI9871320_117);
and \U$26168 ( \26511 , RI9871410_119, \13880 );
nor \U$26169 ( \26512 , \26510 , \26511 );
and \U$26170 ( \26513 , \26512 , \13358 );
not \U$26171 ( \26514 , \26512 );
and \U$26172 ( \26515 , \26514 , \13359 );
nor \U$26173 ( \26516 , \26513 , \26515 );
not \U$26174 ( \26517 , RI9873558_190);
and \U$26175 ( \26518 , \15780 , RI9871500_121);
and \U$26176 ( \26519 , RI9873648_192, RI98715f0_123);
nor \U$26177 ( \26520 , \26518 , \26519 );
not \U$26178 ( \26521 , \26520 );
or \U$26179 ( \26522 , \26517 , \26521 );
or \U$26180 ( \26523 , \26520 , RI9873558_190);
nand \U$26181 ( \26524 , \26522 , \26523 );
xor \U$26182 ( \26525 , \26516 , \26524 );
and \U$26183 ( \26526 , \14937 , RI98716e0_125);
and \U$26184 ( \26527 , RI98717d0_127, \14935 );
nor \U$26185 ( \26528 , \26526 , \26527 );
and \U$26186 ( \26529 , \26528 , \14539 );
not \U$26187 ( \26530 , \26528 );
and \U$26188 ( \26531 , \26530 , \14538 );
nor \U$26189 ( \26532 , \26529 , \26531 );
and \U$26190 ( \26533 , \26525 , \26532 );
and \U$26191 ( \26534 , \26516 , \26524 );
or \U$26192 ( \26535 , \26533 , \26534 );
xor \U$26193 ( \26536 , \26509 , \26535 );
xor \U$26194 ( \26537 , \26420 , \26427 );
and \U$26195 ( \26538 , \26537 , \26435 );
and \U$26196 ( \26539 , \26420 , \26427 );
or \U$26197 ( \26540 , \26538 , \26539 );
xor \U$26198 ( \26541 , \26536 , \26540 );
nand \U$26199 ( \26542 , \26484 , \26541 );
not \U$26200 ( \26543 , \26542 );
and \U$26201 ( \26544 , \26447 , \26543 );
and \U$26202 ( \26545 , \26446 , \26542 );
nor \U$26203 ( \26546 , \26544 , \26545 );
not \U$26204 ( \26547 , \26546 );
and \U$26205 ( \26548 , \8486 , RI986fd90_71);
and \U$26206 ( \26549 , RI986fca0_69, \8484 );
nor \U$26207 ( \26550 , \26548 , \26549 );
and \U$26208 ( \26551 , \26550 , \8050 );
not \U$26209 ( \26552 , \26550 );
and \U$26210 ( \26553 , \26552 , \8051 );
nor \U$26211 ( \26554 , \26551 , \26553 );
and \U$26212 ( \26555 , \7079 , RI98708d0_95);
and \U$26213 ( \26556 , RI98707e0_93, \7077 );
nor \U$26214 ( \26557 , \26555 , \26556 );
and \U$26215 ( \26558 , \26557 , \6710 );
not \U$26216 ( \26559 , \26557 );
and \U$26217 ( \26560 , \26559 , \6709 );
nor \U$26218 ( \26561 , \26558 , \26560 );
xor \U$26219 ( \26562 , \26554 , \26561 );
and \U$26220 ( \26563 , \7729 , RI986fac0_65);
and \U$26221 ( \26564 , RI986fbb0_67, \7727 );
nor \U$26222 ( \26565 , \26563 , \26564 );
and \U$26223 ( \26566 , \26565 , \7480 );
not \U$26224 ( \26567 , \26565 );
and \U$26225 ( \26568 , \26567 , \7733 );
nor \U$26226 ( \26569 , \26566 , \26568 );
and \U$26227 ( \26570 , \26562 , \26569 );
and \U$26228 ( \26571 , \26554 , \26561 );
or \U$26229 ( \26572 , \26570 , \26571 );
and \U$26230 ( \26573 , \5318 , RI9870510_87);
and \U$26231 ( \26574 , RI9870330_83, \5316 );
nor \U$26232 ( \26575 , \26573 , \26574 );
and \U$26233 ( \26576 , \26575 , \5052 );
not \U$26234 ( \26577 , \26575 );
and \U$26235 ( \26578 , \26577 , \5322 );
nor \U$26236 ( \26579 , \26576 , \26578 );
xor \U$26237 ( \26580 , \26572 , \26579 );
and \U$26238 ( \26581 , \5881 , RI9870330_83);
and \U$26239 ( \26582 , RI9870240_81, \5879 );
nor \U$26240 ( \26583 , \26581 , \26582 );
and \U$26241 ( \26584 , \26583 , \5594 );
not \U$26242 ( \26585 , \26583 );
and \U$26243 ( \26586 , \26585 , \5885 );
nor \U$26244 ( \26587 , \26584 , \26586 );
and \U$26245 ( \26588 , \5318 , RI9870420_85);
and \U$26246 ( \26589 , RI9870510_87, \5316 );
nor \U$26247 ( \26590 , \26588 , \26589 );
and \U$26248 ( \26591 , \26590 , \5052 );
not \U$26249 ( \26592 , \26590 );
and \U$26250 ( \26593 , \26592 , \5322 );
nor \U$26251 ( \26594 , \26591 , \26593 );
xor \U$26252 ( \26595 , \26587 , \26594 );
and \U$26253 ( \26596 , \6453 , RI98706f0_91);
and \U$26254 ( \26597 , RI9870600_89, \6451 );
nor \U$26255 ( \26598 , \26596 , \26597 );
and \U$26256 ( \26599 , \26598 , \6190 );
not \U$26257 ( \26600 , \26598 );
and \U$26258 ( \26601 , \26600 , \6180 );
nor \U$26259 ( \26602 , \26599 , \26601 );
and \U$26260 ( \26603 , \26595 , \26602 );
and \U$26261 ( \26604 , \26587 , \26594 );
or \U$26262 ( \26605 , \26603 , \26604 );
xor \U$26263 ( \26606 , \26580 , \26605 );
xor \U$26264 ( \26607 , \26337 , \26344 );
xor \U$26265 ( \26608 , \26607 , \26352 );
nand \U$26266 ( \26609 , RI9870420_85, \4708 );
not \U$26267 ( \26610 , \26609 );
not \U$26268 ( \26611 , \4521 );
or \U$26269 ( \26612 , \26610 , \26611 );
or \U$26270 ( \26613 , \4519 , \26609 );
nand \U$26271 ( \26614 , \26612 , \26613 );
xor \U$26272 ( \26615 , \26608 , \26614 );
xor \U$26273 ( \26616 , \26300 , \26307 );
xor \U$26274 ( \26617 , \26616 , \26315 );
xor \U$26275 ( \26618 , \26615 , \26617 );
and \U$26276 ( \26619 , \26606 , \26618 );
xor \U$26277 ( \26620 , \26225 , \26232 );
xor \U$26278 ( \26621 , \26620 , \26240 );
xor \U$26279 ( \26622 , \26273 , \26280 );
xor \U$26280 ( \26623 , \26622 , \26288 );
xor \U$26281 ( \26624 , \26251 , \4521 );
xor \U$26282 ( \26625 , \26624 , \26259 );
xor \U$26283 ( \26626 , \26623 , \26625 );
xor \U$26284 ( \26627 , \26621 , \26626 );
xor \U$26285 ( \26628 , \26608 , \26614 );
xor \U$26286 ( \26629 , \26628 , \26617 );
and \U$26287 ( \26630 , \26627 , \26629 );
and \U$26288 ( \26631 , \26606 , \26627 );
or \U$26289 ( \26632 , \26619 , \26630 , \26631 );
and \U$26290 ( \26633 , \8486 , RI986fbb0_67);
and \U$26291 ( \26634 , RI986fd90_71, \8484 );
nor \U$26292 ( \26635 , \26633 , \26634 );
and \U$26293 ( \26636 , \26635 , \8050 );
not \U$26294 ( \26637 , \26635 );
and \U$26295 ( \26638 , \26637 , \8051 );
nor \U$26296 ( \26639 , \26636 , \26638 );
and \U$26297 ( \26640 , \7729 , RI98707e0_93);
and \U$26298 ( \26641 , RI986fac0_65, \7727 );
nor \U$26299 ( \26642 , \26640 , \26641 );
and \U$26300 ( \26643 , \26642 , \7480 );
not \U$26301 ( \26644 , \26642 );
and \U$26302 ( \26645 , \26644 , \7733 );
nor \U$26303 ( \26646 , \26643 , \26645 );
xor \U$26304 ( \26647 , \26639 , \26646 );
and \U$26305 ( \26648 , \9237 , RI986fca0_69);
and \U$26306 ( \26649 , RI986ff70_75, \9235 );
nor \U$26307 ( \26650 , \26648 , \26649 );
and \U$26308 ( \26651 , \26650 , \9241 );
not \U$26309 ( \26652 , \26650 );
and \U$26310 ( \26653 , \26652 , \8836 );
nor \U$26311 ( \26654 , \26651 , \26653 );
and \U$26312 ( \26655 , \26647 , \26654 );
and \U$26313 ( \26656 , \26639 , \26646 );
or \U$26314 ( \26657 , \26655 , \26656 );
and \U$26315 ( \26658 , \5881 , RI9870510_87);
and \U$26316 ( \26659 , RI9870330_83, \5879 );
nor \U$26317 ( \26660 , \26658 , \26659 );
and \U$26318 ( \26661 , \26660 , \5594 );
not \U$26319 ( \26662 , \26660 );
and \U$26320 ( \26663 , \26662 , \5885 );
nor \U$26321 ( \26664 , \26661 , \26663 );
and \U$26322 ( \26665 , \6453 , RI9870240_81);
and \U$26323 ( \26666 , RI98706f0_91, \6451 );
nor \U$26324 ( \26667 , \26665 , \26666 );
and \U$26325 ( \26668 , \26667 , \6190 );
not \U$26326 ( \26669 , \26667 );
and \U$26327 ( \26670 , \26669 , \6180 );
nor \U$26328 ( \26671 , \26668 , \26670 );
xor \U$26329 ( \26672 , \26664 , \26671 );
and \U$26330 ( \26673 , \7079 , RI9870600_89);
and \U$26331 ( \26674 , RI98708d0_95, \7077 );
nor \U$26332 ( \26675 , \26673 , \26674 );
and \U$26333 ( \26676 , \26675 , \6710 );
not \U$26334 ( \26677 , \26675 );
and \U$26335 ( \26678 , \26677 , \6709 );
nor \U$26336 ( \26679 , \26676 , \26678 );
and \U$26337 ( \26680 , \26672 , \26679 );
and \U$26338 ( \26681 , \26664 , \26671 );
or \U$26339 ( \26682 , \26680 , \26681 );
xor \U$26340 ( \26683 , \26657 , \26682 );
xor \U$26341 ( \26684 , \26587 , \26594 );
xor \U$26342 ( \26685 , \26684 , \26602 );
and \U$26343 ( \26686 , \26683 , \26685 );
and \U$26344 ( \26687 , \26657 , \26682 );
or \U$26345 ( \26688 , \26686 , \26687 );
and \U$26346 ( \26689 , \11696 , RI9870ab0_99);
and \U$26347 ( \26690 , RI9870d80_105, \11694 );
nor \U$26348 ( \26691 , \26689 , \26690 );
and \U$26349 ( \26692 , \26691 , \10965 );
not \U$26350 ( \26693 , \26691 );
and \U$26351 ( \26694 , \26693 , \11702 );
nor \U$26352 ( \26695 , \26692 , \26694 );
and \U$26353 ( \26696 , \9505 , RI986fe80_73);
and \U$26354 ( \26697 , RI9870060_77, \9503 );
nor \U$26355 ( \26698 , \26696 , \26697 );
and \U$26356 ( \26699 , \26698 , \9510 );
not \U$26357 ( \26700 , \26698 );
and \U$26358 ( \26701 , \26700 , \9513 );
nor \U$26359 ( \26702 , \26699 , \26701 );
xor \U$26360 ( \26703 , \26695 , \26702 );
and \U$26361 ( \26704 , \10424 , RI9870150_79);
and \U$26362 ( \26705 , RI9870f60_109, \10422 );
nor \U$26363 ( \26706 , \26704 , \26705 );
and \U$26364 ( \26707 , \26706 , \9840 );
not \U$26365 ( \26708 , \26706 );
and \U$26366 ( \26709 , \26708 , \10428 );
nor \U$26367 ( \26710 , \26707 , \26709 );
and \U$26368 ( \26711 , \26703 , \26710 );
and \U$26369 ( \26712 , \26695 , \26702 );
or \U$26370 ( \26713 , \26711 , \26712 );
not \U$26371 ( \26714 , RI9873558_190);
and \U$26372 ( \26715 , \15780 , RI9871410_119);
and \U$26373 ( \26716 , RI9873648_192, RI98716e0_125);
nor \U$26374 ( \26717 , \26715 , \26716 );
not \U$26375 ( \26718 , \26717 );
or \U$26376 ( \26719 , \26714 , \26718 );
or \U$26377 ( \26720 , \26717 , RI9873558_190);
nand \U$26378 ( \26721 , \26719 , \26720 );
xor \U$26379 ( \26722 , \26721 , \5322 );
and \U$26380 ( \26723 , \14937 , RI9871140_113);
and \U$26381 ( \26724 , RI9871320_117, \14935 );
nor \U$26382 ( \26725 , \26723 , \26724 );
and \U$26383 ( \26726 , \26725 , \14539 );
not \U$26384 ( \26727 , \26725 );
and \U$26385 ( \26728 , \26727 , \14538 );
nor \U$26386 ( \26729 , \26726 , \26728 );
and \U$26387 ( \26730 , \26722 , \26729 );
and \U$26388 ( \26731 , \26721 , \5322 );
or \U$26389 ( \26732 , \26730 , \26731 );
xor \U$26390 ( \26733 , \26713 , \26732 );
and \U$26391 ( \26734 , \13882 , RI9870c90_103);
and \U$26392 ( \26735 , RI9871230_115, \13880 );
nor \U$26393 ( \26736 , \26734 , \26735 );
and \U$26394 ( \26737 , \26736 , \13358 );
not \U$26395 ( \26738 , \26736 );
and \U$26396 ( \26739 , \26738 , \13359 );
nor \U$26397 ( \26740 , \26737 , \26739 );
and \U$26398 ( \26741 , \12293 , RI98709c0_97);
and \U$26399 ( \26742 , RI9870e70_107, \12291 );
nor \U$26400 ( \26743 , \26741 , \26742 );
and \U$26401 ( \26744 , \26743 , \11687 );
not \U$26402 ( \26745 , \26743 );
and \U$26403 ( \26746 , \26745 , \11686 );
nor \U$26404 ( \26747 , \26744 , \26746 );
xor \U$26405 ( \26748 , \26740 , \26747 );
and \U$26406 ( \26749 , \13045 , RI9870ba0_101);
and \U$26407 ( \26750 , RI9871050_111, \13043 );
nor \U$26408 ( \26751 , \26749 , \26750 );
and \U$26409 ( \26752 , \26751 , \13047 );
not \U$26410 ( \26753 , \26751 );
and \U$26411 ( \26754 , \26753 , \12619 );
nor \U$26412 ( \26755 , \26752 , \26754 );
and \U$26413 ( \26756 , \26748 , \26755 );
and \U$26414 ( \26757 , \26740 , \26747 );
or \U$26415 ( \26758 , \26756 , \26757 );
and \U$26416 ( \26759 , \26733 , \26758 );
and \U$26417 ( \26760 , \26713 , \26732 );
or \U$26418 ( \26761 , \26759 , \26760 );
xor \U$26419 ( \26762 , \26688 , \26761 );
and \U$26420 ( \26763 , \11696 , RI9870d80_105);
and \U$26421 ( \26764 , RI98709c0_97, \11694 );
nor \U$26422 ( \26765 , \26763 , \26764 );
and \U$26423 ( \26766 , \26765 , \11702 );
not \U$26424 ( \26767 , \26765 );
and \U$26425 ( \26768 , \26767 , \10965 );
nor \U$26426 ( \26769 , \26766 , \26768 );
not \U$26427 ( \26770 , \26769 );
and \U$26428 ( \26771 , \12293 , RI9870e70_107);
and \U$26429 ( \26772 , RI9870ba0_101, \12291 );
nor \U$26430 ( \26773 , \26771 , \26772 );
and \U$26431 ( \26774 , \26773 , \11686 );
not \U$26432 ( \26775 , \26773 );
and \U$26433 ( \26776 , \26775 , \11687 );
nor \U$26434 ( \26777 , \26774 , \26776 );
and \U$26435 ( \26778 , \13045 , RI9871050_111);
and \U$26436 ( \26779 , RI9870c90_103, \13043 );
nor \U$26437 ( \26780 , \26778 , \26779 );
and \U$26438 ( \26781 , \26780 , \12619 );
not \U$26439 ( \26782 , \26780 );
and \U$26440 ( \26783 , \26782 , \13047 );
nor \U$26441 ( \26784 , \26781 , \26783 );
xor \U$26442 ( \26785 , \26777 , \26784 );
not \U$26443 ( \26786 , \26785 );
or \U$26444 ( \26787 , \26770 , \26786 );
or \U$26445 ( \26788 , \26785 , \26769 );
nand \U$26446 ( \26789 , \26787 , \26788 );
xor \U$26447 ( \26790 , \26554 , \26561 );
xor \U$26448 ( \26791 , \26790 , \26569 );
xor \U$26449 ( \26792 , \26789 , \26791 );
and \U$26450 ( \26793 , \9237 , RI986ff70_75);
and \U$26451 ( \26794 , RI986fe80_73, \9235 );
nor \U$26452 ( \26795 , \26793 , \26794 );
and \U$26453 ( \26796 , \26795 , \8836 );
not \U$26454 ( \26797 , \26795 );
and \U$26455 ( \26798 , \26797 , \9241 );
nor \U$26456 ( \26799 , \26796 , \26798 );
not \U$26457 ( \26800 , \26799 );
and \U$26458 ( \26801 , \9505 , RI9870060_77);
and \U$26459 ( \26802 , RI9870150_79, \9503 );
nor \U$26460 ( \26803 , \26801 , \26802 );
and \U$26461 ( \26804 , \26803 , \9513 );
not \U$26462 ( \26805 , \26803 );
and \U$26463 ( \26806 , \26805 , \9510 );
nor \U$26464 ( \26807 , \26804 , \26806 );
and \U$26465 ( \26808 , \10424 , RI9870f60_109);
and \U$26466 ( \26809 , RI9870ab0_99, \10422 );
nor \U$26467 ( \26810 , \26808 , \26809 );
and \U$26468 ( \26811 , \26810 , \10428 );
not \U$26469 ( \26812 , \26810 );
and \U$26470 ( \26813 , \26812 , \9840 );
nor \U$26471 ( \26814 , \26811 , \26813 );
xor \U$26472 ( \26815 , \26807 , \26814 );
not \U$26473 ( \26816 , \26815 );
or \U$26474 ( \26817 , \26800 , \26816 );
or \U$26475 ( \26818 , \26815 , \26799 );
nand \U$26476 ( \26819 , \26817 , \26818 );
and \U$26477 ( \26820 , \26792 , \26819 );
and \U$26478 ( \26821 , \26789 , \26791 );
or \U$26479 ( \26822 , \26820 , \26821 );
and \U$26480 ( \26823 , \26762 , \26822 );
and \U$26481 ( \26824 , \26688 , \26761 );
or \U$26482 ( \26825 , \26823 , \26824 );
xor \U$26483 ( \26826 , \26632 , \26825 );
not \U$26484 ( \26827 , \26262 );
not \U$26485 ( \26828 , \26291 );
not \U$26486 ( \26829 , \26243 );
and \U$26487 ( \26830 , \26828 , \26829 );
and \U$26488 ( \26831 , \26291 , \26243 );
nor \U$26489 ( \26832 , \26830 , \26831 );
not \U$26490 ( \26833 , \26832 );
or \U$26491 ( \26834 , \26827 , \26833 );
or \U$26492 ( \26835 , \26832 , \26262 );
nand \U$26493 ( \26836 , \26834 , \26835 );
not \U$26494 ( \26837 , \26327 );
xor \U$26495 ( \26838 , \26318 , \26355 );
not \U$26496 ( \26839 , \26838 );
or \U$26497 ( \26840 , \26837 , \26839 );
or \U$26498 ( \26841 , \26838 , \26327 );
nand \U$26499 ( \26842 , \26840 , \26841 );
xor \U$26500 ( \26843 , \26836 , \26842 );
xor \U$26501 ( \26844 , \26385 , \26412 );
xor \U$26502 ( \26845 , \26844 , \26436 );
xor \U$26503 ( \26846 , \26843 , \26845 );
and \U$26504 ( \26847 , \26826 , \26846 );
and \U$26505 ( \26848 , \26632 , \26825 );
or \U$26506 ( \26849 , \26847 , \26848 );
not \U$26507 ( \26850 , \26799 );
not \U$26508 ( \26851 , \26807 );
and \U$26509 ( \26852 , \26850 , \26851 );
and \U$26510 ( \26853 , \26807 , \26799 );
nor \U$26511 ( \26854 , \26853 , \26814 );
nor \U$26512 ( \26855 , \26852 , \26854 );
not \U$26513 ( \26856 , \26769 );
not \U$26514 ( \26857 , \26784 );
and \U$26515 ( \26858 , \26856 , \26857 );
and \U$26516 ( \26859 , \26784 , \26769 );
nor \U$26517 ( \26860 , \26859 , \26777 );
nor \U$26518 ( \26861 , \26858 , \26860 );
xor \U$26519 ( \26862 , \26855 , \26861 );
and \U$26520 ( \26863 , \14937 , RI9871320_117);
and \U$26521 ( \26864 , RI9871410_119, \14935 );
nor \U$26522 ( \26865 , \26863 , \26864 );
and \U$26523 ( \26866 , \26865 , \14539 );
not \U$26524 ( \26867 , \26865 );
and \U$26525 ( \26868 , \26867 , \14538 );
nor \U$26526 ( \26869 , \26866 , \26868 );
not \U$26527 ( \26870 , RI9873558_190);
and \U$26528 ( \26871 , \15780 , RI98716e0_125);
and \U$26529 ( \26872 , RI9873648_192, RI98717d0_127);
nor \U$26530 ( \26873 , \26871 , \26872 );
not \U$26531 ( \26874 , \26873 );
or \U$26532 ( \26875 , \26870 , \26874 );
or \U$26533 ( \26876 , \26873 , RI9873558_190);
nand \U$26534 ( \26877 , \26875 , \26876 );
xor \U$26535 ( \26878 , \26869 , \26877 );
and \U$26536 ( \26879 , \13882 , RI9871230_115);
and \U$26537 ( \26880 , RI9871140_113, \13880 );
nor \U$26538 ( \26881 , \26879 , \26880 );
and \U$26539 ( \26882 , \26881 , \13358 );
not \U$26540 ( \26883 , \26881 );
and \U$26541 ( \26884 , \26883 , \13359 );
nor \U$26542 ( \26885 , \26882 , \26884 );
and \U$26543 ( \26886 , \26878 , \26885 );
and \U$26544 ( \26887 , \26869 , \26877 );
nor \U$26545 ( \26888 , \26886 , \26887 );
and \U$26546 ( \26889 , \26862 , \26888 );
and \U$26547 ( \26890 , \26855 , \26861 );
nor \U$26548 ( \26891 , \26889 , \26890 );
xor \U$26549 ( \26892 , \26572 , \26579 );
and \U$26550 ( \26893 , \26892 , \26605 );
and \U$26551 ( \26894 , \26572 , \26579 );
or \U$26552 ( \26895 , \26893 , \26894 );
xor \U$26553 ( \26896 , \26891 , \26895 );
xor \U$26554 ( \26897 , \26608 , \26614 );
and \U$26555 ( \26898 , \26897 , \26617 );
and \U$26556 ( \26899 , \26608 , \26614 );
or \U$26557 ( \26900 , \26898 , \26899 );
xor \U$26558 ( \26901 , \26896 , \26900 );
xor \U$26559 ( \26902 , \26491 , \26498 );
xor \U$26560 ( \26903 , \26902 , \26506 );
xor \U$26561 ( \26904 , \26516 , \26524 );
xor \U$26562 ( \26905 , \26904 , \26532 );
xor \U$26563 ( \26906 , \26225 , \26232 );
xor \U$26564 ( \26907 , \26906 , \26240 );
and \U$26565 ( \26908 , \26623 , \26907 );
xor \U$26566 ( \26909 , \26225 , \26232 );
xor \U$26567 ( \26910 , \26909 , \26240 );
and \U$26568 ( \26911 , \26625 , \26910 );
and \U$26569 ( \26912 , \26623 , \26625 );
or \U$26570 ( \26913 , \26908 , \26911 , \26912 );
xor \U$26571 ( \26914 , \26905 , \26913 );
xor \U$26572 ( \26915 , \26903 , \26914 );
and \U$26573 ( \26916 , \26901 , \26915 );
xor \U$26574 ( \26917 , \26849 , \26916 );
not \U$26575 ( \26918 , \26541 );
not \U$26576 ( \26919 , \26483 );
and \U$26577 ( \26920 , \26918 , \26919 );
and \U$26578 ( \26921 , \26541 , \26483 );
nor \U$26579 ( \26922 , \26920 , \26921 );
not \U$26580 ( \26923 , \26922 );
not \U$26581 ( \26924 , \26214 );
xor \U$26582 ( \26925 , \26141 , \26118 );
not \U$26583 ( \26926 , \26925 );
and \U$26584 ( \26927 , \26924 , \26926 );
and \U$26585 ( \26928 , \26214 , \26925 );
nor \U$26586 ( \26929 , \26927 , \26928 );
xor \U$26587 ( \26930 , \26293 , \26357 );
xor \U$26588 ( \26931 , \26930 , \26439 );
xor \U$26589 ( \26932 , \26929 , \26931 );
not \U$26590 ( \26933 , \26932 );
or \U$26591 ( \26934 , \26923 , \26933 );
or \U$26592 ( \26935 , \26932 , \26922 );
nand \U$26593 ( \26936 , \26934 , \26935 );
and \U$26594 ( \26937 , \26917 , \26936 );
and \U$26595 ( \26938 , \26849 , \26916 );
or \U$26596 ( \26939 , \26937 , \26938 );
not \U$26597 ( \26940 , \26939 );
or \U$26598 ( \26941 , \26547 , \26940 );
or \U$26599 ( \26942 , \26939 , \26546 );
nand \U$26600 ( \26943 , \26941 , \26942 );
not \U$26601 ( \26944 , \26943 );
xor \U$26602 ( \26945 , \26891 , \26895 );
and \U$26603 ( \26946 , \26945 , \26900 );
and \U$26604 ( \26947 , \26891 , \26895 );
or \U$26605 ( \26948 , \26946 , \26947 );
xor \U$26606 ( \26949 , \26491 , \26498 );
xor \U$26607 ( \26950 , \26949 , \26506 );
and \U$26608 ( \26951 , \26905 , \26950 );
xor \U$26609 ( \26952 , \26491 , \26498 );
xor \U$26610 ( \26953 , \26952 , \26506 );
and \U$26611 ( \26954 , \26913 , \26953 );
and \U$26612 ( \26955 , \26905 , \26913 );
or \U$26613 ( \26956 , \26951 , \26954 , \26955 );
xor \U$26614 ( \26957 , \26948 , \26956 );
xor \U$26615 ( \26958 , \26836 , \26842 );
and \U$26616 ( \26959 , \26958 , \26845 );
and \U$26617 ( \26960 , \26836 , \26842 );
or \U$26618 ( \26961 , \26959 , \26960 );
and \U$26619 ( \26962 , \26957 , \26961 );
and \U$26620 ( \26963 , \26948 , \26956 );
or \U$26621 ( \26964 , \26962 , \26963 );
not \U$26622 ( \26965 , \26964 );
not \U$26623 ( \26966 , \26931 );
not \U$26624 ( \26967 , \26922 );
and \U$26625 ( \26968 , \26966 , \26967 );
and \U$26626 ( \26969 , \26931 , \26922 );
nor \U$26627 ( \26970 , \26969 , \26929 );
nor \U$26628 ( \26971 , \26968 , \26970 );
not \U$26629 ( \26972 , \26971 );
or \U$26630 ( \26973 , \26965 , \26972 );
or \U$26631 ( \26974 , \26971 , \26964 );
nand \U$26632 ( \26975 , \26973 , \26974 );
not \U$26633 ( \26976 , \26975 );
xor \U$26634 ( \26977 , \26109 , \4207 );
and \U$26635 ( \26978 , \26977 , \26117 );
and \U$26636 ( \26979 , \26109 , \4207 );
or \U$26637 ( \26980 , \26978 , \26979 );
xor \U$26638 ( \26981 , \26196 , \26203 );
and \U$26639 ( \26982 , \26981 , \26211 );
and \U$26640 ( \26983 , \26196 , \26203 );
or \U$26641 ( \26984 , \26982 , \26983 );
xor \U$26642 ( \26985 , \26980 , \26984 );
xor \U$26643 ( \26986 , \26125 , \26132 );
and \U$26644 ( \26987 , \26986 , \26140 );
and \U$26645 ( \26988 , \26125 , \26132 );
or \U$26646 ( \26989 , \26987 , \26988 );
xor \U$26647 ( \26990 , \26985 , \26989 );
xor \U$26648 ( \26991 , \26509 , \26535 );
and \U$26649 ( \26992 , \26991 , \26540 );
and \U$26650 ( \26993 , \26509 , \26535 );
nor \U$26651 ( \26994 , \26992 , \26993 );
xor \U$26652 ( \26995 , \26150 , \26157 );
xor \U$26653 ( \26996 , \26995 , \26165 );
and \U$26654 ( \26997 , \26189 , \26996 );
xor \U$26655 ( \26998 , \26150 , \26157 );
xor \U$26656 ( \26999 , \26998 , \26165 );
and \U$26657 ( \27000 , \26212 , \26999 );
and \U$26658 ( \27001 , \26189 , \26212 );
or \U$26659 ( \27002 , \26997 , \27000 , \27001 );
xor \U$26660 ( \27003 , \26994 , \27002 );
xor \U$26661 ( \27004 , \26453 , \26459 );
and \U$26662 ( \27005 , \27004 , \26482 );
and \U$26663 ( \27006 , \26453 , \26459 );
or \U$26664 ( \27007 , \27005 , \27006 );
xor \U$26665 ( \27008 , \27003 , \27007 );
xor \U$26666 ( \27009 , \26990 , \27008 );
and \U$26667 ( \27010 , \7729 , RI986ff70_75);
and \U$26668 ( \27011 , RI986fe80_73, \7727 );
nor \U$26669 ( \27012 , \27010 , \27011 );
and \U$26670 ( \27013 , \27012 , \7480 );
not \U$26671 ( \27014 , \27012 );
and \U$26672 ( \27015 , \27014 , \7733 );
nor \U$26673 ( \27016 , \27013 , \27015 );
and \U$26674 ( \27017 , \8486 , RI9870060_77);
and \U$26675 ( \27018 , RI9870150_79, \8484 );
nor \U$26676 ( \27019 , \27017 , \27018 );
and \U$26677 ( \27020 , \27019 , \8050 );
not \U$26678 ( \27021 , \27019 );
and \U$26679 ( \27022 , \27021 , \8051 );
nor \U$26680 ( \27023 , \27020 , \27022 );
xor \U$26681 ( \27024 , \27016 , \27023 );
and \U$26682 ( \27025 , \7079 , RI986fd90_71);
and \U$26683 ( \27026 , RI986fca0_69, \7077 );
nor \U$26684 ( \27027 , \27025 , \27026 );
and \U$26685 ( \27028 , \27027 , \6710 );
not \U$26686 ( \27029 , \27027 );
and \U$26687 ( \27030 , \27029 , \6709 );
nor \U$26688 ( \27031 , \27028 , \27030 );
xor \U$26689 ( \27032 , \27024 , \27031 );
and \U$26690 ( \27033 , \6453 , RI986fac0_65);
and \U$26691 ( \27034 , RI986fbb0_67, \6451 );
nor \U$26692 ( \27035 , \27033 , \27034 );
and \U$26693 ( \27036 , \27035 , \6190 );
not \U$26694 ( \27037 , \27035 );
and \U$26695 ( \27038 , \27037 , \6180 );
nor \U$26696 ( \27039 , \27036 , \27038 );
and \U$26697 ( \27040 , \5318 , RI98706f0_91);
and \U$26698 ( \27041 , RI9870600_89, \5316 );
nor \U$26699 ( \27042 , \27040 , \27041 );
and \U$26700 ( \27043 , \27042 , \5052 );
not \U$26701 ( \27044 , \27042 );
and \U$26702 ( \27045 , \27044 , \5322 );
nor \U$26703 ( \27046 , \27043 , \27045 );
xor \U$26704 ( \27047 , \27039 , \27046 );
and \U$26705 ( \27048 , \5881 , RI98708d0_95);
and \U$26706 ( \27049 , RI98707e0_93, \5879 );
nor \U$26707 ( \27050 , \27048 , \27049 );
and \U$26708 ( \27051 , \27050 , \5594 );
not \U$26709 ( \27052 , \27050 );
and \U$26710 ( \27053 , \27052 , \5885 );
nor \U$26711 ( \27054 , \27051 , \27053 );
xor \U$26712 ( \27055 , \27047 , \27054 );
xnor \U$26713 ( \27056 , \27032 , \27055 );
not \U$26714 ( \27057 , \27056 );
and \U$26715 ( \27058 , \4203 , RI9870420_85);
and \U$26716 ( \27059 , RI9870510_87, \4201 );
nor \U$26717 ( \27060 , \27058 , \27059 );
and \U$26718 ( \27061 , \27060 , \3922 );
not \U$26719 ( \27062 , \27060 );
and \U$26720 ( \27063 , \27062 , \4207 );
nor \U$26721 ( \27064 , \27061 , \27063 );
not \U$26722 ( \27065 , \27064 );
not \U$26723 ( \27066 , \4521 );
and \U$26724 ( \27067 , \4710 , RI9870330_83);
and \U$26725 ( \27068 , RI9870240_81, \4708 );
nor \U$26726 ( \27069 , \27067 , \27068 );
not \U$26727 ( \27070 , \27069 );
or \U$26728 ( \27071 , \27066 , \27070 );
or \U$26729 ( \27072 , \27069 , \4521 );
nand \U$26730 ( \27073 , \27071 , \27072 );
not \U$26731 ( \27074 , \27073 );
or \U$26732 ( \27075 , \27065 , \27074 );
or \U$26733 ( \27076 , \27064 , \27073 );
nand \U$26734 ( \27077 , \27075 , \27076 );
not \U$26735 ( \27078 , \27077 );
and \U$26736 ( \27079 , \27057 , \27078 );
and \U$26737 ( \27080 , \27056 , \27077 );
nor \U$26738 ( \27081 , \27079 , \27080 );
xor \U$26739 ( \27082 , \26467 , \26472 );
and \U$26740 ( \27083 , \27082 , \26481 );
and \U$26741 ( \27084 , \26467 , \26472 );
or \U$26742 ( \27085 , \27083 , \27084 );
xor \U$26743 ( \27086 , \26173 , \26180 );
and \U$26744 ( \27087 , \27086 , \26188 );
and \U$26745 ( \27088 , \26173 , \26180 );
or \U$26746 ( \27089 , \27087 , \27088 );
xor \U$26747 ( \27090 , \27085 , \27089 );
xor \U$26748 ( \27091 , \26150 , \26157 );
and \U$26749 ( \27092 , \27091 , \26165 );
and \U$26750 ( \27093 , \26150 , \26157 );
or \U$26751 ( \27094 , \27092 , \27093 );
xor \U$26752 ( \27095 , \27090 , \27094 );
xor \U$26753 ( \27096 , \27081 , \27095 );
and \U$26754 ( \27097 , \9505 , RI9870d80_105);
and \U$26755 ( \27098 , RI98709c0_97, \9503 );
nor \U$26756 ( \27099 , \27097 , \27098 );
and \U$26757 ( \27100 , \27099 , \9513 );
not \U$26758 ( \27101 , \27099 );
and \U$26759 ( \27102 , \27101 , \9510 );
nor \U$26760 ( \27103 , \27100 , \27102 );
and \U$26761 ( \27104 , \9237 , RI9870f60_109);
and \U$26762 ( \27105 , RI9870ab0_99, \9235 );
nor \U$26763 ( \27106 , \27104 , \27105 );
and \U$26764 ( \27107 , \27106 , \8836 );
not \U$26765 ( \27108 , \27106 );
and \U$26766 ( \27109 , \27108 , \9241 );
nor \U$26767 ( \27110 , \27107 , \27109 );
xor \U$26768 ( \27111 , \27103 , \27110 );
and \U$26769 ( \27112 , \10424 , RI9870e70_107);
and \U$26770 ( \27113 , RI9870ba0_101, \10422 );
nor \U$26771 ( \27114 , \27112 , \27113 );
and \U$26772 ( \27115 , \27114 , \10428 );
not \U$26773 ( \27116 , \27114 );
and \U$26774 ( \27117 , \27116 , \9840 );
nor \U$26775 ( \27118 , \27115 , \27117 );
xor \U$26776 ( \27119 , \27111 , \27118 );
and \U$26777 ( \27120 , \13882 , RI98716e0_125);
and \U$26778 ( \27121 , RI98717d0_127, \13880 );
nor \U$26779 ( \27122 , \27120 , \27121 );
and \U$26780 ( \27123 , \27122 , \13359 );
not \U$26781 ( \27124 , \27122 );
and \U$26782 ( \27125 , \27124 , \13358 );
nor \U$26783 ( \27126 , \27123 , \27125 );
and \U$26784 ( \27127 , \15780 , RI986ead0_31);
and \U$26785 ( \27128 , RI9873648_192, RI986e9e0_29);
nor \U$26786 ( \27129 , \27127 , \27128 );
not \U$26787 ( \27130 , \27129 );
not \U$26788 ( \27131 , RI9873558_190);
and \U$26789 ( \27132 , \27130 , \27131 );
and \U$26790 ( \27133 , \27129 , RI9873558_190);
nor \U$26791 ( \27134 , \27132 , \27133 );
xor \U$26792 ( \27135 , \27126 , \27134 );
and \U$26793 ( \27136 , \14937 , RI9871500_121);
and \U$26794 ( \27137 , RI98715f0_123, \14935 );
nor \U$26795 ( \27138 , \27136 , \27137 );
and \U$26796 ( \27139 , \27138 , \14538 );
not \U$26797 ( \27140 , \27138 );
and \U$26798 ( \27141 , \27140 , \14539 );
nor \U$26799 ( \27142 , \27139 , \27141 );
xor \U$26800 ( \27143 , \27135 , \27142 );
xor \U$26801 ( \27144 , \27119 , \27143 );
and \U$26802 ( \27145 , \13045 , RI9871320_117);
and \U$26803 ( \27146 , RI9871410_119, \13043 );
nor \U$26804 ( \27147 , \27145 , \27146 );
and \U$26805 ( \27148 , \27147 , \12619 );
not \U$26806 ( \27149 , \27147 );
and \U$26807 ( \27150 , \27149 , \13047 );
nor \U$26808 ( \27151 , \27148 , \27150 );
and \U$26809 ( \27152 , \11696 , RI9871050_111);
and \U$26810 ( \27153 , RI9870c90_103, \11694 );
nor \U$26811 ( \27154 , \27152 , \27153 );
and \U$26812 ( \27155 , \27154 , \11702 );
not \U$26813 ( \27156 , \27154 );
and \U$26814 ( \27157 , \27156 , \10965 );
nor \U$26815 ( \27158 , \27155 , \27157 );
xor \U$26816 ( \27159 , \27151 , \27158 );
and \U$26817 ( \27160 , \12293 , RI9871230_115);
and \U$26818 ( \27161 , RI9871140_113, \12291 );
nor \U$26819 ( \27162 , \27160 , \27161 );
and \U$26820 ( \27163 , \27162 , \11686 );
not \U$26821 ( \27164 , \27162 );
and \U$26822 ( \27165 , \27164 , \11687 );
nor \U$26823 ( \27166 , \27163 , \27165 );
xor \U$26824 ( \27167 , \27159 , \27166 );
xor \U$26825 ( \27168 , \27144 , \27167 );
xor \U$26826 ( \27169 , \27096 , \27168 );
xor \U$26827 ( \27170 , \27009 , \27169 );
not \U$26828 ( \27171 , \27170 );
and \U$26829 ( \27172 , \26976 , \27171 );
and \U$26830 ( \27173 , \26975 , \27170 );
nor \U$26831 ( \27174 , \27172 , \27173 );
not \U$26832 ( \27175 , \27174 );
and \U$26833 ( \27176 , \26944 , \27175 );
and \U$26834 ( \27177 , \26943 , \27174 );
nor \U$26835 ( \27178 , \27176 , \27177 );
xor \U$26836 ( \27179 , \26849 , \26916 );
xor \U$26837 ( \27180 , \27179 , \26936 );
xor \U$26838 ( \27181 , \26948 , \26956 );
xor \U$26839 ( \27182 , \27181 , \26961 );
xor \U$26840 ( \27183 , \27180 , \27182 );
xor \U$26841 ( \27184 , \26901 , \26915 );
not \U$26842 ( \27185 , \27184 );
xor \U$26843 ( \27186 , \26632 , \26825 );
xor \U$26844 ( \27187 , \27186 , \26846 );
not \U$26845 ( \27188 , \27187 );
or \U$26846 ( \27189 , \27185 , \27188 );
or \U$26847 ( \27190 , \27187 , \27184 );
xor \U$26848 ( \27191 , \26740 , \26747 );
xor \U$26849 ( \27192 , \27191 , \26755 );
xor \U$26850 ( \27193 , \26695 , \26702 );
xor \U$26851 ( \27194 , \27193 , \26710 );
and \U$26852 ( \27195 , \27192 , \27194 );
xor \U$26853 ( \27196 , \26639 , \26646 );
xor \U$26854 ( \27197 , \27196 , \26654 );
xor \U$26855 ( \27198 , \26695 , \26702 );
xor \U$26856 ( \27199 , \27198 , \26710 );
and \U$26857 ( \27200 , \27197 , \27199 );
and \U$26858 ( \27201 , \27192 , \27197 );
or \U$26859 ( \27202 , \27195 , \27200 , \27201 );
not \U$26860 ( \27203 , \27202 );
not \U$26861 ( \27204 , \27203 );
xor \U$26862 ( \27205 , \26664 , \26671 );
xor \U$26863 ( \27206 , \27205 , \26679 );
nand \U$26864 ( \27207 , RI9870420_85, \5316 );
and \U$26865 ( \27208 , \27207 , \5052 );
not \U$26866 ( \27209 , \27207 );
and \U$26867 ( \27210 , \27209 , \5322 );
nor \U$26868 ( \27211 , \27208 , \27210 );
xor \U$26869 ( \27212 , \27206 , \27211 );
and \U$26870 ( \27213 , \7729 , RI98708d0_95);
and \U$26871 ( \27214 , RI98707e0_93, \7727 );
nor \U$26872 ( \27215 , \27213 , \27214 );
and \U$26873 ( \27216 , \27215 , \7480 );
not \U$26874 ( \27217 , \27215 );
and \U$26875 ( \27218 , \27217 , \7733 );
nor \U$26876 ( \27219 , \27216 , \27218 );
and \U$26877 ( \27220 , \7079 , RI98706f0_91);
and \U$26878 ( \27221 , RI9870600_89, \7077 );
nor \U$26879 ( \27222 , \27220 , \27221 );
and \U$26880 ( \27223 , \27222 , \6710 );
not \U$26881 ( \27224 , \27222 );
and \U$26882 ( \27225 , \27224 , \6709 );
nor \U$26883 ( \27226 , \27223 , \27225 );
xor \U$26884 ( \27227 , \27219 , \27226 );
and \U$26885 ( \27228 , \8486 , RI986fac0_65);
and \U$26886 ( \27229 , RI986fbb0_67, \8484 );
nor \U$26887 ( \27230 , \27228 , \27229 );
and \U$26888 ( \27231 , \27230 , \8050 );
not \U$26889 ( \27232 , \27230 );
and \U$26890 ( \27233 , \27232 , \8051 );
nor \U$26891 ( \27234 , \27231 , \27233 );
and \U$26892 ( \27235 , \27227 , \27234 );
and \U$26893 ( \27236 , \27219 , \27226 );
or \U$26894 ( \27237 , \27235 , \27236 );
and \U$26895 ( \27238 , \27212 , \27237 );
and \U$26896 ( \27239 , \27206 , \27211 );
nor \U$26897 ( \27240 , \27238 , \27239 );
not \U$26898 ( \27241 , \27240 );
and \U$26899 ( \27242 , \27204 , \27241 );
and \U$26900 ( \27243 , \27203 , \27240 );
and \U$26901 ( \27244 , \13882 , RI9871050_111);
and \U$26902 ( \27245 , RI9870c90_103, \13880 );
nor \U$26903 ( \27246 , \27244 , \27245 );
and \U$26904 ( \27247 , \27246 , \13359 );
not \U$26905 ( \27248 , \27246 );
and \U$26906 ( \27249 , \27248 , \13358 );
nor \U$26907 ( \27250 , \27247 , \27249 );
not \U$26908 ( \27251 , \27250 );
and \U$26909 ( \27252 , \15780 , RI9871320_117);
and \U$26910 ( \27253 , RI9873648_192, RI9871410_119);
nor \U$26911 ( \27254 , \27252 , \27253 );
not \U$26912 ( \27255 , \27254 );
not \U$26913 ( \27256 , RI9873558_190);
and \U$26914 ( \27257 , \27255 , \27256 );
and \U$26915 ( \27258 , \27254 , RI9873558_190);
nor \U$26916 ( \27259 , \27257 , \27258 );
not \U$26917 ( \27260 , \27259 );
and \U$26918 ( \27261 , \27251 , \27260 );
and \U$26919 ( \27262 , \27250 , \27259 );
and \U$26920 ( \27263 , \14937 , RI9871230_115);
and \U$26921 ( \27264 , RI9871140_113, \14935 );
nor \U$26922 ( \27265 , \27263 , \27264 );
and \U$26923 ( \27266 , \27265 , \14538 );
not \U$26924 ( \27267 , \27265 );
and \U$26925 ( \27268 , \27267 , \14539 );
nor \U$26926 ( \27269 , \27266 , \27268 );
nor \U$26927 ( \27270 , \27262 , \27269 );
nor \U$26928 ( \27271 , \27261 , \27270 );
not \U$26929 ( \27272 , \27271 );
and \U$26930 ( \27273 , \11696 , RI9870f60_109);
and \U$26931 ( \27274 , RI9870ab0_99, \11694 );
nor \U$26932 ( \27275 , \27273 , \27274 );
and \U$26933 ( \27276 , \27275 , \11702 );
not \U$26934 ( \27277 , \27275 );
and \U$26935 ( \27278 , \27277 , \10965 );
nor \U$26936 ( \27279 , \27276 , \27278 );
not \U$26937 ( \27280 , \27279 );
and \U$26938 ( \27281 , \12293 , RI9870d80_105);
and \U$26939 ( \27282 , RI98709c0_97, \12291 );
nor \U$26940 ( \27283 , \27281 , \27282 );
and \U$26941 ( \27284 , \27283 , \11686 );
not \U$26942 ( \27285 , \27283 );
and \U$26943 ( \27286 , \27285 , \11687 );
nor \U$26944 ( \27287 , \27284 , \27286 );
not \U$26945 ( \27288 , \27287 );
and \U$26946 ( \27289 , \27280 , \27288 );
and \U$26947 ( \27290 , \27287 , \27279 );
and \U$26948 ( \27291 , \13045 , RI9870e70_107);
and \U$26949 ( \27292 , RI9870ba0_101, \13043 );
nor \U$26950 ( \27293 , \27291 , \27292 );
and \U$26951 ( \27294 , \27293 , \12619 );
not \U$26952 ( \27295 , \27293 );
and \U$26953 ( \27296 , \27295 , \13047 );
nor \U$26954 ( \27297 , \27294 , \27296 );
nor \U$26955 ( \27298 , \27290 , \27297 );
nor \U$26956 ( \27299 , \27289 , \27298 );
not \U$26957 ( \27300 , \27299 );
and \U$26958 ( \27301 , \27272 , \27300 );
and \U$26959 ( \27302 , \27299 , \27271 );
and \U$26960 ( \27303 , \9237 , RI986fd90_71);
and \U$26961 ( \27304 , RI986fca0_69, \9235 );
nor \U$26962 ( \27305 , \27303 , \27304 );
and \U$26963 ( \27306 , \27305 , \8836 );
not \U$26964 ( \27307 , \27305 );
and \U$26965 ( \27308 , \27307 , \9241 );
nor \U$26966 ( \27309 , \27306 , \27308 );
not \U$26967 ( \27310 , \27309 );
and \U$26968 ( \27311 , \9505 , RI986ff70_75);
and \U$26969 ( \27312 , RI986fe80_73, \9503 );
nor \U$26970 ( \27313 , \27311 , \27312 );
and \U$26971 ( \27314 , \27313 , \9513 );
not \U$26972 ( \27315 , \27313 );
and \U$26973 ( \27316 , \27315 , \9510 );
nor \U$26974 ( \27317 , \27314 , \27316 );
not \U$26975 ( \27318 , \27317 );
and \U$26976 ( \27319 , \27310 , \27318 );
and \U$26977 ( \27320 , \27317 , \27309 );
and \U$26978 ( \27321 , \10424 , RI9870060_77);
and \U$26979 ( \27322 , RI9870150_79, \10422 );
nor \U$26980 ( \27323 , \27321 , \27322 );
and \U$26981 ( \27324 , \27323 , \10428 );
not \U$26982 ( \27325 , \27323 );
and \U$26983 ( \27326 , \27325 , \9840 );
nor \U$26984 ( \27327 , \27324 , \27326 );
nor \U$26985 ( \27328 , \27320 , \27327 );
nor \U$26986 ( \27329 , \27319 , \27328 );
nor \U$26987 ( \27330 , \27302 , \27329 );
nor \U$26988 ( \27331 , \27301 , \27330 );
nor \U$26989 ( \27332 , \27243 , \27331 );
nor \U$26990 ( \27333 , \27242 , \27332 );
xor \U$26991 ( \27334 , \26855 , \26861 );
xor \U$26992 ( \27335 , \27334 , \26888 );
or \U$26993 ( \27336 , \27333 , \27335 );
not \U$26994 ( \27337 , \27335 );
not \U$26995 ( \27338 , \27333 );
or \U$26996 ( \27339 , \27337 , \27338 );
xor \U$26997 ( \27340 , \26869 , \26877 );
xor \U$26998 ( \27341 , \27340 , \26885 );
xor \U$26999 ( \27342 , \26657 , \26682 );
xor \U$27000 ( \27343 , \27342 , \26685 );
and \U$27001 ( \27344 , \27341 , \27343 );
xor \U$27002 ( \27345 , \26789 , \26791 );
xor \U$27003 ( \27346 , \27345 , \26819 );
xor \U$27004 ( \27347 , \26657 , \26682 );
xor \U$27005 ( \27348 , \27347 , \26685 );
and \U$27006 ( \27349 , \27346 , \27348 );
and \U$27007 ( \27350 , \27341 , \27346 );
or \U$27008 ( \27351 , \27344 , \27349 , \27350 );
nand \U$27009 ( \27352 , \27339 , \27351 );
nand \U$27010 ( \27353 , \27336 , \27352 );
nand \U$27011 ( \27354 , \27190 , \27353 );
nand \U$27012 ( \27355 , \27189 , \27354 );
and \U$27013 ( \27356 , \27183 , \27355 );
and \U$27014 ( \27357 , \27180 , \27182 );
nor \U$27015 ( \27358 , \27356 , \27357 );
or \U$27016 ( \27359 , \27178 , \27358 );
xnor \U$27017 ( \27360 , \27358 , \27178 );
xor \U$27018 ( \27361 , \27180 , \27182 );
xor \U$27019 ( \27362 , \27361 , \27355 );
xnor \U$27020 ( \27363 , \27353 , \27187 );
not \U$27021 ( \27364 , \27363 );
not \U$27022 ( \27365 , \27184 );
and \U$27023 ( \27366 , \27364 , \27365 );
and \U$27024 ( \27367 , \27363 , \27184 );
nor \U$27025 ( \27368 , \27366 , \27367 );
not \U$27026 ( \27369 , \27333 );
not \U$27027 ( \27370 , \27351 );
or \U$27028 ( \27371 , \27369 , \27370 );
or \U$27029 ( \27372 , \27351 , \27333 );
nand \U$27030 ( \27373 , \27371 , \27372 );
not \U$27031 ( \27374 , \27373 );
not \U$27032 ( \27375 , \27335 );
and \U$27033 ( \27376 , \27374 , \27375 );
and \U$27034 ( \27377 , \27373 , \27335 );
nor \U$27035 ( \27378 , \27376 , \27377 );
not \U$27036 ( \27379 , \27378 );
xor \U$27037 ( \27380 , \26688 , \26761 );
xor \U$27038 ( \27381 , \27380 , \26822 );
nand \U$27039 ( \27382 , \27379 , \27381 );
or \U$27040 ( \27383 , \27368 , \27382 );
not \U$27041 ( \27384 , \27382 );
not \U$27042 ( \27385 , \27368 );
or \U$27043 ( \27386 , \27384 , \27385 );
not \U$27044 ( \27387 , \27240 );
xor \U$27045 ( \27388 , \27331 , \27203 );
not \U$27046 ( \27389 , \27388 );
or \U$27047 ( \27390 , \27387 , \27389 );
or \U$27048 ( \27391 , \27388 , \27240 );
nand \U$27049 ( \27392 , \27390 , \27391 );
xor \U$27050 ( \27393 , \26657 , \26682 );
xor \U$27051 ( \27394 , \27393 , \26685 );
xor \U$27052 ( \27395 , \27341 , \27346 );
xor \U$27053 ( \27396 , \27394 , \27395 );
and \U$27054 ( \27397 , \27392 , \27396 );
xor \U$27055 ( \27398 , \26608 , \26614 );
xor \U$27056 ( \27399 , \27398 , \26617 );
xor \U$27057 ( \27400 , \26606 , \26627 );
xor \U$27058 ( \27401 , \27399 , \27400 );
xor \U$27059 ( \27402 , \27397 , \27401 );
and \U$27060 ( \27403 , \12293 , RI9870ab0_99);
and \U$27061 ( \27404 , RI9870d80_105, \12291 );
nor \U$27062 ( \27405 , \27403 , \27404 );
and \U$27063 ( \27406 , \27405 , \11687 );
not \U$27064 ( \27407 , \27405 );
and \U$27065 ( \27408 , \27407 , \11686 );
nor \U$27066 ( \27409 , \27406 , \27408 );
and \U$27067 ( \27410 , \13045 , RI98709c0_97);
and \U$27068 ( \27411 , RI9870e70_107, \13043 );
nor \U$27069 ( \27412 , \27410 , \27411 );
and \U$27070 ( \27413 , \27412 , \13047 );
not \U$27071 ( \27414 , \27412 );
and \U$27072 ( \27415 , \27414 , \12619 );
nor \U$27073 ( \27416 , \27413 , \27415 );
xor \U$27074 ( \27417 , \27409 , \27416 );
and \U$27075 ( \27418 , \13882 , RI9870ba0_101);
and \U$27076 ( \27419 , RI9871050_111, \13880 );
nor \U$27077 ( \27420 , \27418 , \27419 );
and \U$27078 ( \27421 , \27420 , \13358 );
not \U$27079 ( \27422 , \27420 );
and \U$27080 ( \27423 , \27422 , \13359 );
nor \U$27081 ( \27424 , \27421 , \27423 );
and \U$27082 ( \27425 , \27417 , \27424 );
and \U$27083 ( \27426 , \27409 , \27416 );
or \U$27084 ( \27427 , \27425 , \27426 );
not \U$27085 ( \27428 , RI9873558_190);
and \U$27086 ( \27429 , \15780 , RI9871140_113);
and \U$27087 ( \27430 , RI9873648_192, RI9871320_117);
nor \U$27088 ( \27431 , \27429 , \27430 );
not \U$27089 ( \27432 , \27431 );
or \U$27090 ( \27433 , \27428 , \27432 );
or \U$27091 ( \27434 , \27431 , RI9873558_190);
nand \U$27092 ( \27435 , \27433 , \27434 );
xor \U$27093 ( \27436 , \27435 , \5885 );
and \U$27094 ( \27437 , \14937 , RI9870c90_103);
and \U$27095 ( \27438 , RI9871230_115, \14935 );
nor \U$27096 ( \27439 , \27437 , \27438 );
and \U$27097 ( \27440 , \27439 , \14539 );
not \U$27098 ( \27441 , \27439 );
and \U$27099 ( \27442 , \27441 , \14538 );
nor \U$27100 ( \27443 , \27440 , \27442 );
and \U$27101 ( \27444 , \27436 , \27443 );
and \U$27102 ( \27445 , \27435 , \5885 );
or \U$27103 ( \27446 , \27444 , \27445 );
xor \U$27104 ( \27447 , \27427 , \27446 );
and \U$27105 ( \27448 , \10424 , RI986fe80_73);
and \U$27106 ( \27449 , RI9870060_77, \10422 );
nor \U$27107 ( \27450 , \27448 , \27449 );
and \U$27108 ( \27451 , \27450 , \9840 );
not \U$27109 ( \27452 , \27450 );
and \U$27110 ( \27453 , \27452 , \10428 );
nor \U$27111 ( \27454 , \27451 , \27453 );
and \U$27112 ( \27455 , \9505 , RI986fca0_69);
and \U$27113 ( \27456 , RI986ff70_75, \9503 );
nor \U$27114 ( \27457 , \27455 , \27456 );
and \U$27115 ( \27458 , \27457 , \9510 );
not \U$27116 ( \27459 , \27457 );
and \U$27117 ( \27460 , \27459 , \9513 );
nor \U$27118 ( \27461 , \27458 , \27460 );
xor \U$27119 ( \27462 , \27454 , \27461 );
and \U$27120 ( \27463 , \11696 , RI9870150_79);
and \U$27121 ( \27464 , RI9870f60_109, \11694 );
nor \U$27122 ( \27465 , \27463 , \27464 );
and \U$27123 ( \27466 , \27465 , \10965 );
not \U$27124 ( \27467 , \27465 );
and \U$27125 ( \27468 , \27467 , \11702 );
nor \U$27126 ( \27469 , \27466 , \27468 );
and \U$27127 ( \27470 , \27462 , \27469 );
and \U$27128 ( \27471 , \27454 , \27461 );
or \U$27129 ( \27472 , \27470 , \27471 );
and \U$27130 ( \27473 , \27447 , \27472 );
and \U$27131 ( \27474 , \27427 , \27446 );
or \U$27132 ( \27475 , \27473 , \27474 );
and \U$27133 ( \27476 , \6453 , RI9870510_87);
and \U$27134 ( \27477 , RI9870330_83, \6451 );
nor \U$27135 ( \27478 , \27476 , \27477 );
and \U$27136 ( \27479 , \27478 , \6190 );
not \U$27137 ( \27480 , \27478 );
and \U$27138 ( \27481 , \27480 , \6180 );
nor \U$27139 ( \27482 , \27479 , \27481 );
nand \U$27140 ( \27483 , RI9870420_85, \5879 );
and \U$27141 ( \27484 , \27483 , \5594 );
not \U$27142 ( \27485 , \27483 );
and \U$27143 ( \27486 , \27485 , \5885 );
nor \U$27144 ( \27487 , \27484 , \27486 );
xor \U$27145 ( \27488 , \27482 , \27487 );
and \U$27146 ( \27489 , \7079 , RI9870240_81);
and \U$27147 ( \27490 , RI98706f0_91, \7077 );
nor \U$27148 ( \27491 , \27489 , \27490 );
and \U$27149 ( \27492 , \27491 , \6710 );
not \U$27150 ( \27493 , \27491 );
and \U$27151 ( \27494 , \27493 , \6709 );
nor \U$27152 ( \27495 , \27492 , \27494 );
and \U$27153 ( \27496 , \27488 , \27495 );
and \U$27154 ( \27497 , \27482 , \27487 );
or \U$27155 ( \27498 , \27496 , \27497 );
and \U$27156 ( \27499 , \6453 , RI9870330_83);
and \U$27157 ( \27500 , RI9870240_81, \6451 );
nor \U$27158 ( \27501 , \27499 , \27500 );
and \U$27159 ( \27502 , \27501 , \6190 );
not \U$27160 ( \27503 , \27501 );
and \U$27161 ( \27504 , \27503 , \6705 );
nor \U$27162 ( \27505 , \27502 , \27504 );
xor \U$27163 ( \27506 , \27498 , \27505 );
and \U$27164 ( \27507 , \9237 , RI986fbb0_67);
and \U$27165 ( \27508 , RI986fd90_71, \9235 );
nor \U$27166 ( \27509 , \27507 , \27508 );
and \U$27167 ( \27510 , \27509 , \9241 );
not \U$27168 ( \27511 , \27509 );
and \U$27169 ( \27512 , \27511 , \8836 );
nor \U$27170 ( \27513 , \27510 , \27512 );
and \U$27171 ( \27514 , \7729 , RI9870600_89);
and \U$27172 ( \27515 , RI98708d0_95, \7727 );
nor \U$27173 ( \27516 , \27514 , \27515 );
and \U$27174 ( \27517 , \27516 , \7480 );
not \U$27175 ( \27518 , \27516 );
and \U$27176 ( \27519 , \27518 , \7733 );
nor \U$27177 ( \27520 , \27517 , \27519 );
xor \U$27178 ( \27521 , \27513 , \27520 );
and \U$27179 ( \27522 , \8486 , RI98707e0_93);
and \U$27180 ( \27523 , RI986fac0_65, \8484 );
nor \U$27181 ( \27524 , \27522 , \27523 );
and \U$27182 ( \27525 , \27524 , \8050 );
not \U$27183 ( \27526 , \27524 );
and \U$27184 ( \27527 , \27526 , \8051 );
nor \U$27185 ( \27528 , \27525 , \27527 );
and \U$27186 ( \27529 , \27521 , \27528 );
and \U$27187 ( \27530 , \27513 , \27520 );
or \U$27188 ( \27531 , \27529 , \27530 );
and \U$27189 ( \27532 , \27506 , \27531 );
and \U$27190 ( \27533 , \27498 , \27505 );
or \U$27191 ( \27534 , \27532 , \27533 );
xor \U$27192 ( \27535 , \27475 , \27534 );
and \U$27193 ( \27536 , \5881 , RI9870420_85);
and \U$27194 ( \27537 , RI9870510_87, \5879 );
nor \U$27195 ( \27538 , \27536 , \27537 );
and \U$27196 ( \27539 , \27538 , \5594 );
not \U$27197 ( \27540 , \27538 );
and \U$27198 ( \27541 , \27540 , \5885 );
nor \U$27199 ( \27542 , \27539 , \27541 );
xor \U$27200 ( \27543 , \27219 , \27226 );
xor \U$27201 ( \27544 , \27543 , \27234 );
and \U$27202 ( \27545 , \27542 , \27544 );
not \U$27203 ( \27546 , \27309 );
xor \U$27204 ( \27547 , \27317 , \27327 );
not \U$27205 ( \27548 , \27547 );
or \U$27206 ( \27549 , \27546 , \27548 );
or \U$27207 ( \27550 , \27547 , \27309 );
nand \U$27208 ( \27551 , \27549 , \27550 );
xor \U$27209 ( \27552 , \27219 , \27226 );
xor \U$27210 ( \27553 , \27552 , \27234 );
and \U$27211 ( \27554 , \27551 , \27553 );
and \U$27212 ( \27555 , \27542 , \27551 );
or \U$27213 ( \27556 , \27545 , \27554 , \27555 );
and \U$27214 ( \27557 , \27535 , \27556 );
and \U$27215 ( \27558 , \27475 , \27534 );
or \U$27216 ( \27559 , \27557 , \27558 );
xor \U$27217 ( \27560 , \26713 , \26732 );
xor \U$27218 ( \27561 , \27560 , \26758 );
xor \U$27219 ( \27562 , \27559 , \27561 );
xor \U$27220 ( \27563 , \27206 , \27211 );
xor \U$27221 ( \27564 , \27563 , \27237 );
xor \U$27222 ( \27565 , \26721 , \5322 );
xor \U$27223 ( \27566 , \27565 , \26729 );
xor \U$27224 ( \27567 , \27564 , \27566 );
xor \U$27225 ( \27568 , \26695 , \26702 );
xor \U$27226 ( \27569 , \27568 , \26710 );
xor \U$27227 ( \27570 , \27192 , \27197 );
xor \U$27228 ( \27571 , \27569 , \27570 );
and \U$27229 ( \27572 , \27567 , \27571 );
and \U$27230 ( \27573 , \27564 , \27566 );
or \U$27231 ( \27574 , \27572 , \27573 );
and \U$27232 ( \27575 , \27562 , \27574 );
and \U$27233 ( \27576 , \27559 , \27561 );
or \U$27234 ( \27577 , \27575 , \27576 );
and \U$27235 ( \27578 , \27402 , \27577 );
and \U$27236 ( \27579 , \27397 , \27401 );
or \U$27237 ( \27580 , \27578 , \27579 );
nand \U$27238 ( \27581 , \27386 , \27580 );
nand \U$27239 ( \27582 , \27383 , \27581 );
and \U$27240 ( \27583 , \27362 , \27582 );
xor \U$27241 ( \27584 , \27582 , \27362 );
not \U$27242 ( \27585 , \27381 );
not \U$27243 ( \27586 , \27378 );
or \U$27244 ( \27587 , \27585 , \27586 );
or \U$27245 ( \27588 , \27378 , \27381 );
nand \U$27246 ( \27589 , \27587 , \27588 );
xor \U$27247 ( \27590 , \27397 , \27401 );
xor \U$27248 ( \27591 , \27590 , \27577 );
xor \U$27249 ( \27592 , \27589 , \27591 );
xor \U$27250 ( \27593 , \27392 , \27396 );
not \U$27251 ( \27594 , \27279 );
xor \U$27252 ( \27595 , \27287 , \27297 );
not \U$27253 ( \27596 , \27595 );
or \U$27254 ( \27597 , \27594 , \27596 );
or \U$27255 ( \27598 , \27595 , \27279 );
nand \U$27256 ( \27599 , \27597 , \27598 );
not \U$27257 ( \27600 , \27250 );
xor \U$27258 ( \27601 , \27259 , \27269 );
not \U$27259 ( \27602 , \27601 );
or \U$27260 ( \27603 , \27600 , \27602 );
or \U$27261 ( \27604 , \27601 , \27250 );
nand \U$27262 ( \27605 , \27603 , \27604 );
xor \U$27263 ( \27606 , \27599 , \27605 );
xor \U$27264 ( \27607 , \27219 , \27226 );
xor \U$27265 ( \27608 , \27607 , \27234 );
xor \U$27266 ( \27609 , \27542 , \27551 );
xor \U$27267 ( \27610 , \27608 , \27609 );
and \U$27268 ( \27611 , \27606 , \27610 );
and \U$27269 ( \27612 , \27599 , \27605 );
or \U$27270 ( \27613 , \27611 , \27612 );
not \U$27271 ( \27614 , \27299 );
xor \U$27272 ( \27615 , \27271 , \27329 );
not \U$27273 ( \27616 , \27615 );
or \U$27274 ( \27617 , \27614 , \27616 );
or \U$27275 ( \27618 , \27615 , \27299 );
nand \U$27276 ( \27619 , \27617 , \27618 );
xor \U$27277 ( \27620 , \27613 , \27619 );
xor \U$27278 ( \27621 , \27482 , \27487 );
xor \U$27279 ( \27622 , \27621 , \27495 );
and \U$27280 ( \27623 , \7079 , RI9870330_83);
and \U$27281 ( \27624 , RI9870240_81, \7077 );
nor \U$27282 ( \27625 , \27623 , \27624 );
and \U$27283 ( \27626 , \27625 , \6710 );
not \U$27284 ( \27627 , \27625 );
and \U$27285 ( \27628 , \27627 , \6709 );
nor \U$27286 ( \27629 , \27626 , \27628 );
and \U$27287 ( \27630 , \7729 , RI98706f0_91);
and \U$27288 ( \27631 , RI9870600_89, \7727 );
nor \U$27289 ( \27632 , \27630 , \27631 );
and \U$27290 ( \27633 , \27632 , \7480 );
not \U$27291 ( \27634 , \27632 );
and \U$27292 ( \27635 , \27634 , \7733 );
nor \U$27293 ( \27636 , \27633 , \27635 );
xor \U$27294 ( \27637 , \27629 , \27636 );
and \U$27295 ( \27638 , \8486 , RI98708d0_95);
and \U$27296 ( \27639 , RI98707e0_93, \8484 );
nor \U$27297 ( \27640 , \27638 , \27639 );
and \U$27298 ( \27641 , \27640 , \8050 );
not \U$27299 ( \27642 , \27640 );
and \U$27300 ( \27643 , \27642 , \8051 );
nor \U$27301 ( \27644 , \27641 , \27643 );
and \U$27302 ( \27645 , \27637 , \27644 );
and \U$27303 ( \27646 , \27629 , \27636 );
or \U$27304 ( \27647 , \27645 , \27646 );
xor \U$27305 ( \27648 , \27622 , \27647 );
xor \U$27306 ( \27649 , \27513 , \27520 );
xor \U$27307 ( \27650 , \27649 , \27528 );
and \U$27308 ( \27651 , \27648 , \27650 );
and \U$27309 ( \27652 , \27622 , \27647 );
or \U$27310 ( \27653 , \27651 , \27652 );
and \U$27311 ( \27654 , \11696 , RI9870060_77);
and \U$27312 ( \27655 , RI9870150_79, \11694 );
nor \U$27313 ( \27656 , \27654 , \27655 );
and \U$27314 ( \27657 , \27656 , \11702 );
not \U$27315 ( \27658 , \27656 );
and \U$27316 ( \27659 , \27658 , \10965 );
nor \U$27317 ( \27660 , \27657 , \27659 );
and \U$27318 ( \27661 , \12293 , RI9870f60_109);
and \U$27319 ( \27662 , RI9870ab0_99, \12291 );
nor \U$27320 ( \27663 , \27661 , \27662 );
and \U$27321 ( \27664 , \27663 , \11686 );
not \U$27322 ( \27665 , \27663 );
and \U$27323 ( \27666 , \27665 , \11687 );
nor \U$27324 ( \27667 , \27664 , \27666 );
or \U$27325 ( \27668 , \27660 , \27667 );
not \U$27326 ( \27669 , \27667 );
not \U$27327 ( \27670 , \27660 );
or \U$27328 ( \27671 , \27669 , \27670 );
and \U$27329 ( \27672 , \13045 , RI9870d80_105);
and \U$27330 ( \27673 , RI98709c0_97, \13043 );
nor \U$27331 ( \27674 , \27672 , \27673 );
and \U$27332 ( \27675 , \27674 , \13047 );
not \U$27333 ( \27676 , \27674 );
and \U$27334 ( \27677 , \27676 , \12619 );
nor \U$27335 ( \27678 , \27675 , \27677 );
nand \U$27336 ( \27679 , \27671 , \27678 );
nand \U$27337 ( \27680 , \27668 , \27679 );
and \U$27338 ( \27681 , \13882 , RI9870e70_107);
and \U$27339 ( \27682 , RI9870ba0_101, \13880 );
nor \U$27340 ( \27683 , \27681 , \27682 );
and \U$27341 ( \27684 , \27683 , \13359 );
not \U$27342 ( \27685 , \27683 );
and \U$27343 ( \27686 , \27685 , \13358 );
nor \U$27344 ( \27687 , \27684 , \27686 );
and \U$27345 ( \27688 , \15780 , RI9871230_115);
and \U$27346 ( \27689 , RI9873648_192, RI9871140_113);
nor \U$27347 ( \27690 , \27688 , \27689 );
not \U$27348 ( \27691 , \27690 );
not \U$27349 ( \27692 , RI9873558_190);
and \U$27350 ( \27693 , \27691 , \27692 );
and \U$27351 ( \27694 , \27690 , RI9873558_190);
nor \U$27352 ( \27695 , \27693 , \27694 );
or \U$27353 ( \27696 , \27687 , \27695 );
not \U$27354 ( \27697 , \27695 );
not \U$27355 ( \27698 , \27687 );
or \U$27356 ( \27699 , \27697 , \27698 );
and \U$27357 ( \27700 , \14937 , RI9871050_111);
and \U$27358 ( \27701 , RI9870c90_103, \14935 );
nor \U$27359 ( \27702 , \27700 , \27701 );
and \U$27360 ( \27703 , \27702 , \14539 );
not \U$27361 ( \27704 , \27702 );
and \U$27362 ( \27705 , \27704 , \14538 );
nor \U$27363 ( \27706 , \27703 , \27705 );
nand \U$27364 ( \27707 , \27699 , \27706 );
nand \U$27365 ( \27708 , \27696 , \27707 );
xor \U$27366 ( \27709 , \27680 , \27708 );
and \U$27367 ( \27710 , \9505 , RI986fd90_71);
and \U$27368 ( \27711 , RI986fca0_69, \9503 );
nor \U$27369 ( \27712 , \27710 , \27711 );
and \U$27370 ( \27713 , \27712 , \9513 );
not \U$27371 ( \27714 , \27712 );
and \U$27372 ( \27715 , \27714 , \9510 );
nor \U$27373 ( \27716 , \27713 , \27715 );
and \U$27374 ( \27717 , \10424 , RI986ff70_75);
and \U$27375 ( \27718 , RI986fe80_73, \10422 );
nor \U$27376 ( \27719 , \27717 , \27718 );
and \U$27377 ( \27720 , \27719 , \10428 );
not \U$27378 ( \27721 , \27719 );
and \U$27379 ( \27722 , \27721 , \9840 );
nor \U$27380 ( \27723 , \27720 , \27722 );
xor \U$27381 ( \27724 , \27716 , \27723 );
and \U$27382 ( \27725 , \9237 , RI986fac0_65);
and \U$27383 ( \27726 , RI986fbb0_67, \9235 );
nor \U$27384 ( \27727 , \27725 , \27726 );
and \U$27385 ( \27728 , \27727 , \8836 );
not \U$27386 ( \27729 , \27727 );
and \U$27387 ( \27730 , \27729 , \9241 );
nor \U$27388 ( \27731 , \27728 , \27730 );
and \U$27389 ( \27732 , \27724 , \27731 );
and \U$27390 ( \27733 , \27716 , \27723 );
nor \U$27391 ( \27734 , \27732 , \27733 );
and \U$27392 ( \27735 , \27709 , \27734 );
and \U$27393 ( \27736 , \27680 , \27708 );
or \U$27394 ( \27737 , \27735 , \27736 );
xor \U$27395 ( \27738 , \27653 , \27737 );
xor \U$27396 ( \27739 , \27454 , \27461 );
xor \U$27397 ( \27740 , \27739 , \27469 );
xor \U$27398 ( \27741 , \27435 , \5885 );
xor \U$27399 ( \27742 , \27741 , \27443 );
and \U$27400 ( \27743 , \27740 , \27742 );
xor \U$27401 ( \27744 , \27409 , \27416 );
xor \U$27402 ( \27745 , \27744 , \27424 );
xor \U$27403 ( \27746 , \27435 , \5885 );
xor \U$27404 ( \27747 , \27746 , \27443 );
and \U$27405 ( \27748 , \27745 , \27747 );
and \U$27406 ( \27749 , \27740 , \27745 );
or \U$27407 ( \27750 , \27743 , \27748 , \27749 );
and \U$27408 ( \27751 , \27738 , \27750 );
and \U$27409 ( \27752 , \27653 , \27737 );
or \U$27410 ( \27753 , \27751 , \27752 );
and \U$27411 ( \27754 , \27620 , \27753 );
and \U$27412 ( \27755 , \27613 , \27619 );
or \U$27413 ( \27756 , \27754 , \27755 );
xor \U$27414 ( \27757 , \27593 , \27756 );
xor \U$27415 ( \27758 , \27559 , \27561 );
xor \U$27416 ( \27759 , \27758 , \27574 );
and \U$27417 ( \27760 , \27757 , \27759 );
and \U$27418 ( \27761 , \27593 , \27756 );
or \U$27419 ( \27762 , \27760 , \27761 );
xor \U$27420 ( \27763 , \27592 , \27762 );
xor \U$27421 ( \27764 , \27475 , \27534 );
xor \U$27422 ( \27765 , \27764 , \27556 );
xor \U$27423 ( \27766 , \27613 , \27619 );
xor \U$27424 ( \27767 , \27766 , \27753 );
and \U$27425 ( \27768 , \27765 , \27767 );
not \U$27426 ( \27769 , \27768 );
xor \U$27427 ( \27770 , \27593 , \27756 );
xor \U$27428 ( \27771 , \27770 , \27759 );
not \U$27429 ( \27772 , \27771 );
or \U$27430 ( \27773 , \27769 , \27772 );
or \U$27431 ( \27774 , \27771 , \27768 );
and \U$27432 ( \27775 , \13882 , RI98709c0_97);
and \U$27433 ( \27776 , RI9870e70_107, \13880 );
nor \U$27434 ( \27777 , \27775 , \27776 );
and \U$27435 ( \27778 , \27777 , \13358 );
not \U$27436 ( \27779 , \27777 );
and \U$27437 ( \27780 , \27779 , \13359 );
nor \U$27438 ( \27781 , \27778 , \27780 );
and \U$27439 ( \27782 , \12293 , RI9870150_79);
and \U$27440 ( \27783 , RI9870f60_109, \12291 );
nor \U$27441 ( \27784 , \27782 , \27783 );
and \U$27442 ( \27785 , \27784 , \11687 );
not \U$27443 ( \27786 , \27784 );
and \U$27444 ( \27787 , \27786 , \11686 );
nor \U$27445 ( \27788 , \27785 , \27787 );
xor \U$27446 ( \27789 , \27781 , \27788 );
and \U$27447 ( \27790 , \13045 , RI9870ab0_99);
and \U$27448 ( \27791 , RI9870d80_105, \13043 );
nor \U$27449 ( \27792 , \27790 , \27791 );
and \U$27450 ( \27793 , \27792 , \13047 );
not \U$27451 ( \27794 , \27792 );
and \U$27452 ( \27795 , \27794 , \12619 );
nor \U$27453 ( \27796 , \27793 , \27795 );
and \U$27454 ( \27797 , \27789 , \27796 );
and \U$27455 ( \27798 , \27781 , \27788 );
or \U$27456 ( \27799 , \27797 , \27798 );
not \U$27457 ( \27800 , RI9873558_190);
and \U$27458 ( \27801 , \15780 , RI9870c90_103);
and \U$27459 ( \27802 , RI9873648_192, RI9871230_115);
nor \U$27460 ( \27803 , \27801 , \27802 );
not \U$27461 ( \27804 , \27803 );
or \U$27462 ( \27805 , \27800 , \27804 );
or \U$27463 ( \27806 , \27803 , RI9873558_190);
nand \U$27464 ( \27807 , \27805 , \27806 );
xor \U$27465 ( \27808 , \27807 , \6180 );
and \U$27466 ( \27809 , \14937 , RI9870ba0_101);
and \U$27467 ( \27810 , RI9871050_111, \14935 );
nor \U$27468 ( \27811 , \27809 , \27810 );
and \U$27469 ( \27812 , \27811 , \14539 );
not \U$27470 ( \27813 , \27811 );
and \U$27471 ( \27814 , \27813 , \14538 );
nor \U$27472 ( \27815 , \27812 , \27814 );
and \U$27473 ( \27816 , \27808 , \27815 );
and \U$27474 ( \27817 , \27807 , \6180 );
or \U$27475 ( \27818 , \27816 , \27817 );
xor \U$27476 ( \27819 , \27799 , \27818 );
and \U$27477 ( \27820 , \10424 , RI986fca0_69);
and \U$27478 ( \27821 , RI986ff70_75, \10422 );
nor \U$27479 ( \27822 , \27820 , \27821 );
and \U$27480 ( \27823 , \27822 , \9840 );
not \U$27481 ( \27824 , \27822 );
and \U$27482 ( \27825 , \27824 , \10428 );
nor \U$27483 ( \27826 , \27823 , \27825 );
and \U$27484 ( \27827 , \9505 , RI986fbb0_67);
and \U$27485 ( \27828 , RI986fd90_71, \9503 );
nor \U$27486 ( \27829 , \27827 , \27828 );
and \U$27487 ( \27830 , \27829 , \9510 );
not \U$27488 ( \27831 , \27829 );
and \U$27489 ( \27832 , \27831 , \9513 );
nor \U$27490 ( \27833 , \27830 , \27832 );
xor \U$27491 ( \27834 , \27826 , \27833 );
and \U$27492 ( \27835 , \11696 , RI986fe80_73);
and \U$27493 ( \27836 , RI9870060_77, \11694 );
nor \U$27494 ( \27837 , \27835 , \27836 );
and \U$27495 ( \27838 , \27837 , \10965 );
not \U$27496 ( \27839 , \27837 );
and \U$27497 ( \27840 , \27839 , \11702 );
nor \U$27498 ( \27841 , \27838 , \27840 );
and \U$27499 ( \27842 , \27834 , \27841 );
and \U$27500 ( \27843 , \27826 , \27833 );
or \U$27501 ( \27844 , \27842 , \27843 );
and \U$27502 ( \27845 , \27819 , \27844 );
and \U$27503 ( \27846 , \27799 , \27818 );
or \U$27504 ( \27847 , \27845 , \27846 );
and \U$27505 ( \27848 , \6453 , RI9870420_85);
and \U$27506 ( \27849 , RI9870510_87, \6451 );
nor \U$27507 ( \27850 , \27848 , \27849 );
and \U$27508 ( \27851 , \27850 , \6190 );
not \U$27509 ( \27852 , \27850 );
and \U$27510 ( \27853 , \27852 , \6705 );
nor \U$27511 ( \27854 , \27851 , \27853 );
not \U$27512 ( \27855 , \27854 );
nand \U$27513 ( \27856 , RI9870420_85, \6451 );
and \U$27514 ( \27857 , \27856 , \6190 );
not \U$27515 ( \27858 , \27856 );
and \U$27516 ( \27859 , \27858 , \6180 );
nor \U$27517 ( \27860 , \27857 , \27859 );
and \U$27518 ( \27861 , \7079 , RI9870510_87);
and \U$27519 ( \27862 , RI9870330_83, \7077 );
nor \U$27520 ( \27863 , \27861 , \27862 );
and \U$27521 ( \27864 , \27863 , \6710 );
not \U$27522 ( \27865 , \27863 );
and \U$27523 ( \27866 , \27865 , \6709 );
nor \U$27524 ( \27867 , \27864 , \27866 );
and \U$27525 ( \27868 , \27860 , \27867 );
not \U$27526 ( \27869 , \27868 );
or \U$27527 ( \27870 , \27855 , \27869 );
or \U$27528 ( \27871 , \27868 , \27854 );
and \U$27529 ( \27872 , \7729 , RI9870240_81);
and \U$27530 ( \27873 , RI98706f0_91, \7727 );
nor \U$27531 ( \27874 , \27872 , \27873 );
and \U$27532 ( \27875 , \27874 , \7480 );
not \U$27533 ( \27876 , \27874 );
and \U$27534 ( \27877 , \27876 , \7733 );
nor \U$27535 ( \27878 , \27875 , \27877 );
and \U$27536 ( \27879 , \8486 , RI9870600_89);
and \U$27537 ( \27880 , RI98708d0_95, \8484 );
nor \U$27538 ( \27881 , \27879 , \27880 );
and \U$27539 ( \27882 , \27881 , \8050 );
not \U$27540 ( \27883 , \27881 );
and \U$27541 ( \27884 , \27883 , \8051 );
nor \U$27542 ( \27885 , \27882 , \27884 );
xor \U$27543 ( \27886 , \27878 , \27885 );
and \U$27544 ( \27887 , \9237 , RI98707e0_93);
and \U$27545 ( \27888 , RI986fac0_65, \9235 );
nor \U$27546 ( \27889 , \27887 , \27888 );
and \U$27547 ( \27890 , \27889 , \9241 );
not \U$27548 ( \27891 , \27889 );
and \U$27549 ( \27892 , \27891 , \8836 );
nor \U$27550 ( \27893 , \27890 , \27892 );
and \U$27551 ( \27894 , \27886 , \27893 );
and \U$27552 ( \27895 , \27878 , \27885 );
or \U$27553 ( \27896 , \27894 , \27895 );
nand \U$27554 ( \27897 , \27871 , \27896 );
nand \U$27555 ( \27898 , \27870 , \27897 );
xor \U$27556 ( \27899 , \27847 , \27898 );
xor \U$27557 ( \27900 , \27716 , \27723 );
xor \U$27558 ( \27901 , \27900 , \27731 );
not \U$27559 ( \27902 , \27667 );
not \U$27560 ( \27903 , \27678 );
or \U$27561 ( \27904 , \27902 , \27903 );
or \U$27562 ( \27905 , \27667 , \27678 );
nand \U$27563 ( \27906 , \27904 , \27905 );
not \U$27564 ( \27907 , \27906 );
not \U$27565 ( \27908 , \27660 );
and \U$27566 ( \27909 , \27907 , \27908 );
and \U$27567 ( \27910 , \27906 , \27660 );
nor \U$27568 ( \27911 , \27909 , \27910 );
or \U$27569 ( \27912 , \27901 , \27911 );
not \U$27570 ( \27913 , \27911 );
not \U$27571 ( \27914 , \27901 );
or \U$27572 ( \27915 , \27913 , \27914 );
xor \U$27573 ( \27916 , \27629 , \27636 );
xor \U$27574 ( \27917 , \27916 , \27644 );
nand \U$27575 ( \27918 , \27915 , \27917 );
nand \U$27576 ( \27919 , \27912 , \27918 );
and \U$27577 ( \27920 , \27899 , \27919 );
and \U$27578 ( \27921 , \27847 , \27898 );
or \U$27579 ( \27922 , \27920 , \27921 );
xor \U$27580 ( \27923 , \27498 , \27505 );
xor \U$27581 ( \27924 , \27923 , \27531 );
xor \U$27582 ( \27925 , \27922 , \27924 );
xor \U$27583 ( \27926 , \27680 , \27708 );
xor \U$27584 ( \27927 , \27926 , \27734 );
xor \U$27585 ( \27928 , \27622 , \27647 );
xor \U$27586 ( \27929 , \27928 , \27650 );
and \U$27587 ( \27930 , \27927 , \27929 );
xor \U$27588 ( \27931 , \27435 , \5885 );
xor \U$27589 ( \27932 , \27931 , \27443 );
xor \U$27590 ( \27933 , \27740 , \27745 );
xor \U$27591 ( \27934 , \27932 , \27933 );
xor \U$27592 ( \27935 , \27622 , \27647 );
xor \U$27593 ( \27936 , \27935 , \27650 );
and \U$27594 ( \27937 , \27934 , \27936 );
and \U$27595 ( \27938 , \27927 , \27934 );
or \U$27596 ( \27939 , \27930 , \27937 , \27938 );
and \U$27597 ( \27940 , \27925 , \27939 );
and \U$27598 ( \27941 , \27922 , \27924 );
or \U$27599 ( \27942 , \27940 , \27941 );
xor \U$27600 ( \27943 , \27564 , \27566 );
xor \U$27601 ( \27944 , \27943 , \27571 );
xor \U$27602 ( \27945 , \27942 , \27944 );
xor \U$27603 ( \27946 , \27599 , \27605 );
xor \U$27604 ( \27947 , \27946 , \27610 );
xor \U$27605 ( \27948 , \27427 , \27446 );
xor \U$27606 ( \27949 , \27948 , \27472 );
xor \U$27607 ( \27950 , \27947 , \27949 );
xor \U$27608 ( \27951 , \27653 , \27737 );
xor \U$27609 ( \27952 , \27951 , \27750 );
and \U$27610 ( \27953 , \27950 , \27952 );
and \U$27611 ( \27954 , \27947 , \27949 );
or \U$27612 ( \27955 , \27953 , \27954 );
and \U$27613 ( \27956 , \27945 , \27955 );
and \U$27614 ( \27957 , \27942 , \27944 );
or \U$27615 ( \27958 , \27956 , \27957 );
nand \U$27616 ( \27959 , \27774 , \27958 );
nand \U$27617 ( \27960 , \27773 , \27959 );
and \U$27618 ( \27961 , \27763 , \27960 );
xor \U$27619 ( \27962 , \27960 , \27763 );
xor \U$27620 ( \27963 , \27947 , \27949 );
xor \U$27621 ( \27964 , \27963 , \27952 );
xor \U$27622 ( \27965 , \27622 , \27647 );
xor \U$27623 ( \27966 , \27965 , \27650 );
xor \U$27624 ( \27967 , \27927 , \27934 );
xor \U$27625 ( \27968 , \27966 , \27967 );
not \U$27626 ( \27969 , \27968 );
xnor \U$27627 ( \27970 , \27896 , \27868 );
not \U$27628 ( \27971 , \27970 );
not \U$27629 ( \27972 , \27854 );
and \U$27630 ( \27973 , \27971 , \27972 );
and \U$27631 ( \27974 , \27970 , \27854 );
nor \U$27632 ( \27975 , \27973 , \27974 );
not \U$27633 ( \27976 , \27695 );
not \U$27634 ( \27977 , \27706 );
or \U$27635 ( \27978 , \27976 , \27977 );
or \U$27636 ( \27979 , \27706 , \27695 );
nand \U$27637 ( \27980 , \27978 , \27979 );
not \U$27638 ( \27981 , \27980 );
not \U$27639 ( \27982 , \27687 );
and \U$27640 ( \27983 , \27981 , \27982 );
and \U$27641 ( \27984 , \27980 , \27687 );
nor \U$27642 ( \27985 , \27983 , \27984 );
xor \U$27643 ( \27986 , \27975 , \27985 );
not \U$27644 ( \27987 , \27911 );
not \U$27645 ( \27988 , \27917 );
or \U$27646 ( \27989 , \27987 , \27988 );
or \U$27647 ( \27990 , \27911 , \27917 );
nand \U$27648 ( \27991 , \27989 , \27990 );
not \U$27649 ( \27992 , \27991 );
not \U$27650 ( \27993 , \27901 );
and \U$27651 ( \27994 , \27992 , \27993 );
and \U$27652 ( \27995 , \27991 , \27901 );
nor \U$27653 ( \27996 , \27994 , \27995 );
and \U$27654 ( \27997 , \27986 , \27996 );
and \U$27655 ( \27998 , \27975 , \27985 );
or \U$27656 ( \27999 , \27997 , \27998 );
or \U$27657 ( \28000 , \27969 , \27999 );
not \U$27658 ( \28001 , \27999 );
not \U$27659 ( \28002 , \27969 );
or \U$27660 ( \28003 , \28001 , \28002 );
and \U$27661 ( \28004 , \7079 , RI9870420_85);
and \U$27662 ( \28005 , RI9870510_87, \7077 );
nor \U$27663 ( \28006 , \28004 , \28005 );
and \U$27664 ( \28007 , \28006 , \6710 );
not \U$27665 ( \28008 , \28006 );
and \U$27666 ( \28009 , \28008 , \6709 );
nor \U$27667 ( \28010 , \28007 , \28009 );
and \U$27668 ( \28011 , \7729 , RI9870330_83);
and \U$27669 ( \28012 , RI9870240_81, \7727 );
nor \U$27670 ( \28013 , \28011 , \28012 );
and \U$27671 ( \28014 , \28013 , \7480 );
not \U$27672 ( \28015 , \28013 );
and \U$27673 ( \28016 , \28015 , \7733 );
nor \U$27674 ( \28017 , \28014 , \28016 );
xor \U$27675 ( \28018 , \28010 , \28017 );
and \U$27676 ( \28019 , \8486 , RI98706f0_91);
and \U$27677 ( \28020 , RI9870600_89, \8484 );
nor \U$27678 ( \28021 , \28019 , \28020 );
and \U$27679 ( \28022 , \28021 , \8050 );
not \U$27680 ( \28023 , \28021 );
and \U$27681 ( \28024 , \28023 , \8051 );
nor \U$27682 ( \28025 , \28022 , \28024 );
and \U$27683 ( \28026 , \28018 , \28025 );
and \U$27684 ( \28027 , \28010 , \28017 );
or \U$27685 ( \28028 , \28026 , \28027 );
xor \U$27686 ( \28029 , \27860 , \27867 );
xor \U$27687 ( \28030 , \28028 , \28029 );
xor \U$27688 ( \28031 , \27878 , \27885 );
xor \U$27689 ( \28032 , \28031 , \27893 );
and \U$27690 ( \28033 , \28030 , \28032 );
and \U$27691 ( \28034 , \28028 , \28029 );
or \U$27692 ( \28035 , \28033 , \28034 );
and \U$27693 ( \28036 , \9505 , RI986fac0_65);
and \U$27694 ( \28037 , RI986fbb0_67, \9503 );
nor \U$27695 ( \28038 , \28036 , \28037 );
and \U$27696 ( \28039 , \28038 , \9510 );
not \U$27697 ( \28040 , \28038 );
and \U$27698 ( \28041 , \28040 , \9513 );
nor \U$27699 ( \28042 , \28039 , \28041 );
and \U$27700 ( \28043 , \9237 , RI98708d0_95);
and \U$27701 ( \28044 , RI98707e0_93, \9235 );
nor \U$27702 ( \28045 , \28043 , \28044 );
and \U$27703 ( \28046 , \28045 , \9241 );
not \U$27704 ( \28047 , \28045 );
and \U$27705 ( \28048 , \28047 , \8836 );
nor \U$27706 ( \28049 , \28046 , \28048 );
xor \U$27707 ( \28050 , \28042 , \28049 );
and \U$27708 ( \28051 , \10424 , RI986fd90_71);
and \U$27709 ( \28052 , RI986fca0_69, \10422 );
nor \U$27710 ( \28053 , \28051 , \28052 );
and \U$27711 ( \28054 , \28053 , \9840 );
not \U$27712 ( \28055 , \28053 );
and \U$27713 ( \28056 , \28055 , \10428 );
nor \U$27714 ( \28057 , \28054 , \28056 );
and \U$27715 ( \28058 , \28050 , \28057 );
and \U$27716 ( \28059 , \28042 , \28049 );
or \U$27717 ( \28060 , \28058 , \28059 );
and \U$27718 ( \28061 , \13882 , RI9870d80_105);
and \U$27719 ( \28062 , RI98709c0_97, \13880 );
nor \U$27720 ( \28063 , \28061 , \28062 );
and \U$27721 ( \28064 , \28063 , \13358 );
not \U$27722 ( \28065 , \28063 );
and \U$27723 ( \28066 , \28065 , \13359 );
nor \U$27724 ( \28067 , \28064 , \28066 );
not \U$27725 ( \28068 , RI9873558_190);
and \U$27726 ( \28069 , \15780 , RI9871050_111);
and \U$27727 ( \28070 , RI9873648_192, RI9870c90_103);
nor \U$27728 ( \28071 , \28069 , \28070 );
not \U$27729 ( \28072 , \28071 );
or \U$27730 ( \28073 , \28068 , \28072 );
or \U$27731 ( \28074 , \28071 , RI9873558_190);
nand \U$27732 ( \28075 , \28073 , \28074 );
xor \U$27733 ( \28076 , \28067 , \28075 );
and \U$27734 ( \28077 , \14937 , RI9870e70_107);
and \U$27735 ( \28078 , RI9870ba0_101, \14935 );
nor \U$27736 ( \28079 , \28077 , \28078 );
and \U$27737 ( \28080 , \28079 , \14539 );
not \U$27738 ( \28081 , \28079 );
and \U$27739 ( \28082 , \28081 , \14538 );
nor \U$27740 ( \28083 , \28080 , \28082 );
and \U$27741 ( \28084 , \28076 , \28083 );
and \U$27742 ( \28085 , \28067 , \28075 );
or \U$27743 ( \28086 , \28084 , \28085 );
xor \U$27744 ( \28087 , \28060 , \28086 );
and \U$27745 ( \28088 , \11696 , RI986ff70_75);
and \U$27746 ( \28089 , RI986fe80_73, \11694 );
nor \U$27747 ( \28090 , \28088 , \28089 );
and \U$27748 ( \28091 , \28090 , \10965 );
not \U$27749 ( \28092 , \28090 );
and \U$27750 ( \28093 , \28092 , \11702 );
nor \U$27751 ( \28094 , \28091 , \28093 );
and \U$27752 ( \28095 , \12293 , RI9870060_77);
and \U$27753 ( \28096 , RI9870150_79, \12291 );
nor \U$27754 ( \28097 , \28095 , \28096 );
and \U$27755 ( \28098 , \28097 , \11687 );
not \U$27756 ( \28099 , \28097 );
and \U$27757 ( \28100 , \28099 , \11686 );
nor \U$27758 ( \28101 , \28098 , \28100 );
xor \U$27759 ( \28102 , \28094 , \28101 );
and \U$27760 ( \28103 , \13045 , RI9870f60_109);
and \U$27761 ( \28104 , RI9870ab0_99, \13043 );
nor \U$27762 ( \28105 , \28103 , \28104 );
and \U$27763 ( \28106 , \28105 , \13047 );
not \U$27764 ( \28107 , \28105 );
and \U$27765 ( \28108 , \28107 , \12619 );
nor \U$27766 ( \28109 , \28106 , \28108 );
and \U$27767 ( \28110 , \28102 , \28109 );
and \U$27768 ( \28111 , \28094 , \28101 );
or \U$27769 ( \28112 , \28110 , \28111 );
and \U$27770 ( \28113 , \28087 , \28112 );
and \U$27771 ( \28114 , \28060 , \28086 );
or \U$27772 ( \28115 , \28113 , \28114 );
xor \U$27773 ( \28116 , \28035 , \28115 );
xor \U$27774 ( \28117 , \27826 , \27833 );
xor \U$27775 ( \28118 , \28117 , \27841 );
xor \U$27776 ( \28119 , \27781 , \27788 );
xor \U$27777 ( \28120 , \28119 , \27796 );
and \U$27778 ( \28121 , \28118 , \28120 );
xor \U$27779 ( \28122 , \27807 , \6180 );
xor \U$27780 ( \28123 , \28122 , \27815 );
xor \U$27781 ( \28124 , \27781 , \27788 );
xor \U$27782 ( \28125 , \28124 , \27796 );
and \U$27783 ( \28126 , \28123 , \28125 );
and \U$27784 ( \28127 , \28118 , \28123 );
or \U$27785 ( \28128 , \28121 , \28126 , \28127 );
and \U$27786 ( \28129 , \28116 , \28128 );
and \U$27787 ( \28130 , \28035 , \28115 );
or \U$27788 ( \28131 , \28129 , \28130 );
nand \U$27789 ( \28132 , \28003 , \28131 );
nand \U$27790 ( \28133 , \28000 , \28132 );
xor \U$27791 ( \28134 , \27922 , \27924 );
xor \U$27792 ( \28135 , \28134 , \27939 );
xor \U$27793 ( \28136 , \28133 , \28135 );
xor \U$27794 ( \28137 , \27964 , \28136 );
not \U$27795 ( \28138 , \28137 );
xor \U$27796 ( \28139 , \27847 , \27898 );
xor \U$27797 ( \28140 , \28139 , \27919 );
not \U$27798 ( \28141 , \28140 );
xor \U$27799 ( \28142 , \27975 , \27985 );
xor \U$27800 ( \28143 , \28142 , \27996 );
not \U$27801 ( \28144 , \28143 );
xor \U$27802 ( \28145 , \28035 , \28115 );
xor \U$27803 ( \28146 , \28145 , \28128 );
nand \U$27804 ( \28147 , \28144 , \28146 );
nand \U$27805 ( \28148 , \28141 , \28147 );
and \U$27806 ( \28149 , \9505 , RI98707e0_93);
and \U$27807 ( \28150 , RI986fac0_65, \9503 );
nor \U$27808 ( \28151 , \28149 , \28150 );
and \U$27809 ( \28152 , \28151 , \9510 );
not \U$27810 ( \28153 , \28151 );
and \U$27811 ( \28154 , \28153 , \9513 );
nor \U$27812 ( \28155 , \28152 , \28154 );
and \U$27813 ( \28156 , \10424 , RI986fbb0_67);
and \U$27814 ( \28157 , RI986fd90_71, \10422 );
nor \U$27815 ( \28158 , \28156 , \28157 );
and \U$27816 ( \28159 , \28158 , \9840 );
not \U$27817 ( \28160 , \28158 );
and \U$27818 ( \28161 , \28160 , \10428 );
nor \U$27819 ( \28162 , \28159 , \28161 );
xor \U$27820 ( \28163 , \28155 , \28162 );
and \U$27821 ( \28164 , \11696 , RI986fca0_69);
and \U$27822 ( \28165 , RI986ff70_75, \11694 );
nor \U$27823 ( \28166 , \28164 , \28165 );
and \U$27824 ( \28167 , \28166 , \10965 );
not \U$27825 ( \28168 , \28166 );
and \U$27826 ( \28169 , \28168 , \11702 );
nor \U$27827 ( \28170 , \28167 , \28169 );
and \U$27828 ( \28171 , \28163 , \28170 );
and \U$27829 ( \28172 , \28155 , \28162 );
or \U$27830 ( \28173 , \28171 , \28172 );
not \U$27831 ( \28174 , RI9873558_190);
and \U$27832 ( \28175 , \15780 , RI9870ba0_101);
and \U$27833 ( \28176 , RI9873648_192, RI9871050_111);
nor \U$27834 ( \28177 , \28175 , \28176 );
not \U$27835 ( \28178 , \28177 );
or \U$27836 ( \28179 , \28174 , \28178 );
or \U$27837 ( \28180 , \28177 , RI9873558_190);
nand \U$27838 ( \28181 , \28179 , \28180 );
xor \U$27839 ( \28182 , \28181 , \6709 );
and \U$27840 ( \28183 , \14937 , RI98709c0_97);
and \U$27841 ( \28184 , RI9870e70_107, \14935 );
nor \U$27842 ( \28185 , \28183 , \28184 );
and \U$27843 ( \28186 , \28185 , \14539 );
not \U$27844 ( \28187 , \28185 );
and \U$27845 ( \28188 , \28187 , \14538 );
nor \U$27846 ( \28189 , \28186 , \28188 );
and \U$27847 ( \28190 , \28182 , \28189 );
and \U$27848 ( \28191 , \28181 , \6709 );
or \U$27849 ( \28192 , \28190 , \28191 );
xor \U$27850 ( \28193 , \28173 , \28192 );
and \U$27851 ( \28194 , \13045 , RI9870150_79);
and \U$27852 ( \28195 , RI9870f60_109, \13043 );
nor \U$27853 ( \28196 , \28194 , \28195 );
and \U$27854 ( \28197 , \28196 , \12619 );
not \U$27855 ( \28198 , \28196 );
and \U$27856 ( \28199 , \28198 , \13047 );
nor \U$27857 ( \28200 , \28197 , \28199 );
and \U$27858 ( \28201 , \13882 , RI9870ab0_99);
and \U$27859 ( \28202 , RI9870d80_105, \13880 );
nor \U$27860 ( \28203 , \28201 , \28202 );
and \U$27861 ( \28204 , \28203 , \13359 );
not \U$27862 ( \28205 , \28203 );
and \U$27863 ( \28206 , \28205 , \13358 );
nor \U$27864 ( \28207 , \28204 , \28206 );
xor \U$27865 ( \28208 , \28200 , \28207 );
and \U$27866 ( \28209 , \12293 , RI986fe80_73);
and \U$27867 ( \28210 , RI9870060_77, \12291 );
nor \U$27868 ( \28211 , \28209 , \28210 );
and \U$27869 ( \28212 , \28211 , \11686 );
not \U$27870 ( \28213 , \28211 );
and \U$27871 ( \28214 , \28213 , \11687 );
nor \U$27872 ( \28215 , \28212 , \28214 );
and \U$27873 ( \28216 , \28208 , \28215 );
and \U$27874 ( \28217 , \28200 , \28207 );
nor \U$27875 ( \28218 , \28216 , \28217 );
and \U$27876 ( \28219 , \28193 , \28218 );
and \U$27877 ( \28220 , \28173 , \28192 );
or \U$27878 ( \28221 , \28219 , \28220 );
xor \U$27879 ( \28222 , \28094 , \28101 );
xor \U$27880 ( \28223 , \28222 , \28109 );
xor \U$27881 ( \28224 , \28067 , \28075 );
xor \U$27882 ( \28225 , \28224 , \28083 );
and \U$27883 ( \28226 , \28223 , \28225 );
xor \U$27884 ( \28227 , \28221 , \28226 );
and \U$27885 ( \28228 , \8486 , RI9870240_81);
and \U$27886 ( \28229 , RI98706f0_91, \8484 );
nor \U$27887 ( \28230 , \28228 , \28229 );
and \U$27888 ( \28231 , \28230 , \8050 );
not \U$27889 ( \28232 , \28230 );
and \U$27890 ( \28233 , \28232 , \8051 );
nor \U$27891 ( \28234 , \28231 , \28233 );
and \U$27892 ( \28235 , \7729 , RI9870510_87);
and \U$27893 ( \28236 , RI9870330_83, \7727 );
nor \U$27894 ( \28237 , \28235 , \28236 );
and \U$27895 ( \28238 , \28237 , \7480 );
not \U$27896 ( \28239 , \28237 );
and \U$27897 ( \28240 , \28239 , \7733 );
nor \U$27898 ( \28241 , \28238 , \28240 );
xor \U$27899 ( \28242 , \28234 , \28241 );
and \U$27900 ( \28243 , \9237 , RI9870600_89);
and \U$27901 ( \28244 , RI98708d0_95, \9235 );
nor \U$27902 ( \28245 , \28243 , \28244 );
and \U$27903 ( \28246 , \28245 , \9241 );
not \U$27904 ( \28247 , \28245 );
and \U$27905 ( \28248 , \28247 , \8836 );
nor \U$27906 ( \28249 , \28246 , \28248 );
and \U$27907 ( \28250 , \28242 , \28249 );
and \U$27908 ( \28251 , \28234 , \28241 );
or \U$27909 ( \28252 , \28250 , \28251 );
xor \U$27910 ( \28253 , \28010 , \28017 );
xor \U$27911 ( \28254 , \28253 , \28025 );
and \U$27912 ( \28255 , \28252 , \28254 );
xor \U$27913 ( \28256 , \28042 , \28049 );
xor \U$27914 ( \28257 , \28256 , \28057 );
xor \U$27915 ( \28258 , \28010 , \28017 );
xor \U$27916 ( \28259 , \28258 , \28025 );
and \U$27917 ( \28260 , \28257 , \28259 );
and \U$27918 ( \28261 , \28252 , \28257 );
or \U$27919 ( \28262 , \28255 , \28260 , \28261 );
and \U$27920 ( \28263 , \28227 , \28262 );
and \U$27921 ( \28264 , \28221 , \28226 );
or \U$27922 ( \28265 , \28263 , \28264 );
xor \U$27923 ( \28266 , \27799 , \27818 );
xor \U$27924 ( \28267 , \28266 , \27844 );
xor \U$27925 ( \28268 , \28265 , \28267 );
xor \U$27926 ( \28269 , \28060 , \28086 );
xor \U$27927 ( \28270 , \28269 , \28112 );
xor \U$27928 ( \28271 , \28028 , \28029 );
xor \U$27929 ( \28272 , \28271 , \28032 );
and \U$27930 ( \28273 , \28270 , \28272 );
xor \U$27931 ( \28274 , \27781 , \27788 );
xor \U$27932 ( \28275 , \28274 , \27796 );
xor \U$27933 ( \28276 , \28118 , \28123 );
xor \U$27934 ( \28277 , \28275 , \28276 );
xor \U$27935 ( \28278 , \28028 , \28029 );
xor \U$27936 ( \28279 , \28278 , \28032 );
and \U$27937 ( \28280 , \28277 , \28279 );
and \U$27938 ( \28281 , \28270 , \28277 );
or \U$27939 ( \28282 , \28273 , \28280 , \28281 );
and \U$27940 ( \28283 , \28268 , \28282 );
and \U$27941 ( \28284 , \28265 , \28267 );
or \U$27942 ( \28285 , \28283 , \28284 );
and \U$27943 ( \28286 , \28148 , \28285 );
not \U$27944 ( \28287 , \28147 );
and \U$27945 ( \28288 , \28140 , \28287 );
nor \U$27946 ( \28289 , \28286 , \28288 );
not \U$27947 ( \28290 , \28289 );
and \U$27948 ( \28291 , \28138 , \28290 );
and \U$27949 ( \28292 , \28137 , \28289 );
nor \U$27950 ( \28293 , \28291 , \28292 );
not \U$27951 ( \28294 , \27999 );
not \U$27952 ( \28295 , \28131 );
and \U$27953 ( \28296 , \28294 , \28295 );
and \U$27954 ( \28297 , \27999 , \28131 );
nor \U$27955 ( \28298 , \28296 , \28297 );
not \U$27956 ( \28299 , \28298 );
not \U$27957 ( \28300 , \27968 );
and \U$27958 ( \28301 , \28299 , \28300 );
and \U$27959 ( \28302 , \28298 , \27968 );
nor \U$27960 ( \28303 , \28301 , \28302 );
not \U$27961 ( \28304 , \28303 );
not \U$27962 ( \28305 , \28140 );
not \U$27963 ( \28306 , \28285 );
not \U$27964 ( \28307 , \28147 );
and \U$27965 ( \28308 , \28306 , \28307 );
and \U$27966 ( \28309 , \28285 , \28147 );
nor \U$27967 ( \28310 , \28308 , \28309 );
not \U$27968 ( \28311 , \28310 );
or \U$27969 ( \28312 , \28305 , \28311 );
or \U$27970 ( \28313 , \28310 , \28140 );
nand \U$27971 ( \28314 , \28312 , \28313 );
nand \U$27972 ( \28315 , \28304 , \28314 );
or \U$27973 ( \28316 , \28293 , \28315 );
xnor \U$27974 ( \28317 , \28315 , \28293 );
and \U$27975 ( \28318 , \9505 , RI98706f0_91);
and \U$27976 ( \28319 , RI9870600_89, \9503 );
nor \U$27977 ( \28320 , \28318 , \28319 );
and \U$27978 ( \28321 , \28320 , \9510 );
not \U$27979 ( \28322 , \28320 );
and \U$27980 ( \28323 , \28322 , \9513 );
nor \U$27981 ( \28324 , \28321 , \28323 );
and \U$27982 ( \28325 , \9237 , RI9870330_83);
and \U$27983 ( \28326 , RI9870240_81, \9235 );
nor \U$27984 ( \28327 , \28325 , \28326 );
and \U$27985 ( \28328 , \28327 , \9241 );
not \U$27986 ( \28329 , \28327 );
and \U$27987 ( \28330 , \28329 , \8836 );
nor \U$27988 ( \28331 , \28328 , \28330 );
xor \U$27989 ( \28332 , \28324 , \28331 );
and \U$27990 ( \28333 , \10424 , RI98708d0_95);
and \U$27991 ( \28334 , RI98707e0_93, \10422 );
nor \U$27992 ( \28335 , \28333 , \28334 );
and \U$27993 ( \28336 , \28335 , \9840 );
not \U$27994 ( \28337 , \28335 );
and \U$27995 ( \28338 , \28337 , \10428 );
nor \U$27996 ( \28339 , \28336 , \28338 );
and \U$27997 ( \28340 , \28332 , \28339 );
and \U$27998 ( \28341 , \28324 , \28331 );
or \U$27999 ( \28342 , \28340 , \28341 );
and \U$28000 ( \28343 , \13882 , RI9870060_77);
and \U$28001 ( \28344 , RI9870150_79, \13880 );
nor \U$28002 ( \28345 , \28343 , \28344 );
and \U$28003 ( \28346 , \28345 , \13358 );
not \U$28004 ( \28347 , \28345 );
and \U$28005 ( \28348 , \28347 , \13359 );
nor \U$28006 ( \28349 , \28346 , \28348 );
not \U$28007 ( \28350 , RI9873558_190);
and \U$28008 ( \28351 , \15780 , RI9870d80_105);
and \U$28009 ( \28352 , RI9873648_192, RI98709c0_97);
nor \U$28010 ( \28353 , \28351 , \28352 );
not \U$28011 ( \28354 , \28353 );
or \U$28012 ( \28355 , \28350 , \28354 );
or \U$28013 ( \28356 , \28353 , RI9873558_190);
nand \U$28014 ( \28357 , \28355 , \28356 );
xor \U$28015 ( \28358 , \28349 , \28357 );
and \U$28016 ( \28359 , \14937 , RI9870f60_109);
and \U$28017 ( \28360 , RI9870ab0_99, \14935 );
nor \U$28018 ( \28361 , \28359 , \28360 );
and \U$28019 ( \28362 , \28361 , \14539 );
not \U$28020 ( \28363 , \28361 );
and \U$28021 ( \28364 , \28363 , \14538 );
nor \U$28022 ( \28365 , \28362 , \28364 );
and \U$28023 ( \28366 , \28358 , \28365 );
and \U$28024 ( \28367 , \28349 , \28357 );
or \U$28025 ( \28368 , \28366 , \28367 );
xor \U$28026 ( \28369 , \28342 , \28368 );
and \U$28027 ( \28370 , \11696 , RI986fac0_65);
and \U$28028 ( \28371 , RI986fbb0_67, \11694 );
nor \U$28029 ( \28372 , \28370 , \28371 );
and \U$28030 ( \28373 , \28372 , \10965 );
not \U$28031 ( \28374 , \28372 );
and \U$28032 ( \28375 , \28374 , \11702 );
nor \U$28033 ( \28376 , \28373 , \28375 );
and \U$28034 ( \28377 , \12293 , RI986fd90_71);
and \U$28035 ( \28378 , RI986fca0_69, \12291 );
nor \U$28036 ( \28379 , \28377 , \28378 );
and \U$28037 ( \28380 , \28379 , \11687 );
not \U$28038 ( \28381 , \28379 );
and \U$28039 ( \28382 , \28381 , \11686 );
nor \U$28040 ( \28383 , \28380 , \28382 );
xor \U$28041 ( \28384 , \28376 , \28383 );
and \U$28042 ( \28385 , \13045 , RI986ff70_75);
and \U$28043 ( \28386 , RI986fe80_73, \13043 );
nor \U$28044 ( \28387 , \28385 , \28386 );
and \U$28045 ( \28388 , \28387 , \13047 );
not \U$28046 ( \28389 , \28387 );
and \U$28047 ( \28390 , \28389 , \12619 );
nor \U$28048 ( \28391 , \28388 , \28390 );
and \U$28049 ( \28392 , \28384 , \28391 );
and \U$28050 ( \28393 , \28376 , \28383 );
or \U$28051 ( \28394 , \28392 , \28393 );
and \U$28052 ( \28395 , \28369 , \28394 );
and \U$28053 ( \28396 , \28342 , \28368 );
nor \U$28054 ( \28397 , \28395 , \28396 );
and \U$28055 ( \28398 , \8486 , RI9870510_87);
and \U$28056 ( \28399 , RI9870330_83, \8484 );
nor \U$28057 ( \28400 , \28398 , \28399 );
and \U$28058 ( \28401 , \28400 , \8050 );
not \U$28059 ( \28402 , \28400 );
and \U$28060 ( \28403 , \28402 , \8051 );
nor \U$28061 ( \28404 , \28401 , \28403 );
nand \U$28062 ( \28405 , RI9870420_85, \7727 );
and \U$28063 ( \28406 , \28405 , \7480 );
not \U$28064 ( \28407 , \28405 );
and \U$28065 ( \28408 , \28407 , \7733 );
nor \U$28066 ( \28409 , \28406 , \28408 );
xor \U$28067 ( \28410 , \28404 , \28409 );
and \U$28068 ( \28411 , \9237 , RI9870240_81);
and \U$28069 ( \28412 , RI98706f0_91, \9235 );
nor \U$28070 ( \28413 , \28411 , \28412 );
and \U$28071 ( \28414 , \28413 , \9241 );
not \U$28072 ( \28415 , \28413 );
and \U$28073 ( \28416 , \28415 , \8836 );
nor \U$28074 ( \28417 , \28414 , \28416 );
xor \U$28075 ( \28418 , \28410 , \28417 );
and \U$28076 ( \28419 , \13045 , RI986fe80_73);
and \U$28077 ( \28420 , RI9870060_77, \13043 );
nor \U$28078 ( \28421 , \28419 , \28420 );
and \U$28079 ( \28422 , \28421 , \13047 );
not \U$28080 ( \28423 , \28421 );
and \U$28081 ( \28424 , \28423 , \12619 );
nor \U$28082 ( \28425 , \28422 , \28424 );
and \U$28083 ( \28426 , \12293 , RI986fca0_69);
and \U$28084 ( \28427 , RI986ff70_75, \12291 );
nor \U$28085 ( \28428 , \28426 , \28427 );
and \U$28086 ( \28429 , \28428 , \11687 );
not \U$28087 ( \28430 , \28428 );
and \U$28088 ( \28431 , \28430 , \11686 );
nor \U$28089 ( \28432 , \28429 , \28431 );
xor \U$28090 ( \28433 , \28425 , \28432 );
and \U$28091 ( \28434 , \13882 , RI9870150_79);
and \U$28092 ( \28435 , RI9870f60_109, \13880 );
nor \U$28093 ( \28436 , \28434 , \28435 );
and \U$28094 ( \28437 , \28436 , \13358 );
not \U$28095 ( \28438 , \28436 );
and \U$28096 ( \28439 , \28438 , \13359 );
nor \U$28097 ( \28440 , \28437 , \28439 );
xor \U$28098 ( \28441 , \28433 , \28440 );
and \U$28099 ( \28442 , \28418 , \28441 );
and \U$28100 ( \28443 , \9505 , RI9870600_89);
and \U$28101 ( \28444 , RI98708d0_95, \9503 );
nor \U$28102 ( \28445 , \28443 , \28444 );
and \U$28103 ( \28446 , \28445 , \9510 );
not \U$28104 ( \28447 , \28445 );
and \U$28105 ( \28448 , \28447 , \9513 );
nor \U$28106 ( \28449 , \28446 , \28448 );
and \U$28107 ( \28450 , \10424 , RI98707e0_93);
and \U$28108 ( \28451 , RI986fac0_65, \10422 );
nor \U$28109 ( \28452 , \28450 , \28451 );
and \U$28110 ( \28453 , \28452 , \9840 );
not \U$28111 ( \28454 , \28452 );
and \U$28112 ( \28455 , \28454 , \10428 );
nor \U$28113 ( \28456 , \28453 , \28455 );
xor \U$28114 ( \28457 , \28449 , \28456 );
and \U$28115 ( \28458 , \11696 , RI986fbb0_67);
and \U$28116 ( \28459 , RI986fd90_71, \11694 );
nor \U$28117 ( \28460 , \28458 , \28459 );
and \U$28118 ( \28461 , \28460 , \10965 );
not \U$28119 ( \28462 , \28460 );
and \U$28120 ( \28463 , \28462 , \11702 );
nor \U$28121 ( \28464 , \28461 , \28463 );
xor \U$28122 ( \28465 , \28457 , \28464 );
xor \U$28123 ( \28466 , \28425 , \28432 );
xor \U$28124 ( \28467 , \28466 , \28440 );
and \U$28125 ( \28468 , \28465 , \28467 );
and \U$28126 ( \28469 , \28418 , \28465 );
or \U$28127 ( \28470 , \28442 , \28468 , \28469 );
not \U$28128 ( \28471 , \28470 );
xor \U$28129 ( \28472 , \28397 , \28471 );
and \U$28130 ( \28473 , \15780 , RI9870e70_107);
and \U$28131 ( \28474 , RI9873648_192, RI9870ba0_101);
nor \U$28132 ( \28475 , \28473 , \28474 );
not \U$28133 ( \28476 , \28475 );
not \U$28134 ( \28477 , RI9873558_190);
and \U$28135 ( \28478 , \28476 , \28477 );
and \U$28136 ( \28479 , \28475 , RI9873558_190);
nor \U$28137 ( \28480 , \28478 , \28479 );
and \U$28138 ( \28481 , \14937 , RI9870d80_105);
and \U$28139 ( \28482 , RI98709c0_97, \14935 );
nor \U$28140 ( \28483 , \28481 , \28482 );
and \U$28141 ( \28484 , \28483 , \14538 );
not \U$28142 ( \28485 , \28483 );
and \U$28143 ( \28486 , \28485 , \14539 );
nor \U$28144 ( \28487 , \28484 , \28486 );
xor \U$28145 ( \28488 , \28480 , \28487 );
and \U$28146 ( \28489 , \13882 , RI9870f60_109);
and \U$28147 ( \28490 , RI9870ab0_99, \13880 );
nor \U$28148 ( \28491 , \28489 , \28490 );
and \U$28149 ( \28492 , \28491 , \13359 );
not \U$28150 ( \28493 , \28491 );
and \U$28151 ( \28494 , \28493 , \13358 );
nor \U$28152 ( \28495 , \28492 , \28494 );
xor \U$28153 ( \28496 , \28488 , \28495 );
and \U$28154 ( \28497 , \9505 , RI98708d0_95);
and \U$28155 ( \28498 , RI98707e0_93, \9503 );
nor \U$28156 ( \28499 , \28497 , \28498 );
and \U$28157 ( \28500 , \28499 , \9513 );
not \U$28158 ( \28501 , \28499 );
and \U$28159 ( \28502 , \28501 , \9510 );
nor \U$28160 ( \28503 , \28500 , \28502 );
and \U$28161 ( \28504 , \10424 , RI986fac0_65);
and \U$28162 ( \28505 , RI986fbb0_67, \10422 );
nor \U$28163 ( \28506 , \28504 , \28505 );
and \U$28164 ( \28507 , \28506 , \10428 );
not \U$28165 ( \28508 , \28506 );
and \U$28166 ( \28509 , \28508 , \9840 );
nor \U$28167 ( \28510 , \28507 , \28509 );
xor \U$28168 ( \28511 , \28503 , \28510 );
and \U$28169 ( \28512 , \9237 , RI98706f0_91);
and \U$28170 ( \28513 , RI9870600_89, \9235 );
nor \U$28171 ( \28514 , \28512 , \28513 );
and \U$28172 ( \28515 , \28514 , \8836 );
not \U$28173 ( \28516 , \28514 );
and \U$28174 ( \28517 , \28516 , \9241 );
nor \U$28175 ( \28518 , \28515 , \28517 );
xor \U$28176 ( \28519 , \28511 , \28518 );
xor \U$28177 ( \28520 , \28496 , \28519 );
and \U$28178 ( \28521 , \12293 , RI986ff70_75);
and \U$28179 ( \28522 , RI986fe80_73, \12291 );
nor \U$28180 ( \28523 , \28521 , \28522 );
and \U$28181 ( \28524 , \28523 , \11686 );
not \U$28182 ( \28525 , \28523 );
and \U$28183 ( \28526 , \28525 , \11687 );
nor \U$28184 ( \28527 , \28524 , \28526 );
and \U$28185 ( \28528 , \13045 , RI9870060_77);
and \U$28186 ( \28529 , RI9870150_79, \13043 );
nor \U$28187 ( \28530 , \28528 , \28529 );
and \U$28188 ( \28531 , \28530 , \12619 );
not \U$28189 ( \28532 , \28530 );
and \U$28190 ( \28533 , \28532 , \13047 );
nor \U$28191 ( \28534 , \28531 , \28533 );
xor \U$28192 ( \28535 , \28527 , \28534 );
and \U$28193 ( \28536 , \11696 , RI986fd90_71);
and \U$28194 ( \28537 , RI986fca0_69, \11694 );
nor \U$28195 ( \28538 , \28536 , \28537 );
and \U$28196 ( \28539 , \28538 , \11702 );
not \U$28197 ( \28540 , \28538 );
and \U$28198 ( \28541 , \28540 , \10965 );
nor \U$28199 ( \28542 , \28539 , \28541 );
xor \U$28200 ( \28543 , \28535 , \28542 );
xor \U$28201 ( \28544 , \28520 , \28543 );
and \U$28202 ( \28545 , \28472 , \28544 );
and \U$28203 ( \28546 , \28397 , \28471 );
nor \U$28204 ( \28547 , \28545 , \28546 );
xor \U$28205 ( \28548 , \28449 , \28456 );
and \U$28206 ( \28549 , \28548 , \28464 );
and \U$28207 ( \28550 , \28449 , \28456 );
or \U$28208 ( \28551 , \28549 , \28550 );
not \U$28209 ( \28552 , RI9873558_190);
and \U$28210 ( \28553 , \15780 , RI98709c0_97);
and \U$28211 ( \28554 , RI9873648_192, RI9870e70_107);
nor \U$28212 ( \28555 , \28553 , \28554 );
not \U$28213 ( \28556 , \28555 );
or \U$28214 ( \28557 , \28552 , \28556 );
or \U$28215 ( \28558 , \28555 , RI9873558_190);
nand \U$28216 ( \28559 , \28557 , \28558 );
xor \U$28217 ( \28560 , \28559 , \7733 );
and \U$28218 ( \28561 , \14937 , RI9870ab0_99);
and \U$28219 ( \28562 , RI9870d80_105, \14935 );
nor \U$28220 ( \28563 , \28561 , \28562 );
and \U$28221 ( \28564 , \28563 , \14539 );
not \U$28222 ( \28565 , \28563 );
and \U$28223 ( \28566 , \28565 , \14538 );
nor \U$28224 ( \28567 , \28564 , \28566 );
and \U$28225 ( \28568 , \28560 , \28567 );
and \U$28226 ( \28569 , \28559 , \7733 );
or \U$28227 ( \28570 , \28568 , \28569 );
xor \U$28228 ( \28571 , \28551 , \28570 );
xor \U$28229 ( \28572 , \28425 , \28432 );
and \U$28230 ( \28573 , \28572 , \28440 );
and \U$28231 ( \28574 , \28425 , \28432 );
or \U$28232 ( \28575 , \28573 , \28574 );
and \U$28233 ( \28576 , \28571 , \28575 );
and \U$28234 ( \28577 , \28551 , \28570 );
or \U$28235 ( \28578 , \28576 , \28577 );
and \U$28236 ( \28579 , \7729 , RI9870420_85);
and \U$28237 ( \28580 , RI9870510_87, \7727 );
nor \U$28238 ( \28581 , \28579 , \28580 );
and \U$28239 ( \28582 , \28581 , \7733 );
not \U$28240 ( \28583 , \28581 );
and \U$28241 ( \28584 , \28583 , \7480 );
nor \U$28242 ( \28585 , \28582 , \28584 );
and \U$28243 ( \28586 , \8486 , RI9870330_83);
and \U$28244 ( \28587 , RI9870240_81, \8484 );
nor \U$28245 ( \28588 , \28586 , \28587 );
and \U$28246 ( \28589 , \28588 , \8051 );
not \U$28247 ( \28590 , \28588 );
and \U$28248 ( \28591 , \28590 , \8050 );
nor \U$28249 ( \28592 , \28589 , \28591 );
or \U$28250 ( \28593 , \28585 , \28592 );
not \U$28251 ( \28594 , \28592 );
not \U$28252 ( \28595 , \28585 );
or \U$28253 ( \28596 , \28594 , \28595 );
xor \U$28254 ( \28597 , \28404 , \28409 );
and \U$28255 ( \28598 , \28597 , \28417 );
and \U$28256 ( \28599 , \28404 , \28409 );
or \U$28257 ( \28600 , \28598 , \28599 );
nand \U$28258 ( \28601 , \28596 , \28600 );
nand \U$28259 ( \28602 , \28593 , \28601 );
xor \U$28260 ( \28603 , \28578 , \28602 );
xor \U$28261 ( \28604 , \28496 , \28519 );
and \U$28262 ( \28605 , \28604 , \28543 );
and \U$28263 ( \28606 , \28496 , \28519 );
nor \U$28264 ( \28607 , \28605 , \28606 );
xor \U$28265 ( \28608 , \28603 , \28607 );
and \U$28266 ( \28609 , \28547 , \28608 );
xor \U$28267 ( \28610 , \28503 , \28510 );
and \U$28268 ( \28611 , \28610 , \28518 );
and \U$28269 ( \28612 , \28503 , \28510 );
nor \U$28270 ( \28613 , \28611 , \28612 );
xor \U$28271 ( \28614 , \28480 , \28487 );
and \U$28272 ( \28615 , \28614 , \28495 );
and \U$28273 ( \28616 , \28480 , \28487 );
nor \U$28274 ( \28617 , \28615 , \28616 );
xor \U$28275 ( \28618 , \28613 , \28617 );
xor \U$28276 ( \28619 , \28527 , \28534 );
and \U$28277 ( \28620 , \28619 , \28542 );
and \U$28278 ( \28621 , \28527 , \28534 );
nor \U$28279 ( \28622 , \28620 , \28621 );
xor \U$28280 ( \28623 , \28618 , \28622 );
xor \U$28281 ( \28624 , \28200 , \28207 );
xor \U$28282 ( \28625 , \28624 , \28215 );
not \U$28283 ( \28626 , \28625 );
xor \U$28284 ( \28627 , \28181 , \6709 );
xor \U$28285 ( \28628 , \28627 , \28189 );
not \U$28286 ( \28629 , \28628 );
or \U$28287 ( \28630 , \28626 , \28629 );
or \U$28288 ( \28631 , \28628 , \28625 );
nand \U$28289 ( \28632 , \28630 , \28631 );
xor \U$28290 ( \28633 , \28155 , \28162 );
xor \U$28291 ( \28634 , \28633 , \28170 );
nand \U$28292 ( \28635 , RI9870420_85, \7077 );
and \U$28293 ( \28636 , \28635 , \6710 );
not \U$28294 ( \28637 , \28635 );
and \U$28295 ( \28638 , \28637 , \6709 );
nor \U$28296 ( \28639 , \28636 , \28638 );
xor \U$28297 ( \28640 , \28234 , \28241 );
xor \U$28298 ( \28641 , \28640 , \28249 );
xor \U$28299 ( \28642 , \28639 , \28641 );
xor \U$28300 ( \28643 , \28634 , \28642 );
xor \U$28301 ( \28644 , \28632 , \28643 );
xor \U$28302 ( \28645 , \28623 , \28644 );
xor \U$28303 ( \28646 , \28578 , \28602 );
xor \U$28304 ( \28647 , \28646 , \28607 );
and \U$28305 ( \28648 , \28645 , \28647 );
and \U$28306 ( \28649 , \28547 , \28645 );
or \U$28307 ( \28650 , \28609 , \28648 , \28649 );
not \U$28308 ( \28651 , \28650 );
xor \U$28309 ( \28652 , \28613 , \28617 );
and \U$28310 ( \28653 , \28652 , \28622 );
and \U$28311 ( \28654 , \28613 , \28617 );
or \U$28312 ( \28655 , \28653 , \28654 );
not \U$28313 ( \28656 , \28655 );
xor \U$28314 ( \28657 , \28155 , \28162 );
xor \U$28315 ( \28658 , \28657 , \28170 );
and \U$28316 ( \28659 , \28639 , \28658 );
xor \U$28317 ( \28660 , \28155 , \28162 );
xor \U$28318 ( \28661 , \28660 , \28170 );
and \U$28319 ( \28662 , \28641 , \28661 );
and \U$28320 ( \28663 , \28639 , \28641 );
or \U$28321 ( \28664 , \28659 , \28662 , \28663 );
not \U$28322 ( \28665 , \28664 );
not \U$28323 ( \28666 , \28665 );
or \U$28324 ( \28667 , \28656 , \28666 );
or \U$28325 ( \28668 , \28665 , \28655 );
nand \U$28326 ( \28669 , \28667 , \28668 );
not \U$28327 ( \28670 , \28669 );
not \U$28328 ( \28671 , \28625 );
nand \U$28329 ( \28672 , \28671 , \28628 );
not \U$28330 ( \28673 , \28672 );
and \U$28331 ( \28674 , \28670 , \28673 );
and \U$28332 ( \28675 , \28669 , \28672 );
nor \U$28333 ( \28676 , \28674 , \28675 );
not \U$28334 ( \28677 , \28676 );
and \U$28335 ( \28678 , \28651 , \28677 );
and \U$28336 ( \28679 , \28650 , \28676 );
nor \U$28337 ( \28680 , \28678 , \28679 );
not \U$28338 ( \28681 , \28680 );
xor \U$28339 ( \28682 , \28613 , \28617 );
xor \U$28340 ( \28683 , \28682 , \28622 );
and \U$28341 ( \28684 , \28632 , \28683 );
xor \U$28342 ( \28685 , \28613 , \28617 );
xor \U$28343 ( \28686 , \28685 , \28622 );
and \U$28344 ( \28687 , \28643 , \28686 );
and \U$28345 ( \28688 , \28632 , \28643 );
or \U$28346 ( \28689 , \28684 , \28687 , \28688 );
xor \U$28347 ( \28690 , \28578 , \28602 );
and \U$28348 ( \28691 , \28690 , \28607 );
and \U$28349 ( \28692 , \28578 , \28602 );
or \U$28350 ( \28693 , \28691 , \28692 );
xor \U$28351 ( \28694 , \28689 , \28693 );
xor \U$28352 ( \28695 , \28173 , \28192 );
xor \U$28353 ( \28696 , \28695 , \28218 );
xor \U$28354 ( \28697 , \28223 , \28225 );
xor \U$28355 ( \28698 , \28010 , \28017 );
xor \U$28356 ( \28699 , \28698 , \28025 );
xor \U$28357 ( \28700 , \28252 , \28257 );
xor \U$28358 ( \28701 , \28699 , \28700 );
xor \U$28359 ( \28702 , \28697 , \28701 );
xor \U$28360 ( \28703 , \28696 , \28702 );
xor \U$28361 ( \28704 , \28694 , \28703 );
not \U$28362 ( \28705 , \28704 );
and \U$28363 ( \28706 , \28681 , \28705 );
and \U$28364 ( \28707 , \28680 , \28704 );
nor \U$28365 ( \28708 , \28706 , \28707 );
xor \U$28366 ( \28709 , \28578 , \28602 );
xor \U$28367 ( \28710 , \28709 , \28607 );
xor \U$28368 ( \28711 , \28547 , \28645 );
xor \U$28369 ( \28712 , \28710 , \28711 );
xor \U$28370 ( \28713 , \28551 , \28570 );
xor \U$28371 ( \28714 , \28713 , \28575 );
not \U$28372 ( \28715 , \28714 );
xor \U$28373 ( \28716 , \28397 , \28471 );
xor \U$28374 ( \28717 , \28716 , \28544 );
nor \U$28375 ( \28718 , \28715 , \28717 );
xor \U$28376 ( \28719 , \28712 , \28718 );
xor \U$28377 ( \28720 , \28559 , \7733 );
xor \U$28378 ( \28721 , \28720 , \28567 );
and \U$28379 ( \28722 , \12293 , RI986fbb0_67);
and \U$28380 ( \28723 , RI986fd90_71, \12291 );
nor \U$28381 ( \28724 , \28722 , \28723 );
and \U$28382 ( \28725 , \28724 , \11687 );
not \U$28383 ( \28726 , \28724 );
and \U$28384 ( \28727 , \28726 , \11686 );
nor \U$28385 ( \28728 , \28725 , \28727 );
and \U$28386 ( \28729 , \13045 , RI986fca0_69);
and \U$28387 ( \28730 , RI986ff70_75, \13043 );
nor \U$28388 ( \28731 , \28729 , \28730 );
and \U$28389 ( \28732 , \28731 , \13047 );
not \U$28390 ( \28733 , \28731 );
and \U$28391 ( \28734 , \28733 , \12619 );
nor \U$28392 ( \28735 , \28732 , \28734 );
xor \U$28393 ( \28736 , \28728 , \28735 );
and \U$28394 ( \28737 , \13882 , RI986fe80_73);
and \U$28395 ( \28738 , RI9870060_77, \13880 );
nor \U$28396 ( \28739 , \28737 , \28738 );
and \U$28397 ( \28740 , \28739 , \13358 );
not \U$28398 ( \28741 , \28739 );
and \U$28399 ( \28742 , \28741 , \13359 );
nor \U$28400 ( \28743 , \28740 , \28742 );
and \U$28401 ( \28744 , \28736 , \28743 );
and \U$28402 ( \28745 , \28728 , \28735 );
or \U$28403 ( \28746 , \28744 , \28745 );
not \U$28404 ( \28747 , RI9873558_190);
and \U$28405 ( \28748 , \15780 , RI9870ab0_99);
and \U$28406 ( \28749 , RI9873648_192, RI9870d80_105);
nor \U$28407 ( \28750 , \28748 , \28749 );
not \U$28408 ( \28751 , \28750 );
or \U$28409 ( \28752 , \28747 , \28751 );
or \U$28410 ( \28753 , \28750 , RI9873558_190);
nand \U$28411 ( \28754 , \28752 , \28753 );
xor \U$28412 ( \28755 , \28754 , \8051 );
and \U$28413 ( \28756 , \14937 , RI9870150_79);
and \U$28414 ( \28757 , RI9870f60_109, \14935 );
nor \U$28415 ( \28758 , \28756 , \28757 );
and \U$28416 ( \28759 , \28758 , \14539 );
not \U$28417 ( \28760 , \28758 );
and \U$28418 ( \28761 , \28760 , \14538 );
nor \U$28419 ( \28762 , \28759 , \28761 );
and \U$28420 ( \28763 , \28755 , \28762 );
and \U$28421 ( \28764 , \28754 , \8051 );
or \U$28422 ( \28765 , \28763 , \28764 );
xor \U$28423 ( \28766 , \28746 , \28765 );
and \U$28424 ( \28767 , \9505 , RI9870240_81);
and \U$28425 ( \28768 , RI98706f0_91, \9503 );
nor \U$28426 ( \28769 , \28767 , \28768 );
and \U$28427 ( \28770 , \28769 , \9510 );
not \U$28428 ( \28771 , \28769 );
and \U$28429 ( \28772 , \28771 , \9513 );
nor \U$28430 ( \28773 , \28770 , \28772 );
and \U$28431 ( \28774 , \10424 , RI9870600_89);
and \U$28432 ( \28775 , RI98708d0_95, \10422 );
nor \U$28433 ( \28776 , \28774 , \28775 );
and \U$28434 ( \28777 , \28776 , \9840 );
not \U$28435 ( \28778 , \28776 );
and \U$28436 ( \28779 , \28778 , \10428 );
nor \U$28437 ( \28780 , \28777 , \28779 );
xor \U$28438 ( \28781 , \28773 , \28780 );
and \U$28439 ( \28782 , \11696 , RI98707e0_93);
and \U$28440 ( \28783 , RI986fac0_65, \11694 );
nor \U$28441 ( \28784 , \28782 , \28783 );
and \U$28442 ( \28785 , \28784 , \10965 );
not \U$28443 ( \28786 , \28784 );
and \U$28444 ( \28787 , \28786 , \11702 );
nor \U$28445 ( \28788 , \28785 , \28787 );
and \U$28446 ( \28789 , \28781 , \28788 );
and \U$28447 ( \28790 , \28773 , \28780 );
or \U$28448 ( \28791 , \28789 , \28790 );
and \U$28449 ( \28792 , \28766 , \28791 );
and \U$28450 ( \28793 , \28746 , \28765 );
or \U$28451 ( \28794 , \28792 , \28793 );
xor \U$28452 ( \28795 , \28721 , \28794 );
and \U$28453 ( \28796 , \8486 , RI9870420_85);
and \U$28454 ( \28797 , RI9870510_87, \8484 );
nor \U$28455 ( \28798 , \28796 , \28797 );
and \U$28456 ( \28799 , \28798 , \8050 );
not \U$28457 ( \28800 , \28798 );
and \U$28458 ( \28801 , \28800 , \8051 );
nor \U$28459 ( \28802 , \28799 , \28801 );
xor \U$28460 ( \28803 , \28324 , \28331 );
xor \U$28461 ( \28804 , \28803 , \28339 );
and \U$28462 ( \28805 , \28802 , \28804 );
xor \U$28463 ( \28806 , \28376 , \28383 );
xor \U$28464 ( \28807 , \28806 , \28391 );
xor \U$28465 ( \28808 , \28324 , \28331 );
xor \U$28466 ( \28809 , \28808 , \28339 );
and \U$28467 ( \28810 , \28807 , \28809 );
and \U$28468 ( \28811 , \28802 , \28807 );
or \U$28469 ( \28812 , \28805 , \28810 , \28811 );
and \U$28470 ( \28813 , \28795 , \28812 );
and \U$28471 ( \28814 , \28721 , \28794 );
nor \U$28472 ( \28815 , \28813 , \28814 );
not \U$28473 ( \28816 , \28592 );
not \U$28474 ( \28817 , \28600 );
or \U$28475 ( \28818 , \28816 , \28817 );
or \U$28476 ( \28819 , \28600 , \28592 );
nand \U$28477 ( \28820 , \28818 , \28819 );
not \U$28478 ( \28821 , \28820 );
not \U$28479 ( \28822 , \28585 );
and \U$28480 ( \28823 , \28821 , \28822 );
and \U$28481 ( \28824 , \28820 , \28585 );
nor \U$28482 ( \28825 , \28823 , \28824 );
or \U$28483 ( \28826 , \28815 , \28825 );
not \U$28484 ( \28827 , \28825 );
not \U$28485 ( \28828 , \28815 );
or \U$28486 ( \28829 , \28827 , \28828 );
xor \U$28487 ( \28830 , \28342 , \28368 );
xor \U$28488 ( \28831 , \28830 , \28394 );
xor \U$28489 ( \28832 , \28425 , \28432 );
xor \U$28490 ( \28833 , \28832 , \28440 );
xor \U$28491 ( \28834 , \28418 , \28465 );
xor \U$28492 ( \28835 , \28833 , \28834 );
and \U$28493 ( \28836 , \28831 , \28835 );
nand \U$28494 ( \28837 , \28829 , \28836 );
nand \U$28495 ( \28838 , \28826 , \28837 );
and \U$28496 ( \28839 , \28719 , \28838 );
and \U$28497 ( \28840 , \28712 , \28718 );
nor \U$28498 ( \28841 , \28839 , \28840 );
or \U$28499 ( \28842 , \28708 , \28841 );
xnor \U$28500 ( \28843 , \28841 , \28708 );
not \U$28501 ( \28844 , RI9873558_190);
and \U$28502 ( \28845 , \15780 , RI986fe80_73);
and \U$28503 ( \28846 , RI9873648_192, RI9870060_77);
nor \U$28504 ( \28847 , \28845 , \28846 );
not \U$28505 ( \28848 , \28847 );
or \U$28506 ( \28849 , \28844 , \28848 );
or \U$28507 ( \28850 , \28847 , RI9873558_190);
nand \U$28508 ( \28851 , \28849 , \28850 );
and \U$28509 ( \28852 , \28851 , \9513 );
not \U$28510 ( \28853 , \28851 );
not \U$28511 ( \28854 , \9513 );
and \U$28512 ( \28855 , \28853 , \28854 );
and \U$28513 ( \28856 , \14937 , RI986fca0_69);
and \U$28514 ( \28857 , RI986ff70_75, \14935 );
nor \U$28515 ( \28858 , \28856 , \28857 );
and \U$28516 ( \28859 , \28858 , \14538 );
not \U$28517 ( \28860 , \28858 );
and \U$28518 ( \28861 , \28860 , \14539 );
nor \U$28519 ( \28862 , \28859 , \28861 );
nor \U$28520 ( \28863 , \28855 , \28862 );
nor \U$28521 ( \28864 , \28852 , \28863 );
and \U$28522 ( \28865 , \11696 , RI9870240_81);
and \U$28523 ( \28866 , RI98706f0_91, \11694 );
nor \U$28524 ( \28867 , \28865 , \28866 );
and \U$28525 ( \28868 , \28867 , \11702 );
not \U$28526 ( \28869 , \28867 );
and \U$28527 ( \28870 , \28869 , \10965 );
nor \U$28528 ( \28871 , \28868 , \28870 );
not \U$28529 ( \28872 , \28871 );
nand \U$28530 ( \28873 , RI9870420_85, \9503 );
and \U$28531 ( \28874 , \28873 , \9513 );
not \U$28532 ( \28875 , \28873 );
and \U$28533 ( \28876 , \28875 , \9510 );
nor \U$28534 ( \28877 , \28874 , \28876 );
not \U$28535 ( \28878 , \28877 );
and \U$28536 ( \28879 , \28872 , \28878 );
and \U$28537 ( \28880 , \28871 , \28877 );
and \U$28538 ( \28881 , \10424 , RI9870510_87);
and \U$28539 ( \28882 , RI9870330_83, \10422 );
nor \U$28540 ( \28883 , \28881 , \28882 );
and \U$28541 ( \28884 , \28883 , \10428 );
not \U$28542 ( \28885 , \28883 );
and \U$28543 ( \28886 , \28885 , \9840 );
nor \U$28544 ( \28887 , \28884 , \28886 );
nor \U$28545 ( \28888 , \28880 , \28887 );
nor \U$28546 ( \28889 , \28879 , \28888 );
xor \U$28547 ( \28890 , \28864 , \28889 );
and \U$28548 ( \28891 , \12293 , RI9870600_89);
and \U$28549 ( \28892 , RI98708d0_95, \12291 );
nor \U$28550 ( \28893 , \28891 , \28892 );
and \U$28551 ( \28894 , \28893 , \11686 );
not \U$28552 ( \28895 , \28893 );
and \U$28553 ( \28896 , \28895 , \11687 );
nor \U$28554 ( \28897 , \28894 , \28896 );
and \U$28555 ( \28898 , \13045 , RI98707e0_93);
and \U$28556 ( \28899 , RI986fac0_65, \13043 );
nor \U$28557 ( \28900 , \28898 , \28899 );
and \U$28558 ( \28901 , \28900 , \12619 );
not \U$28559 ( \28902 , \28900 );
and \U$28560 ( \28903 , \28902 , \13047 );
nor \U$28561 ( \28904 , \28901 , \28903 );
xor \U$28562 ( \28905 , \28897 , \28904 );
and \U$28563 ( \28906 , \13882 , RI986fbb0_67);
and \U$28564 ( \28907 , RI986fd90_71, \13880 );
nor \U$28565 ( \28908 , \28906 , \28907 );
and \U$28566 ( \28909 , \28908 , \13359 );
not \U$28567 ( \28910 , \28908 );
and \U$28568 ( \28911 , \28910 , \13358 );
nor \U$28569 ( \28912 , \28909 , \28911 );
and \U$28570 ( \28913 , \28905 , \28912 );
and \U$28571 ( \28914 , \28897 , \28904 );
or \U$28572 ( \28915 , \28913 , \28914 );
and \U$28573 ( \28916 , \28890 , \28915 );
and \U$28574 ( \28917 , \28864 , \28889 );
nor \U$28575 ( \28918 , \28916 , \28917 );
not \U$28576 ( \28919 , RI9873558_190);
and \U$28577 ( \28920 , \15780 , RI9870150_79);
and \U$28578 ( \28921 , RI9873648_192, RI9870f60_109);
nor \U$28579 ( \28922 , \28920 , \28921 );
not \U$28580 ( \28923 , \28922 );
or \U$28581 ( \28924 , \28919 , \28923 );
or \U$28582 ( \28925 , \28922 , RI9873558_190);
nand \U$28583 ( \28926 , \28924 , \28925 );
xor \U$28584 ( \28927 , \28926 , \8836 );
and \U$28585 ( \28928 , \14937 , RI986fe80_73);
and \U$28586 ( \28929 , RI9870060_77, \14935 );
nor \U$28587 ( \28930 , \28928 , \28929 );
and \U$28588 ( \28931 , \28930 , \14539 );
not \U$28589 ( \28932 , \28930 );
and \U$28590 ( \28933 , \28932 , \14538 );
nor \U$28591 ( \28934 , \28931 , \28933 );
xor \U$28592 ( \28935 , \28927 , \28934 );
xor \U$28593 ( \28936 , \28918 , \28935 );
and \U$28594 ( \28937 , \9505 , RI9870420_85);
and \U$28595 ( \28938 , RI9870510_87, \9503 );
nor \U$28596 ( \28939 , \28937 , \28938 );
and \U$28597 ( \28940 , \28939 , \9513 );
not \U$28598 ( \28941 , \28939 );
and \U$28599 ( \28942 , \28941 , \9510 );
nor \U$28600 ( \28943 , \28940 , \28942 );
not \U$28601 ( \28944 , \28943 );
and \U$28602 ( \28945 , \10424 , RI9870330_83);
and \U$28603 ( \28946 , RI9870240_81, \10422 );
nor \U$28604 ( \28947 , \28945 , \28946 );
and \U$28605 ( \28948 , \28947 , \9840 );
not \U$28606 ( \28949 , \28947 );
and \U$28607 ( \28950 , \28949 , \10428 );
nor \U$28608 ( \28951 , \28948 , \28950 );
not \U$28609 ( \28952 , \28951 );
or \U$28610 ( \28953 , \28944 , \28952 );
or \U$28611 ( \28954 , \28943 , \28951 );
nand \U$28612 ( \28955 , \28953 , \28954 );
not \U$28613 ( \28956 , \28955 );
and \U$28614 ( \28957 , \12293 , RI98708d0_95);
and \U$28615 ( \28958 , RI98707e0_93, \12291 );
nor \U$28616 ( \28959 , \28957 , \28958 );
and \U$28617 ( \28960 , \28959 , \11687 );
not \U$28618 ( \28961 , \28959 );
and \U$28619 ( \28962 , \28961 , \11686 );
nor \U$28620 ( \28963 , \28960 , \28962 );
and \U$28621 ( \28964 , \13045 , RI986fac0_65);
and \U$28622 ( \28965 , RI986fbb0_67, \13043 );
nor \U$28623 ( \28966 , \28964 , \28965 );
and \U$28624 ( \28967 , \28966 , \13047 );
not \U$28625 ( \28968 , \28966 );
and \U$28626 ( \28969 , \28968 , \12619 );
nor \U$28627 ( \28970 , \28967 , \28969 );
xor \U$28628 ( \28971 , \28963 , \28970 );
and \U$28629 ( \28972 , \11696 , RI98706f0_91);
and \U$28630 ( \28973 , RI9870600_89, \11694 );
nor \U$28631 ( \28974 , \28972 , \28973 );
and \U$28632 ( \28975 , \28974 , \10965 );
not \U$28633 ( \28976 , \28974 );
and \U$28634 ( \28977 , \28976 , \11702 );
nor \U$28635 ( \28978 , \28975 , \28977 );
xor \U$28636 ( \28979 , \28971 , \28978 );
not \U$28637 ( \28980 , \28979 );
or \U$28638 ( \28981 , \28956 , \28980 );
or \U$28639 ( \28982 , \28979 , \28955 );
and \U$28640 ( \28983 , \14937 , RI986ff70_75);
and \U$28641 ( \28984 , RI986fe80_73, \14935 );
nor \U$28642 ( \28985 , \28983 , \28984 );
and \U$28643 ( \28986 , \28985 , \14539 );
not \U$28644 ( \28987 , \28985 );
and \U$28645 ( \28988 , \28987 , \14538 );
nor \U$28646 ( \28989 , \28986 , \28988 );
not \U$28647 ( \28990 , RI9873558_190);
and \U$28648 ( \28991 , \15780 , RI9870060_77);
and \U$28649 ( \28992 , RI9873648_192, RI9870150_79);
nor \U$28650 ( \28993 , \28991 , \28992 );
not \U$28651 ( \28994 , \28993 );
or \U$28652 ( \28995 , \28990 , \28994 );
or \U$28653 ( \28996 , \28993 , RI9873558_190);
nand \U$28654 ( \28997 , \28995 , \28996 );
xor \U$28655 ( \28998 , \28989 , \28997 );
and \U$28656 ( \28999 , \13882 , RI986fd90_71);
and \U$28657 ( \29000 , RI986fca0_69, \13880 );
nor \U$28658 ( \29001 , \28999 , \29000 );
and \U$28659 ( \29002 , \29001 , \13358 );
not \U$28660 ( \29003 , \29001 );
and \U$28661 ( \29004 , \29003 , \13359 );
nor \U$28662 ( \29005 , \29002 , \29004 );
xor \U$28663 ( \29006 , \28998 , \29005 );
nand \U$28664 ( \29007 , \28982 , \29006 );
nand \U$28665 ( \29008 , \28981 , \29007 );
and \U$28666 ( \29009 , \28936 , \29008 );
and \U$28667 ( \29010 , \28918 , \28935 );
or \U$28668 ( \29011 , \29009 , \29010 );
and \U$28669 ( \29012 , \13045 , RI986fbb0_67);
and \U$28670 ( \29013 , RI986fd90_71, \13043 );
nor \U$28671 ( \29014 , \29012 , \29013 );
and \U$28672 ( \29015 , \29014 , \13047 );
not \U$28673 ( \29016 , \29014 );
and \U$28674 ( \29017 , \29016 , \12619 );
nor \U$28675 ( \29018 , \29015 , \29017 );
and \U$28676 ( \29019 , \12293 , RI98707e0_93);
and \U$28677 ( \29020 , RI986fac0_65, \12291 );
nor \U$28678 ( \29021 , \29019 , \29020 );
and \U$28679 ( \29022 , \29021 , \11687 );
not \U$28680 ( \29023 , \29021 );
and \U$28681 ( \29024 , \29023 , \11686 );
nor \U$28682 ( \29025 , \29022 , \29024 );
xor \U$28683 ( \29026 , \29018 , \29025 );
and \U$28684 ( \29027 , \13882 , RI986fca0_69);
and \U$28685 ( \29028 , RI986ff70_75, \13880 );
nor \U$28686 ( \29029 , \29027 , \29028 );
and \U$28687 ( \29030 , \29029 , \13358 );
not \U$28688 ( \29031 , \29029 );
and \U$28689 ( \29032 , \29031 , \13359 );
nor \U$28690 ( \29033 , \29030 , \29032 );
and \U$28691 ( \29034 , \29026 , \29033 );
and \U$28692 ( \29035 , \29018 , \29025 );
or \U$28693 ( \29036 , \29034 , \29035 );
xor \U$28694 ( \29037 , \28926 , \8836 );
and \U$28695 ( \29038 , \29037 , \28934 );
and \U$28696 ( \29039 , \28926 , \8836 );
or \U$28697 ( \29040 , \29038 , \29039 );
xor \U$28698 ( \29041 , \29036 , \29040 );
and \U$28699 ( \29042 , \9505 , RI9870510_87);
and \U$28700 ( \29043 , RI9870330_83, \9503 );
nor \U$28701 ( \29044 , \29042 , \29043 );
and \U$28702 ( \29045 , \29044 , \9510 );
not \U$28703 ( \29046 , \29044 );
and \U$28704 ( \29047 , \29046 , \9513 );
nor \U$28705 ( \29048 , \29045 , \29047 );
and \U$28706 ( \29049 , \10424 , RI9870240_81);
and \U$28707 ( \29050 , RI98706f0_91, \10422 );
nor \U$28708 ( \29051 , \29049 , \29050 );
and \U$28709 ( \29052 , \29051 , \9840 );
not \U$28710 ( \29053 , \29051 );
and \U$28711 ( \29054 , \29053 , \10428 );
nor \U$28712 ( \29055 , \29052 , \29054 );
xor \U$28713 ( \29056 , \29048 , \29055 );
and \U$28714 ( \29057 , \11696 , RI9870600_89);
and \U$28715 ( \29058 , RI98708d0_95, \11694 );
nor \U$28716 ( \29059 , \29057 , \29058 );
and \U$28717 ( \29060 , \29059 , \10965 );
not \U$28718 ( \29061 , \29059 );
and \U$28719 ( \29062 , \29061 , \11702 );
nor \U$28720 ( \29063 , \29060 , \29062 );
and \U$28721 ( \29064 , \29056 , \29063 );
and \U$28722 ( \29065 , \29048 , \29055 );
or \U$28723 ( \29066 , \29064 , \29065 );
xor \U$28724 ( \29067 , \29041 , \29066 );
xor \U$28725 ( \29068 , \29011 , \29067 );
not \U$28726 ( \29069 , \28943 );
nand \U$28727 ( \29070 , \29069 , \28951 );
not \U$28728 ( \29071 , \29070 );
xor \U$28729 ( \29072 , \28989 , \28997 );
and \U$28730 ( \29073 , \29072 , \29005 );
and \U$28731 ( \29074 , \28989 , \28997 );
nor \U$28732 ( \29075 , \29073 , \29074 );
xor \U$28733 ( \29076 , \28963 , \28970 );
and \U$28734 ( \29077 , \29076 , \28978 );
and \U$28735 ( \29078 , \28963 , \28970 );
nor \U$28736 ( \29079 , \29077 , \29078 );
xor \U$28737 ( \29080 , \29075 , \29079 );
not \U$28738 ( \29081 , \29080 );
or \U$28739 ( \29082 , \29071 , \29081 );
or \U$28740 ( \29083 , \29080 , \29070 );
nand \U$28741 ( \29084 , \29082 , \29083 );
xor \U$28742 ( \29085 , \29048 , \29055 );
xor \U$28743 ( \29086 , \29085 , \29063 );
nand \U$28744 ( \29087 , RI9870420_85, \9235 );
and \U$28745 ( \29088 , \29087 , \9241 );
not \U$28746 ( \29089 , \29087 );
and \U$28747 ( \29090 , \29089 , \8836 );
nor \U$28748 ( \29091 , \29088 , \29090 );
xor \U$28749 ( \29092 , \29086 , \29091 );
xor \U$28750 ( \29093 , \29018 , \29025 );
xor \U$28751 ( \29094 , \29093 , \29033 );
xor \U$28752 ( \29095 , \29092 , \29094 );
and \U$28753 ( \29096 , \29084 , \29095 );
and \U$28754 ( \29097 , \29068 , \29096 );
and \U$28755 ( \29098 , \29011 , \29067 );
or \U$28756 ( \29099 , \29097 , \29098 );
not \U$28757 ( \29100 , \29099 );
not \U$28758 ( \29101 , \29075 );
not \U$28759 ( \29102 , \29070 );
and \U$28760 ( \29103 , \29101 , \29102 );
and \U$28761 ( \29104 , \29075 , \29070 );
nor \U$28762 ( \29105 , \29104 , \29079 );
nor \U$28763 ( \29106 , \29103 , \29105 );
xor \U$28764 ( \29107 , \29086 , \29091 );
and \U$28765 ( \29108 , \29107 , \29094 );
and \U$28766 ( \29109 , \29086 , \29091 );
nor \U$28767 ( \29110 , \29108 , \29109 );
xor \U$28768 ( \29111 , \29106 , \29110 );
and \U$28769 ( \29112 , \11696 , RI98708d0_95);
and \U$28770 ( \29113 , RI98707e0_93, \11694 );
nor \U$28771 ( \29114 , \29112 , \29113 );
and \U$28772 ( \29115 , \29114 , \10965 );
not \U$28773 ( \29116 , \29114 );
and \U$28774 ( \29117 , \29116 , \11702 );
nor \U$28775 ( \29118 , \29115 , \29117 );
and \U$28776 ( \29119 , \12293 , RI986fac0_65);
and \U$28777 ( \29120 , RI986fbb0_67, \12291 );
nor \U$28778 ( \29121 , \29119 , \29120 );
and \U$28779 ( \29122 , \29121 , \11687 );
not \U$28780 ( \29123 , \29121 );
and \U$28781 ( \29124 , \29123 , \11686 );
nor \U$28782 ( \29125 , \29122 , \29124 );
xor \U$28783 ( \29126 , \29118 , \29125 );
and \U$28784 ( \29127 , \13045 , RI986fd90_71);
and \U$28785 ( \29128 , RI986fca0_69, \13043 );
nor \U$28786 ( \29129 , \29127 , \29128 );
and \U$28787 ( \29130 , \29129 , \13047 );
not \U$28788 ( \29131 , \29129 );
and \U$28789 ( \29132 , \29131 , \12619 );
nor \U$28790 ( \29133 , \29130 , \29132 );
xor \U$28791 ( \29134 , \29126 , \29133 );
not \U$28792 ( \29135 , \29134 );
and \U$28793 ( \29136 , \15780 , RI9870f60_109);
and \U$28794 ( \29137 , RI9873648_192, RI9870ab0_99);
nor \U$28795 ( \29138 , \29136 , \29137 );
not \U$28796 ( \29139 , \29138 );
not \U$28797 ( \29140 , RI9873558_190);
and \U$28798 ( \29141 , \29139 , \29140 );
and \U$28799 ( \29142 , \29138 , RI9873558_190);
nor \U$28800 ( \29143 , \29141 , \29142 );
and \U$28801 ( \29144 , \14937 , RI9870060_77);
and \U$28802 ( \29145 , RI9870150_79, \14935 );
nor \U$28803 ( \29146 , \29144 , \29145 );
and \U$28804 ( \29147 , \29146 , \14538 );
not \U$28805 ( \29148 , \29146 );
and \U$28806 ( \29149 , \29148 , \14539 );
nor \U$28807 ( \29150 , \29147 , \29149 );
xor \U$28808 ( \29151 , \29143 , \29150 );
and \U$28809 ( \29152 , \13882 , RI986ff70_75);
and \U$28810 ( \29153 , RI986fe80_73, \13880 );
nor \U$28811 ( \29154 , \29152 , \29153 );
and \U$28812 ( \29155 , \29154 , \13359 );
not \U$28813 ( \29156 , \29154 );
and \U$28814 ( \29157 , \29156 , \13358 );
nor \U$28815 ( \29158 , \29155 , \29157 );
xor \U$28816 ( \29159 , \29151 , \29158 );
not \U$28817 ( \29160 , \29159 );
or \U$28818 ( \29161 , \29135 , \29160 );
or \U$28819 ( \29162 , \29159 , \29134 );
nand \U$28820 ( \29163 , \29161 , \29162 );
not \U$28821 ( \29164 , \29163 );
and \U$28822 ( \29165 , \9505 , RI9870330_83);
and \U$28823 ( \29166 , RI9870240_81, \9503 );
nor \U$28824 ( \29167 , \29165 , \29166 );
and \U$28825 ( \29168 , \29167 , \9513 );
not \U$28826 ( \29169 , \29167 );
and \U$28827 ( \29170 , \29169 , \9510 );
nor \U$28828 ( \29171 , \29168 , \29170 );
and \U$28829 ( \29172 , \10424 , RI98706f0_91);
and \U$28830 ( \29173 , RI9870600_89, \10422 );
nor \U$28831 ( \29174 , \29172 , \29173 );
and \U$28832 ( \29175 , \29174 , \10428 );
not \U$28833 ( \29176 , \29174 );
and \U$28834 ( \29177 , \29176 , \9840 );
nor \U$28835 ( \29178 , \29175 , \29177 );
xor \U$28836 ( \29179 , \29171 , \29178 );
and \U$28837 ( \29180 , \9237 , RI9870420_85);
and \U$28838 ( \29181 , RI9870510_87, \9235 );
nor \U$28839 ( \29182 , \29180 , \29181 );
and \U$28840 ( \29183 , \29182 , \8836 );
not \U$28841 ( \29184 , \29182 );
and \U$28842 ( \29185 , \29184 , \9241 );
nor \U$28843 ( \29186 , \29183 , \29185 );
xor \U$28844 ( \29187 , \29179 , \29186 );
not \U$28845 ( \29188 , \29187 );
and \U$28846 ( \29189 , \29164 , \29188 );
and \U$28847 ( \29190 , \29163 , \29187 );
nor \U$28848 ( \29191 , \29189 , \29190 );
and \U$28849 ( \29192 , \29111 , \29191 );
and \U$28850 ( \29193 , \29106 , \29110 );
nor \U$28851 ( \29194 , \29192 , \29193 );
xor \U$28852 ( \29195 , \29036 , \29040 );
and \U$28853 ( \29196 , \29195 , \29066 );
and \U$28854 ( \29197 , \29036 , \29040 );
or \U$28855 ( \29198 , \29196 , \29197 );
xor \U$28856 ( \29199 , \28728 , \28735 );
xor \U$28857 ( \29200 , \29199 , \28743 );
xor \U$28858 ( \29201 , \29198 , \29200 );
or \U$28859 ( \29202 , \29159 , \29187 );
not \U$28860 ( \29203 , \29187 );
not \U$28861 ( \29204 , \29159 );
or \U$28862 ( \29205 , \29203 , \29204 );
nand \U$28863 ( \29206 , \29205 , \29134 );
nand \U$28864 ( \29207 , \29202 , \29206 );
xor \U$28865 ( \29208 , \29201 , \29207 );
xnor \U$28866 ( \29209 , \29194 , \29208 );
not \U$28867 ( \29210 , \29209 );
and \U$28868 ( \29211 , \9237 , RI9870510_87);
and \U$28869 ( \29212 , RI9870330_83, \9235 );
nor \U$28870 ( \29213 , \29211 , \29212 );
and \U$28871 ( \29214 , \29213 , \9241 );
not \U$28872 ( \29215 , \29213 );
and \U$28873 ( \29216 , \29215 , \8836 );
nor \U$28874 ( \29217 , \29214 , \29216 );
nand \U$28875 ( \29218 , RI9870420_85, \8484 );
and \U$28876 ( \29219 , \29218 , \8050 );
not \U$28877 ( \29220 , \29218 );
and \U$28878 ( \29221 , \29220 , \8051 );
nor \U$28879 ( \29222 , \29219 , \29221 );
xor \U$28880 ( \29223 , \29217 , \29222 );
xor \U$28881 ( \29224 , \28773 , \28780 );
xor \U$28882 ( \29225 , \29224 , \28788 );
xor \U$28883 ( \29226 , \29223 , \29225 );
xor \U$28884 ( \29227 , \28754 , \8051 );
xor \U$28885 ( \29228 , \29227 , \28762 );
xor \U$28886 ( \29229 , \29118 , \29125 );
and \U$28887 ( \29230 , \29229 , \29133 );
and \U$28888 ( \29231 , \29118 , \29125 );
or \U$28889 ( \29232 , \29230 , \29231 );
xor \U$28890 ( \29233 , \29143 , \29150 );
and \U$28891 ( \29234 , \29233 , \29158 );
and \U$28892 ( \29235 , \29143 , \29150 );
nor \U$28893 ( \29236 , \29234 , \29235 );
xor \U$28894 ( \29237 , \29232 , \29236 );
xor \U$28895 ( \29238 , \29171 , \29178 );
and \U$28896 ( \29239 , \29238 , \29186 );
and \U$28897 ( \29240 , \29171 , \29178 );
nor \U$28898 ( \29241 , \29239 , \29240 );
xor \U$28899 ( \29242 , \29237 , \29241 );
xor \U$28900 ( \29243 , \29228 , \29242 );
xor \U$28901 ( \29244 , \29226 , \29243 );
not \U$28902 ( \29245 , \29244 );
and \U$28903 ( \29246 , \29210 , \29245 );
and \U$28904 ( \29247 , \29209 , \29244 );
nor \U$28905 ( \29248 , \29246 , \29247 );
not \U$28906 ( \29249 , \29248 );
or \U$28907 ( \29250 , \29100 , \29249 );
or \U$28908 ( \29251 , \29248 , \29099 );
nand \U$28909 ( \29252 , \29250 , \29251 );
xor \U$28910 ( \29253 , \29011 , \29067 );
xor \U$28911 ( \29254 , \29253 , \29096 );
not \U$28912 ( \29255 , \29254 );
xor \U$28913 ( \29256 , \29106 , \29110 );
xor \U$28914 ( \29257 , \29256 , \29191 );
nor \U$28915 ( \29258 , \29255 , \29257 );
and \U$28916 ( \29259 , \29252 , \29258 );
xor \U$28917 ( \29260 , \29258 , \29252 );
and \U$28918 ( \29261 , \13882 , RI986fac0_65);
and \U$28919 ( \29262 , RI986fbb0_67, \13880 );
nor \U$28920 ( \29263 , \29261 , \29262 );
and \U$28921 ( \29264 , \29263 , \13358 );
not \U$28922 ( \29265 , \29263 );
and \U$28923 ( \29266 , \29265 , \13359 );
nor \U$28924 ( \29267 , \29264 , \29266 );
not \U$28925 ( \29268 , RI9873558_190);
and \U$28926 ( \29269 , \15780 , RI986ff70_75);
and \U$28927 ( \29270 , RI9873648_192, RI986fe80_73);
nor \U$28928 ( \29271 , \29269 , \29270 );
not \U$28929 ( \29272 , \29271 );
or \U$28930 ( \29273 , \29268 , \29272 );
or \U$28931 ( \29274 , \29271 , RI9873558_190);
nand \U$28932 ( \29275 , \29273 , \29274 );
xor \U$28933 ( \29276 , \29267 , \29275 );
and \U$28934 ( \29277 , \14937 , RI986fd90_71);
and \U$28935 ( \29278 , RI986fca0_69, \14935 );
nor \U$28936 ( \29279 , \29277 , \29278 );
and \U$28937 ( \29280 , \29279 , \14539 );
not \U$28938 ( \29281 , \29279 );
and \U$28939 ( \29282 , \29281 , \14538 );
nor \U$28940 ( \29283 , \29280 , \29282 );
xor \U$28941 ( \29284 , \29276 , \29283 );
not \U$28942 ( \29285 , RI9873558_190);
and \U$28943 ( \29286 , \15780 , RI986fca0_69);
and \U$28944 ( \29287 , RI9873648_192, RI986ff70_75);
nor \U$28945 ( \29288 , \29286 , \29287 );
not \U$28946 ( \29289 , \29288 );
or \U$28947 ( \29290 , \29285 , \29289 );
or \U$28948 ( \29291 , \29288 , RI9873558_190);
nand \U$28949 ( \29292 , \29290 , \29291 );
xor \U$28950 ( \29293 , \29292 , \10428 );
and \U$28951 ( \29294 , \14937 , RI986fbb0_67);
and \U$28952 ( \29295 , RI986fd90_71, \14935 );
nor \U$28953 ( \29296 , \29294 , \29295 );
and \U$28954 ( \29297 , \29296 , \14539 );
not \U$28955 ( \29298 , \29296 );
and \U$28956 ( \29299 , \29298 , \14538 );
nor \U$28957 ( \29300 , \29297 , \29299 );
and \U$28958 ( \29301 , \29293 , \29300 );
and \U$28959 ( \29302 , \29292 , \10428 );
or \U$28960 ( \29303 , \29301 , \29302 );
and \U$28961 ( \29304 , \10424 , RI9870420_85);
and \U$28962 ( \29305 , RI9870510_87, \10422 );
nor \U$28963 ( \29306 , \29304 , \29305 );
and \U$28964 ( \29307 , \29306 , \9840 );
not \U$28965 ( \29308 , \29306 );
and \U$28966 ( \29309 , \29308 , \10428 );
nor \U$28967 ( \29310 , \29307 , \29309 );
xor \U$28968 ( \29311 , \29303 , \29310 );
and \U$28969 ( \29312 , \13045 , RI9870600_89);
and \U$28970 ( \29313 , RI98708d0_95, \13043 );
nor \U$28971 ( \29314 , \29312 , \29313 );
and \U$28972 ( \29315 , \29314 , \13047 );
not \U$28973 ( \29316 , \29314 );
and \U$28974 ( \29317 , \29316 , \12619 );
nor \U$28975 ( \29318 , \29315 , \29317 );
and \U$28976 ( \29319 , \12293 , RI9870240_81);
and \U$28977 ( \29320 , RI98706f0_91, \12291 );
nor \U$28978 ( \29321 , \29319 , \29320 );
and \U$28979 ( \29322 , \29321 , \11687 );
not \U$28980 ( \29323 , \29321 );
and \U$28981 ( \29324 , \29323 , \11686 );
nor \U$28982 ( \29325 , \29322 , \29324 );
xor \U$28983 ( \29326 , \29318 , \29325 );
and \U$28984 ( \29327 , \13882 , RI98707e0_93);
and \U$28985 ( \29328 , RI986fac0_65, \13880 );
nor \U$28986 ( \29329 , \29327 , \29328 );
and \U$28987 ( \29330 , \29329 , \13358 );
not \U$28988 ( \29331 , \29329 );
and \U$28989 ( \29332 , \29331 , \13359 );
nor \U$28990 ( \29333 , \29330 , \29332 );
and \U$28991 ( \29334 , \29326 , \29333 );
and \U$28992 ( \29335 , \29318 , \29325 );
or \U$28993 ( \29336 , \29334 , \29335 );
xor \U$28994 ( \29337 , \29311 , \29336 );
xor \U$28995 ( \29338 , \29284 , \29337 );
not \U$28996 ( \29339 , \29338 );
and \U$28997 ( \29340 , \15780 , RI986fd90_71);
and \U$28998 ( \29341 , RI9873648_192, RI986fca0_69);
nor \U$28999 ( \29342 , \29340 , \29341 );
not \U$29000 ( \29343 , \29342 );
not \U$29001 ( \29344 , RI9873558_190);
and \U$29002 ( \29345 , \29343 , \29344 );
and \U$29003 ( \29346 , \29342 , RI9873558_190);
nor \U$29004 ( \29347 , \29345 , \29346 );
and \U$29005 ( \29348 , \14937 , RI986fac0_65);
and \U$29006 ( \29349 , RI986fbb0_67, \14935 );
nor \U$29007 ( \29350 , \29348 , \29349 );
and \U$29008 ( \29351 , \29350 , \14538 );
not \U$29009 ( \29352 , \29350 );
and \U$29010 ( \29353 , \29352 , \14539 );
nor \U$29011 ( \29354 , \29351 , \29353 );
xor \U$29012 ( \29355 , \29347 , \29354 );
and \U$29013 ( \29356 , \13882 , RI98708d0_95);
and \U$29014 ( \29357 , RI98707e0_93, \13880 );
nor \U$29015 ( \29358 , \29356 , \29357 );
and \U$29016 ( \29359 , \29358 , \13359 );
not \U$29017 ( \29360 , \29358 );
and \U$29018 ( \29361 , \29360 , \13358 );
nor \U$29019 ( \29362 , \29359 , \29361 );
and \U$29020 ( \29363 , \29355 , \29362 );
and \U$29021 ( \29364 , \29347 , \29354 );
nor \U$29022 ( \29365 , \29363 , \29364 );
and \U$29023 ( \29366 , \11696 , RI9870510_87);
and \U$29024 ( \29367 , RI9870330_83, \11694 );
nor \U$29025 ( \29368 , \29366 , \29367 );
and \U$29026 ( \29369 , \29368 , \10965 );
not \U$29027 ( \29370 , \29368 );
and \U$29028 ( \29371 , \29370 , \11702 );
nor \U$29029 ( \29372 , \29369 , \29371 );
xor \U$29030 ( \29373 , \29365 , \29372 );
and \U$29031 ( \29374 , \12293 , RI9870330_83);
and \U$29032 ( \29375 , RI9870240_81, \12291 );
nor \U$29033 ( \29376 , \29374 , \29375 );
and \U$29034 ( \29377 , \29376 , \11686 );
not \U$29035 ( \29378 , \29376 );
and \U$29036 ( \29379 , \29378 , \11687 );
nor \U$29037 ( \29380 , \29377 , \29379 );
and \U$29038 ( \29381 , \13045 , RI98706f0_91);
and \U$29039 ( \29382 , RI9870600_89, \13043 );
nor \U$29040 ( \29383 , \29381 , \29382 );
and \U$29041 ( \29384 , \29383 , \12619 );
not \U$29042 ( \29385 , \29383 );
and \U$29043 ( \29386 , \29385 , \13047 );
nor \U$29044 ( \29387 , \29384 , \29386 );
xor \U$29045 ( \29388 , \29380 , \29387 );
and \U$29046 ( \29389 , \11696 , RI9870420_85);
and \U$29047 ( \29390 , RI9870510_87, \11694 );
nor \U$29048 ( \29391 , \29389 , \29390 );
and \U$29049 ( \29392 , \29391 , \11702 );
not \U$29050 ( \29393 , \29391 );
and \U$29051 ( \29394 , \29393 , \10965 );
nor \U$29052 ( \29395 , \29392 , \29394 );
and \U$29053 ( \29396 , \29388 , \29395 );
and \U$29054 ( \29397 , \29380 , \29387 );
nor \U$29055 ( \29398 , \29396 , \29397 );
and \U$29056 ( \29399 , \29373 , \29398 );
and \U$29057 ( \29400 , \29365 , \29372 );
or \U$29058 ( \29401 , \29399 , \29400 );
and \U$29059 ( \29402 , \11696 , RI9870330_83);
and \U$29060 ( \29403 , RI9870240_81, \11694 );
nor \U$29061 ( \29404 , \29402 , \29403 );
and \U$29062 ( \29405 , \29404 , \10965 );
not \U$29063 ( \29406 , \29404 );
and \U$29064 ( \29407 , \29406 , \11702 );
nor \U$29065 ( \29408 , \29405 , \29407 );
and \U$29066 ( \29409 , \12293 , RI98706f0_91);
and \U$29067 ( \29410 , RI9870600_89, \12291 );
nor \U$29068 ( \29411 , \29409 , \29410 );
and \U$29069 ( \29412 , \29411 , \11687 );
not \U$29070 ( \29413 , \29411 );
and \U$29071 ( \29414 , \29413 , \11686 );
nor \U$29072 ( \29415 , \29412 , \29414 );
xor \U$29073 ( \29416 , \29408 , \29415 );
and \U$29074 ( \29417 , \13045 , RI98708d0_95);
and \U$29075 ( \29418 , RI98707e0_93, \13043 );
nor \U$29076 ( \29419 , \29417 , \29418 );
and \U$29077 ( \29420 , \29419 , \13047 );
not \U$29078 ( \29421 , \29419 );
and \U$29079 ( \29422 , \29421 , \12619 );
nor \U$29080 ( \29423 , \29420 , \29422 );
xor \U$29081 ( \29424 , \29416 , \29423 );
xor \U$29082 ( \29425 , \29401 , \29424 );
nand \U$29083 ( \29426 , RI9870420_85, \10422 );
and \U$29084 ( \29427 , \29426 , \9840 );
not \U$29085 ( \29428 , \29426 );
and \U$29086 ( \29429 , \29428 , \10428 );
nor \U$29087 ( \29430 , \29427 , \29429 );
xor \U$29088 ( \29431 , \29318 , \29325 );
xor \U$29089 ( \29432 , \29431 , \29333 );
and \U$29090 ( \29433 , \29430 , \29432 );
xor \U$29091 ( \29434 , \29292 , \10428 );
xor \U$29092 ( \29435 , \29434 , \29300 );
xor \U$29093 ( \29436 , \29318 , \29325 );
xor \U$29094 ( \29437 , \29436 , \29333 );
and \U$29095 ( \29438 , \29435 , \29437 );
and \U$29096 ( \29439 , \29430 , \29435 );
or \U$29097 ( \29440 , \29433 , \29438 , \29439 );
xor \U$29098 ( \29441 , \29425 , \29440 );
not \U$29099 ( \29442 , \29441 );
or \U$29100 ( \29443 , \29339 , \29442 );
or \U$29101 ( \29444 , \29441 , \29338 );
xor \U$29102 ( \29445 , \29380 , \29387 );
xor \U$29103 ( \29446 , \29445 , \29395 );
not \U$29104 ( \29447 , RI9873558_190);
and \U$29105 ( \29448 , \15780 , RI986fbb0_67);
and \U$29106 ( \29449 , RI9873648_192, RI986fd90_71);
nor \U$29107 ( \29450 , \29448 , \29449 );
not \U$29108 ( \29451 , \29450 );
or \U$29109 ( \29452 , \29447 , \29451 );
or \U$29110 ( \29453 , \29450 , RI9873558_190);
nand \U$29111 ( \29454 , \29452 , \29453 );
and \U$29112 ( \29455 , \29454 , \11702 );
not \U$29113 ( \29456 , \29454 );
not \U$29114 ( \29457 , \11702 );
and \U$29115 ( \29458 , \29456 , \29457 );
and \U$29116 ( \29459 , \14937 , RI98707e0_93);
and \U$29117 ( \29460 , RI986fac0_65, \14935 );
nor \U$29118 ( \29461 , \29459 , \29460 );
and \U$29119 ( \29462 , \29461 , \14538 );
not \U$29120 ( \29463 , \29461 );
and \U$29121 ( \29464 , \29463 , \14539 );
nor \U$29122 ( \29465 , \29462 , \29464 );
nor \U$29123 ( \29466 , \29458 , \29465 );
nor \U$29124 ( \29467 , \29455 , \29466 );
or \U$29125 ( \29468 , \29446 , \29467 );
not \U$29126 ( \29469 , \29467 );
not \U$29127 ( \29470 , \29446 );
or \U$29128 ( \29471 , \29469 , \29470 );
and \U$29129 ( \29472 , \12293 , RI9870510_87);
and \U$29130 ( \29473 , RI9870330_83, \12291 );
nor \U$29131 ( \29474 , \29472 , \29473 );
and \U$29132 ( \29475 , \29474 , \11686 );
not \U$29133 ( \29476 , \29474 );
and \U$29134 ( \29477 , \29476 , \11687 );
nor \U$29135 ( \29478 , \29475 , \29477 );
and \U$29136 ( \29479 , \13045 , RI9870240_81);
and \U$29137 ( \29480 , RI98706f0_91, \13043 );
nor \U$29138 ( \29481 , \29479 , \29480 );
and \U$29139 ( \29482 , \29481 , \12619 );
not \U$29140 ( \29483 , \29481 );
and \U$29141 ( \29484 , \29483 , \13047 );
nor \U$29142 ( \29485 , \29482 , \29484 );
or \U$29143 ( \29486 , \29478 , \29485 );
not \U$29144 ( \29487 , \29485 );
not \U$29145 ( \29488 , \29478 );
or \U$29146 ( \29489 , \29487 , \29488 );
and \U$29147 ( \29490 , \13882 , RI9870600_89);
and \U$29148 ( \29491 , RI98708d0_95, \13880 );
nor \U$29149 ( \29492 , \29490 , \29491 );
and \U$29150 ( \29493 , \29492 , \13358 );
not \U$29151 ( \29494 , \29492 );
and \U$29152 ( \29495 , \29494 , \13359 );
nor \U$29153 ( \29496 , \29493 , \29495 );
nand \U$29154 ( \29497 , \29489 , \29496 );
nand \U$29155 ( \29498 , \29486 , \29497 );
nand \U$29156 ( \29499 , \29471 , \29498 );
nand \U$29157 ( \29500 , \29468 , \29499 );
xor \U$29158 ( \29501 , \29365 , \29372 );
xor \U$29159 ( \29502 , \29501 , \29398 );
and \U$29160 ( \29503 , \29500 , \29502 );
xor \U$29161 ( \29504 , \29318 , \29325 );
xor \U$29162 ( \29505 , \29504 , \29333 );
xor \U$29163 ( \29506 , \29430 , \29435 );
xor \U$29164 ( \29507 , \29505 , \29506 );
xor \U$29165 ( \29508 , \29365 , \29372 );
xor \U$29166 ( \29509 , \29508 , \29398 );
and \U$29167 ( \29510 , \29507 , \29509 );
and \U$29168 ( \29511 , \29500 , \29507 );
or \U$29169 ( \29512 , \29503 , \29510 , \29511 );
nand \U$29170 ( \29513 , \29444 , \29512 );
nand \U$29171 ( \29514 , \29443 , \29513 );
xor \U$29172 ( \29515 , \28897 , \28904 );
xor \U$29173 ( \29516 , \29515 , \28912 );
not \U$29174 ( \29517 , \29516 );
not \U$29175 ( \29518 , \9510 );
not \U$29176 ( \29519 , \28851 );
not \U$29177 ( \29520 , \28862 );
or \U$29178 ( \29521 , \29519 , \29520 );
or \U$29179 ( \29522 , \28862 , \28851 );
nand \U$29180 ( \29523 , \29521 , \29522 );
not \U$29181 ( \29524 , \29523 );
or \U$29182 ( \29525 , \29518 , \29524 );
or \U$29183 ( \29526 , \29523 , \9510 );
nand \U$29184 ( \29527 , \29525 , \29526 );
not \U$29185 ( \29528 , \29527 );
or \U$29186 ( \29529 , \29517 , \29528 );
or \U$29187 ( \29530 , \29527 , \29516 );
nand \U$29188 ( \29531 , \29529 , \29530 );
xor \U$29189 ( \29532 , \29303 , \29310 );
and \U$29190 ( \29533 , \29532 , \29336 );
and \U$29191 ( \29534 , \29303 , \29310 );
or \U$29192 ( \29535 , \29533 , \29534 );
xor \U$29193 ( \29536 , \29531 , \29535 );
xor \U$29194 ( \29537 , \29408 , \29415 );
and \U$29195 ( \29538 , \29537 , \29423 );
and \U$29196 ( \29539 , \29408 , \29415 );
or \U$29197 ( \29540 , \29538 , \29539 );
xor \U$29198 ( \29541 , \29267 , \29275 );
and \U$29199 ( \29542 , \29541 , \29283 );
and \U$29200 ( \29543 , \29267 , \29275 );
or \U$29201 ( \29544 , \29542 , \29543 );
xor \U$29202 ( \29545 , \29540 , \29544 );
not \U$29203 ( \29546 , \28877 );
xor \U$29204 ( \29547 , \28887 , \28871 );
not \U$29205 ( \29548 , \29547 );
or \U$29206 ( \29549 , \29546 , \29548 );
or \U$29207 ( \29550 , \29547 , \28877 );
nand \U$29208 ( \29551 , \29549 , \29550 );
xor \U$29209 ( \29552 , \29545 , \29551 );
xor \U$29210 ( \29553 , \29536 , \29552 );
and \U$29211 ( \29554 , \29284 , \29337 );
xor \U$29212 ( \29555 , \29553 , \29554 );
xor \U$29213 ( \29556 , \29401 , \29424 );
and \U$29214 ( \29557 , \29556 , \29440 );
and \U$29215 ( \29558 , \29401 , \29424 );
or \U$29216 ( \29559 , \29557 , \29558 );
xor \U$29217 ( \29560 , \29555 , \29559 );
and \U$29218 ( \29561 , \29514 , \29560 );
xor \U$29219 ( \29562 , \29560 , \29514 );
and \U$29220 ( \29563 , \13882 , RI98706f0_91);
and \U$29221 ( \29564 , RI9870600_89, \13880 );
nor \U$29222 ( \29565 , \29563 , \29564 );
and \U$29223 ( \29566 , \29565 , \13359 );
not \U$29224 ( \29567 , \29565 );
and \U$29225 ( \29568 , \29567 , \13358 );
nor \U$29226 ( \29569 , \29566 , \29568 );
not \U$29227 ( \29570 , \29569 );
and \U$29228 ( \29571 , \15780 , RI986fac0_65);
and \U$29229 ( \29572 , RI9873648_192, RI986fbb0_67);
nor \U$29230 ( \29573 , \29571 , \29572 );
not \U$29231 ( \29574 , \29573 );
not \U$29232 ( \29575 , RI9873558_190);
and \U$29233 ( \29576 , \29574 , \29575 );
and \U$29234 ( \29577 , \29573 , RI9873558_190);
nor \U$29235 ( \29578 , \29576 , \29577 );
not \U$29236 ( \29579 , \29578 );
and \U$29237 ( \29580 , \29570 , \29579 );
and \U$29238 ( \29581 , \29569 , \29578 );
and \U$29239 ( \29582 , \14937 , RI98708d0_95);
and \U$29240 ( \29583 , RI98707e0_93, \14935 );
nor \U$29241 ( \29584 , \29582 , \29583 );
and \U$29242 ( \29585 , \29584 , \14538 );
not \U$29243 ( \29586 , \29584 );
and \U$29244 ( \29587 , \29586 , \14539 );
nor \U$29245 ( \29588 , \29585 , \29587 );
nor \U$29246 ( \29589 , \29581 , \29588 );
nor \U$29247 ( \29590 , \29580 , \29589 );
nand \U$29248 ( \29591 , RI9870420_85, \11694 );
and \U$29249 ( \29592 , \29591 , \11702 );
not \U$29250 ( \29593 , \29591 );
and \U$29251 ( \29594 , \29593 , \10965 );
nor \U$29252 ( \29595 , \29592 , \29594 );
xor \U$29253 ( \29596 , \29590 , \29595 );
not \U$29254 ( \29597 , \29485 );
not \U$29255 ( \29598 , \29496 );
or \U$29256 ( \29599 , \29597 , \29598 );
or \U$29257 ( \29600 , \29485 , \29496 );
nand \U$29258 ( \29601 , \29599 , \29600 );
not \U$29259 ( \29602 , \29601 );
not \U$29260 ( \29603 , \29478 );
and \U$29261 ( \29604 , \29602 , \29603 );
and \U$29262 ( \29605 , \29601 , \29478 );
nor \U$29263 ( \29606 , \29604 , \29605 );
and \U$29264 ( \29607 , \29596 , \29606 );
and \U$29265 ( \29608 , \29590 , \29595 );
or \U$29266 ( \29609 , \29607 , \29608 );
xor \U$29267 ( \29610 , \29347 , \29354 );
xor \U$29268 ( \29611 , \29610 , \29362 );
xor \U$29269 ( \29612 , \29609 , \29611 );
not \U$29270 ( \29613 , \29467 );
not \U$29271 ( \29614 , \29498 );
or \U$29272 ( \29615 , \29613 , \29614 );
or \U$29273 ( \29616 , \29498 , \29467 );
nand \U$29274 ( \29617 , \29615 , \29616 );
not \U$29275 ( \29618 , \29617 );
not \U$29276 ( \29619 , \29446 );
and \U$29277 ( \29620 , \29618 , \29619 );
and \U$29278 ( \29621 , \29617 , \29446 );
nor \U$29279 ( \29622 , \29620 , \29621 );
xor \U$29280 ( \29623 , \29612 , \29622 );
not \U$29281 ( \29624 , \29623 );
not \U$29282 ( \29625 , RI9873558_190);
and \U$29283 ( \29626 , \15780 , RI98707e0_93);
and \U$29284 ( \29627 , RI9873648_192, RI986fac0_65);
nor \U$29285 ( \29628 , \29626 , \29627 );
not \U$29286 ( \29629 , \29628 );
or \U$29287 ( \29630 , \29625 , \29629 );
or \U$29288 ( \29631 , \29628 , RI9873558_190);
nand \U$29289 ( \29632 , \29630 , \29631 );
and \U$29290 ( \29633 , \29632 , \11686 );
not \U$29291 ( \29634 , \29632 );
not \U$29292 ( \29635 , \11686 );
and \U$29293 ( \29636 , \29634 , \29635 );
and \U$29294 ( \29637 , \14937 , RI9870600_89);
and \U$29295 ( \29638 , RI98708d0_95, \14935 );
nor \U$29296 ( \29639 , \29637 , \29638 );
and \U$29297 ( \29640 , \29639 , \14538 );
not \U$29298 ( \29641 , \29639 );
and \U$29299 ( \29642 , \29641 , \14539 );
nor \U$29300 ( \29643 , \29640 , \29642 );
nor \U$29301 ( \29644 , \29636 , \29643 );
nor \U$29302 ( \29645 , \29633 , \29644 );
and \U$29303 ( \29646 , \13045 , RI9870330_83);
and \U$29304 ( \29647 , RI9870240_81, \13043 );
nor \U$29305 ( \29648 , \29646 , \29647 );
and \U$29306 ( \29649 , \29648 , \12619 );
not \U$29307 ( \29650 , \29648 );
and \U$29308 ( \29651 , \29650 , \13047 );
nor \U$29309 ( \29652 , \29649 , \29651 );
or \U$29310 ( \29653 , \29645 , \29652 );
not \U$29311 ( \29654 , \29652 );
not \U$29312 ( \29655 , \29645 );
or \U$29313 ( \29656 , \29654 , \29655 );
and \U$29314 ( \29657 , \13882 , RI9870240_81);
and \U$29315 ( \29658 , RI98706f0_91, \13880 );
nor \U$29316 ( \29659 , \29657 , \29658 );
and \U$29317 ( \29660 , \29659 , \13358 );
not \U$29318 ( \29661 , \29659 );
and \U$29319 ( \29662 , \29661 , \13359 );
nor \U$29320 ( \29663 , \29660 , \29662 );
nand \U$29321 ( \29664 , RI9870420_85, \12291 );
and \U$29322 ( \29665 , \29664 , \11687 );
not \U$29323 ( \29666 , \29664 );
and \U$29324 ( \29667 , \29666 , \11686 );
nor \U$29325 ( \29668 , \29665 , \29667 );
xor \U$29326 ( \29669 , \29663 , \29668 );
and \U$29327 ( \29670 , \13045 , RI9870510_87);
and \U$29328 ( \29671 , RI9870330_83, \13043 );
nor \U$29329 ( \29672 , \29670 , \29671 );
and \U$29330 ( \29673 , \29672 , \13047 );
not \U$29331 ( \29674 , \29672 );
and \U$29332 ( \29675 , \29674 , \12619 );
nor \U$29333 ( \29676 , \29673 , \29675 );
and \U$29334 ( \29677 , \29669 , \29676 );
and \U$29335 ( \29678 , \29663 , \29668 );
or \U$29336 ( \29679 , \29677 , \29678 );
nand \U$29337 ( \29680 , \29656 , \29679 );
nand \U$29338 ( \29681 , \29653 , \29680 );
not \U$29339 ( \29682 , \10965 );
not \U$29340 ( \29683 , \29454 );
not \U$29341 ( \29684 , \29465 );
or \U$29342 ( \29685 , \29683 , \29684 );
or \U$29343 ( \29686 , \29465 , \29454 );
nand \U$29344 ( \29687 , \29685 , \29686 );
not \U$29345 ( \29688 , \29687 );
or \U$29346 ( \29689 , \29682 , \29688 );
or \U$29347 ( \29690 , \29687 , \10965 );
nand \U$29348 ( \29691 , \29689 , \29690 );
xor \U$29349 ( \29692 , \29681 , \29691 );
and \U$29350 ( \29693 , \12293 , RI9870420_85);
and \U$29351 ( \29694 , RI9870510_87, \12291 );
nor \U$29352 ( \29695 , \29693 , \29694 );
and \U$29353 ( \29696 , \29695 , \11687 );
not \U$29354 ( \29697 , \29695 );
and \U$29355 ( \29698 , \29697 , \11686 );
nor \U$29356 ( \29699 , \29696 , \29698 );
not \U$29357 ( \29700 , \29569 );
xor \U$29358 ( \29701 , \29578 , \29588 );
not \U$29359 ( \29702 , \29701 );
or \U$29360 ( \29703 , \29700 , \29702 );
or \U$29361 ( \29704 , \29701 , \29569 );
nand \U$29362 ( \29705 , \29703 , \29704 );
and \U$29363 ( \29706 , \29699 , \29705 );
and \U$29364 ( \29707 , \29692 , \29706 );
and \U$29365 ( \29708 , \29681 , \29691 );
or \U$29366 ( \29709 , \29707 , \29708 );
not \U$29367 ( \29710 , \29709 );
and \U$29368 ( \29711 , \29624 , \29710 );
and \U$29369 ( \29712 , \29623 , \29709 );
nor \U$29370 ( \29713 , \29711 , \29712 );
xor \U$29371 ( \29714 , \29590 , \29595 );
xor \U$29372 ( \29715 , \29714 , \29606 );
not \U$29373 ( \29716 , \29715 );
xor \U$29374 ( \29717 , \29681 , \29691 );
xor \U$29375 ( \29718 , \29717 , \29706 );
nand \U$29376 ( \29719 , \29716 , \29718 );
or \U$29377 ( \29720 , \29713 , \29719 );
xnor \U$29378 ( \29721 , \29719 , \29713 );
and \U$29379 ( \29722 , \13882 , RI9870510_87);
and \U$29380 ( \29723 , RI9870330_83, \13880 );
nor \U$29381 ( \29724 , \29722 , \29723 );
and \U$29382 ( \29725 , \29724 , \13359 );
not \U$29383 ( \29726 , \29724 );
and \U$29384 ( \29727 , \29726 , \13358 );
nor \U$29385 ( \29728 , \29725 , \29727 );
not \U$29386 ( \29729 , \29728 );
nand \U$29387 ( \29730 , RI9870420_85, \13043 );
and \U$29388 ( \29731 , \29730 , \13047 );
not \U$29389 ( \29732 , \29730 );
and \U$29390 ( \29733 , \29732 , \12619 );
nor \U$29391 ( \29734 , \29731 , \29733 );
nand \U$29392 ( \29735 , \29729 , \29734 );
not \U$29393 ( \29736 , \29735 );
and \U$29394 ( \29737 , \13045 , RI9870420_85);
and \U$29395 ( \29738 , RI9870510_87, \13043 );
nor \U$29396 ( \29739 , \29737 , \29738 );
and \U$29397 ( \29740 , \29739 , \12619 );
not \U$29398 ( \29741 , \29739 );
and \U$29399 ( \29742 , \29741 , \13047 );
nor \U$29400 ( \29743 , \29740 , \29742 );
not \U$29401 ( \29744 , \29743 );
and \U$29402 ( \29745 , \29736 , \29744 );
and \U$29403 ( \29746 , \29735 , \29743 );
not \U$29404 ( \29747 , RI9873558_190);
and \U$29405 ( \29748 , \15780 , RI9870600_89);
and \U$29406 ( \29749 , RI9873648_192, RI98708d0_95);
nor \U$29407 ( \29750 , \29748 , \29749 );
not \U$29408 ( \29751 , \29750 );
or \U$29409 ( \29752 , \29747 , \29751 );
or \U$29410 ( \29753 , \29750 , RI9873558_190);
nand \U$29411 ( \29754 , \29752 , \29753 );
xor \U$29412 ( \29755 , \29754 , \12619 );
and \U$29413 ( \29756 , \14937 , RI9870240_81);
and \U$29414 ( \29757 , RI98706f0_91, \14935 );
nor \U$29415 ( \29758 , \29756 , \29757 );
and \U$29416 ( \29759 , \29758 , \14539 );
not \U$29417 ( \29760 , \29758 );
and \U$29418 ( \29761 , \29760 , \14538 );
nor \U$29419 ( \29762 , \29759 , \29761 );
and \U$29420 ( \29763 , \29755 , \29762 );
and \U$29421 ( \29764 , \29754 , \12619 );
or \U$29422 ( \29765 , \29763 , \29764 );
not \U$29423 ( \29766 , \29765 );
nor \U$29424 ( \29767 , \29746 , \29766 );
nor \U$29425 ( \29768 , \29745 , \29767 );
not \U$29426 ( \29769 , \29768 );
not \U$29427 ( \29770 , \29632 );
not \U$29428 ( \29771 , \29643 );
or \U$29429 ( \29772 , \29770 , \29771 );
or \U$29430 ( \29773 , \29643 , \29632 );
nand \U$29431 ( \29774 , \29772 , \29773 );
and \U$29432 ( \29775 , \29774 , \11686 );
not \U$29433 ( \29776 , \29774 );
and \U$29434 ( \29777 , \29776 , \11687 );
nor \U$29435 ( \29778 , \29775 , \29777 );
and \U$29436 ( \29779 , \15780 , RI98708d0_95);
and \U$29437 ( \29780 , RI9873648_192, RI98707e0_93);
nor \U$29438 ( \29781 , \29779 , \29780 );
not \U$29439 ( \29782 , \29781 );
not \U$29440 ( \29783 , RI9873558_190);
and \U$29441 ( \29784 , \29782 , \29783 );
and \U$29442 ( \29785 , \29781 , RI9873558_190);
nor \U$29443 ( \29786 , \29784 , \29785 );
and \U$29444 ( \29787 , \14937 , RI98706f0_91);
and \U$29445 ( \29788 , RI9870600_89, \14935 );
nor \U$29446 ( \29789 , \29787 , \29788 );
and \U$29447 ( \29790 , \29789 , \14538 );
not \U$29448 ( \29791 , \29789 );
and \U$29449 ( \29792 , \29791 , \14539 );
nor \U$29450 ( \29793 , \29790 , \29792 );
xor \U$29451 ( \29794 , \29786 , \29793 );
and \U$29452 ( \29795 , \13882 , RI9870330_83);
and \U$29453 ( \29796 , RI9870240_81, \13880 );
nor \U$29454 ( \29797 , \29795 , \29796 );
and \U$29455 ( \29798 , \29797 , \13359 );
not \U$29456 ( \29799 , \29797 );
and \U$29457 ( \29800 , \29799 , \13358 );
nor \U$29458 ( \29801 , \29798 , \29800 );
and \U$29459 ( \29802 , \29794 , \29801 );
and \U$29460 ( \29803 , \29786 , \29793 );
nor \U$29461 ( \29804 , \29802 , \29803 );
xor \U$29462 ( \29805 , \29778 , \29804 );
xor \U$29463 ( \29806 , \29663 , \29668 );
xor \U$29464 ( \29807 , \29806 , \29676 );
xor \U$29465 ( \29808 , \29805 , \29807 );
nand \U$29466 ( \29809 , \29769 , \29808 );
not \U$29467 ( \29810 , \29645 );
not \U$29468 ( \29811 , \29679 );
or \U$29469 ( \29812 , \29810 , \29811 );
or \U$29470 ( \29813 , \29679 , \29645 );
nand \U$29471 ( \29814 , \29812 , \29813 );
not \U$29472 ( \29815 , \29814 );
not \U$29473 ( \29816 , \29652 );
and \U$29474 ( \29817 , \29815 , \29816 );
and \U$29475 ( \29818 , \29814 , \29652 );
nor \U$29476 ( \29819 , \29817 , \29818 );
not \U$29477 ( \29820 , \29819 );
xor \U$29478 ( \29821 , \29778 , \29804 );
and \U$29479 ( \29822 , \29821 , \29807 );
and \U$29480 ( \29823 , \29778 , \29804 );
or \U$29481 ( \29824 , \29822 , \29823 );
not \U$29482 ( \29825 , \29824 );
and \U$29483 ( \29826 , \29820 , \29825 );
and \U$29484 ( \29827 , \29819 , \29824 );
nor \U$29485 ( \29828 , \29826 , \29827 );
not \U$29486 ( \29829 , \29828 );
xor \U$29487 ( \29830 , \29699 , \29705 );
not \U$29488 ( \29831 , \29830 );
and \U$29489 ( \29832 , \29829 , \29831 );
and \U$29490 ( \29833 , \29828 , \29830 );
nor \U$29491 ( \29834 , \29832 , \29833 );
xor \U$29492 ( \29835 , \29809 , \29834 );
xor \U$29493 ( \29836 , \29754 , \12619 );
xor \U$29494 ( \29837 , \29836 , \29762 );
not \U$29495 ( \29838 , \29734 );
not \U$29496 ( \29839 , \29728 );
or \U$29497 ( \29840 , \29838 , \29839 );
or \U$29498 ( \29841 , \29728 , \29734 );
nand \U$29499 ( \29842 , \29840 , \29841 );
and \U$29500 ( \29843 , \29837 , \29842 );
not \U$29501 ( \29844 , \29837 );
not \U$29502 ( \29845 , \29842 );
and \U$29503 ( \29846 , \29844 , \29845 );
and \U$29504 ( \29847 , \13882 , RI9870420_85);
and \U$29505 ( \29848 , RI9870510_87, \13880 );
nor \U$29506 ( \29849 , \29847 , \29848 );
and \U$29507 ( \29850 , \29849 , \13359 );
not \U$29508 ( \29851 , \29849 );
and \U$29509 ( \29852 , \29851 , \13358 );
nor \U$29510 ( \29853 , \29850 , \29852 );
and \U$29511 ( \29854 , \15780 , RI98706f0_91);
and \U$29512 ( \29855 , RI9873648_192, RI9870600_89);
nor \U$29513 ( \29856 , \29854 , \29855 );
not \U$29514 ( \29857 , \29856 );
not \U$29515 ( \29858 , RI9873558_190);
and \U$29516 ( \29859 , \29857 , \29858 );
and \U$29517 ( \29860 , \29856 , RI9873558_190);
nor \U$29518 ( \29861 , \29859 , \29860 );
xor \U$29519 ( \29862 , \29853 , \29861 );
and \U$29520 ( \29863 , \14937 , RI9870330_83);
and \U$29521 ( \29864 , RI9870240_81, \14935 );
nor \U$29522 ( \29865 , \29863 , \29864 );
and \U$29523 ( \29866 , \29865 , \14538 );
not \U$29524 ( \29867 , \29865 );
and \U$29525 ( \29868 , \29867 , \14539 );
nor \U$29526 ( \29869 , \29866 , \29868 );
and \U$29527 ( \29870 , \29862 , \29869 );
and \U$29528 ( \29871 , \29853 , \29861 );
or \U$29529 ( \29872 , \29870 , \29871 );
nor \U$29530 ( \29873 , \29846 , \29872 );
nor \U$29531 ( \29874 , \29843 , \29873 );
not \U$29532 ( \29875 , \29743 );
not \U$29533 ( \29876 , \29735 );
not \U$29534 ( \29877 , \29765 );
or \U$29535 ( \29878 , \29876 , \29877 );
or \U$29536 ( \29879 , \29765 , \29735 );
nand \U$29537 ( \29880 , \29878 , \29879 );
not \U$29538 ( \29881 , \29880 );
or \U$29539 ( \29882 , \29875 , \29881 );
or \U$29540 ( \29883 , \29880 , \29743 );
nand \U$29541 ( \29884 , \29882 , \29883 );
not \U$29542 ( \29885 , \29884 );
xor \U$29543 ( \29886 , \29786 , \29793 );
xor \U$29544 ( \29887 , \29886 , \29801 );
not \U$29545 ( \29888 , \29887 );
and \U$29546 ( \29889 , \29885 , \29888 );
and \U$29547 ( \29890 , \29884 , \29887 );
nor \U$29548 ( \29891 , \29889 , \29890 );
xor \U$29549 ( \29892 , \29874 , \29891 );
nand \U$29550 ( \29893 , RI9870420_85, \13880 );
and \U$29551 ( \29894 , \29893 , \13359 );
not \U$29552 ( \29895 , \29893 );
and \U$29553 ( \29896 , \29895 , \13358 );
nor \U$29554 ( \29897 , \29894 , \29896 );
not \U$29555 ( \29898 , \29897 );
not \U$29556 ( \29899 , RI9873558_190);
and \U$29557 ( \29900 , \15780 , RI9870240_81);
and \U$29558 ( \29901 , RI9873648_192, RI98706f0_91);
nor \U$29559 ( \29902 , \29900 , \29901 );
not \U$29560 ( \29903 , \29902 );
or \U$29561 ( \29904 , \29899 , \29903 );
or \U$29562 ( \29905 , \29902 , RI9873558_190);
nand \U$29563 ( \29906 , \29904 , \29905 );
xor \U$29564 ( \29907 , \29906 , \13359 );
and \U$29565 ( \29908 , \14937 , RI9870510_87);
and \U$29566 ( \29909 , RI9870330_83, \14935 );
nor \U$29567 ( \29910 , \29908 , \29909 );
and \U$29568 ( \29911 , \29910 , \14539 );
not \U$29569 ( \29912 , \29910 );
and \U$29570 ( \29913 , \29912 , \14538 );
nor \U$29571 ( \29914 , \29911 , \29913 );
xor \U$29572 ( \29915 , \29907 , \29914 );
nand \U$29573 ( \29916 , \29898 , \29915 );
xor \U$29574 ( \29917 , \29853 , \29861 );
xor \U$29575 ( \29918 , \29917 , \29869 );
not \U$29576 ( \29919 , \29918 );
xor \U$29577 ( \29920 , \29906 , \13359 );
and \U$29578 ( \29921 , \29920 , \29914 );
and \U$29579 ( \29922 , \29906 , \13359 );
or \U$29580 ( \29923 , \29921 , \29922 );
not \U$29581 ( \29924 , \29923 );
and \U$29582 ( \29925 , \29919 , \29924 );
and \U$29583 ( \29926 , \29918 , \29923 );
nor \U$29584 ( \29927 , \29925 , \29926 );
xor \U$29585 ( \29928 , \29916 , \29927 );
and \U$29586 ( \29929 , \14937 , RI9870420_85);
and \U$29587 ( \29930 , RI9870510_87, \14935 );
nor \U$29588 ( \29931 , \29929 , \29930 );
and \U$29589 ( \29932 , \29931 , \14539 );
not \U$29590 ( \29933 , \29931 );
and \U$29591 ( \29934 , \29933 , \14538 );
nor \U$29592 ( \29935 , \29932 , \29934 );
not \U$29593 ( \29936 , \29935 );
and \U$29594 ( \29937 , \15780 , RI9870330_83);
and \U$29595 ( \29938 , RI9873648_192, RI9870240_81);
nor \U$29596 ( \29939 , \29937 , \29938 );
not \U$29597 ( \29940 , \29939 );
not \U$29598 ( \29941 , RI9873558_190);
and \U$29599 ( \29942 , \29940 , \29941 );
and \U$29600 ( \29943 , \29939 , RI9873558_190);
nor \U$29601 ( \29944 , \29942 , \29943 );
nor \U$29602 ( \29945 , \29936 , \29944 );
not \U$29603 ( \29946 , \29897 );
not \U$29604 ( \29947 , \29915 );
or \U$29605 ( \29948 , \29946 , \29947 );
or \U$29606 ( \29949 , \29915 , \29897 );
nand \U$29607 ( \29950 , \29948 , \29949 );
xor \U$29608 ( \29951 , \29945 , \29950 );
not \U$29609 ( \29952 , RI9873558_190);
and \U$29610 ( \29953 , \15780 , RI9870510_87);
and \U$29611 ( \29954 , RI9873648_192, RI9870330_83);
nor \U$29612 ( \29955 , \29953 , \29954 );
not \U$29613 ( \29956 , \29955 );
or \U$29614 ( \29957 , \29952 , \29956 );
or \U$29615 ( \29958 , \29955 , RI9873558_190);
nand \U$29616 ( \29959 , \29957 , \29958 );
nand \U$29617 ( \29960 , \14538 , \29959 );
not \U$29618 ( \29961 , \29935 );
not \U$29619 ( \29962 , \29944 );
and \U$29620 ( \29963 , \29961 , \29962 );
and \U$29621 ( \29964 , \29935 , \29944 );
nor \U$29622 ( \29965 , \29963 , \29964 );
xnor \U$29623 ( \29966 , \29960 , \29965 );
nand \U$29624 ( \29967 , RI9870420_85, \14935 );
and \U$29625 ( \29968 , \29967 , \14539 );
not \U$29626 ( \29969 , \29967 );
and \U$29627 ( \29970 , \29969 , \14538 );
nor \U$29628 ( \29971 , \29968 , \29970 );
and \U$29629 ( \29972 , \29959 , \14538 );
not \U$29630 ( \29973 , \29959 );
and \U$29631 ( \29974 , \29973 , \14539 );
nor \U$29632 ( \29975 , \29972 , \29974 );
xor \U$29633 ( \29976 , \29971 , \29975 );
and \U$29634 ( \29977 , \15780 , RI9870420_85);
and \U$29635 ( \29978 , RI9873648_192, RI9870510_87);
nor \U$29636 ( \29979 , \29977 , \29978 );
not \U$29637 ( \29980 , \29979 );
not \U$29638 ( \29981 , RI9873558_190);
and \U$29639 ( \29982 , \29980 , \29981 );
and \U$29640 ( \29983 , \29979 , RI9873558_190);
nor \U$29641 ( \29984 , \29982 , \29983 );
nand \U$29642 ( \29985 , RI9870420_85, RI9873648_192);
nand \U$29643 ( \29986 , RI9873558_190, \29985 );
nor \U$29644 ( \29987 , \29984 , \29986 );
and \U$29645 ( \29988 , \29976 , \29987 );
and \U$29646 ( \29989 , \29971 , \29975 );
nor \U$29647 ( \29990 , \29988 , \29989 );
or \U$29648 ( \29991 , \29966 , \29990 );
or \U$29649 ( \29992 , \29960 , \29965 );
nand \U$29650 ( \29993 , \29991 , \29992 );
and \U$29651 ( \29994 , \29951 , \29993 );
and \U$29652 ( \29995 , \29945 , \29950 );
nor \U$29653 ( \29996 , \29994 , \29995 );
and \U$29654 ( \29997 , \29928 , \29996 );
and \U$29655 ( \29998 , \29916 , \29927 );
nor \U$29656 ( \29999 , \29997 , \29998 );
not \U$29657 ( \30000 , \29923 );
nor \U$29658 ( \30001 , \30000 , \29918 );
not \U$29659 ( \30002 , \29842 );
not \U$29660 ( \30003 , \29837 );
not \U$29661 ( \30004 , \29872 );
and \U$29662 ( \30005 , \30003 , \30004 );
and \U$29663 ( \30006 , \29837 , \29872 );
nor \U$29664 ( \30007 , \30005 , \30006 );
not \U$29665 ( \30008 , \30007 );
or \U$29666 ( \30009 , \30002 , \30008 );
or \U$29667 ( \30010 , \30007 , \29842 );
nand \U$29668 ( \30011 , \30009 , \30010 );
xor \U$29669 ( \30012 , \30001 , \30011 );
and \U$29670 ( \30013 , \29999 , \30012 );
and \U$29671 ( \30014 , \30001 , \30011 );
nor \U$29672 ( \30015 , \30013 , \30014 );
and \U$29673 ( \30016 , \29892 , \30015 );
and \U$29674 ( \30017 , \29874 , \29891 );
nor \U$29675 ( \30018 , \30016 , \30017 );
not \U$29676 ( \30019 , \29884 );
nor \U$29677 ( \30020 , \30019 , \29887 );
not \U$29678 ( \30021 , \29768 );
not \U$29679 ( \30022 , \29808 );
or \U$29680 ( \30023 , \30021 , \30022 );
or \U$29681 ( \30024 , \29808 , \29768 );
nand \U$29682 ( \30025 , \30023 , \30024 );
xor \U$29683 ( \30026 , \30020 , \30025 );
and \U$29684 ( \30027 , \30018 , \30026 );
and \U$29685 ( \30028 , \30020 , \30025 );
nor \U$29686 ( \30029 , \30027 , \30028 );
and \U$29687 ( \30030 , \29835 , \30029 );
and \U$29688 ( \30031 , \29809 , \29834 );
nor \U$29689 ( \30032 , \30030 , \30031 );
not \U$29690 ( \30033 , \29830 );
or \U$29691 ( \30034 , \29819 , \30033 );
not \U$29692 ( \30035 , \30033 );
not \U$29693 ( \30036 , \29819 );
or \U$29694 ( \30037 , \30035 , \30036 );
nand \U$29695 ( \30038 , \30037 , \29824 );
nand \U$29696 ( \30039 , \30034 , \30038 );
not \U$29697 ( \30040 , \29715 );
not \U$29698 ( \30041 , \29718 );
or \U$29699 ( \30042 , \30040 , \30041 );
or \U$29700 ( \30043 , \29718 , \29715 );
nand \U$29701 ( \30044 , \30042 , \30043 );
xor \U$29702 ( \30045 , \30039 , \30044 );
and \U$29703 ( \30046 , \30032 , \30045 );
and \U$29704 ( \30047 , \30039 , \30044 );
nor \U$29705 ( \30048 , \30046 , \30047 );
or \U$29706 ( \30049 , \29721 , \30048 );
nand \U$29707 ( \30050 , \29720 , \30049 );
not \U$29708 ( \30051 , \29709 );
nor \U$29709 ( \30052 , \30051 , \29623 );
xor \U$29710 ( \30053 , \29609 , \29611 );
and \U$29711 ( \30054 , \30053 , \29622 );
and \U$29712 ( \30055 , \29609 , \29611 );
or \U$29713 ( \30056 , \30054 , \30055 );
not \U$29714 ( \30057 , \30056 );
xor \U$29715 ( \30058 , \29365 , \29372 );
xor \U$29716 ( \30059 , \30058 , \29398 );
xor \U$29717 ( \30060 , \29500 , \29507 );
xor \U$29718 ( \30061 , \30059 , \30060 );
not \U$29719 ( \30062 , \30061 );
or \U$29720 ( \30063 , \30057 , \30062 );
or \U$29721 ( \30064 , \30061 , \30056 );
nand \U$29722 ( \30065 , \30063 , \30064 );
xor \U$29723 ( \30066 , \30052 , \30065 );
and \U$29724 ( \30067 , \30050 , \30066 );
and \U$29725 ( \30068 , \30052 , \30065 );
nor \U$29726 ( \30069 , \30067 , \30068 );
not \U$29727 ( \30070 , \30056 );
nand \U$29728 ( \30071 , \30070 , \30061 );
xnor \U$29729 ( \30072 , \29512 , \29441 );
not \U$29730 ( \30073 , \30072 );
not \U$29731 ( \30074 , \29338 );
and \U$29732 ( \30075 , \30073 , \30074 );
and \U$29733 ( \30076 , \30072 , \29338 );
nor \U$29734 ( \30077 , \30075 , \30076 );
xnor \U$29735 ( \30078 , \30071 , \30077 );
or \U$29736 ( \30079 , \30069 , \30078 );
or \U$29737 ( \30080 , \30071 , \30077 );
nand \U$29738 ( \30081 , \30079 , \30080 );
and \U$29739 ( \30082 , \29562 , \30081 );
nor \U$29740 ( \30083 , \29561 , \30082 );
xor \U$29741 ( \30084 , \28864 , \28889 );
xor \U$29742 ( \30085 , \30084 , \28915 );
not \U$29743 ( \30086 , \30085 );
xor \U$29744 ( \30087 , \29531 , \29535 );
and \U$29745 ( \30088 , \30087 , \29552 );
and \U$29746 ( \30089 , \29531 , \29535 );
or \U$29747 ( \30090 , \30088 , \30089 );
not \U$29748 ( \30091 , \30090 );
or \U$29749 ( \30092 , \30086 , \30091 );
or \U$29750 ( \30093 , \30090 , \30085 );
nand \U$29751 ( \30094 , \30092 , \30093 );
not \U$29752 ( \30095 , \30094 );
xor \U$29753 ( \30096 , \29540 , \29544 );
and \U$29754 ( \30097 , \30096 , \29551 );
and \U$29755 ( \30098 , \29540 , \29544 );
nor \U$29756 ( \30099 , \30097 , \30098 );
not \U$29757 ( \30100 , \29516 );
nand \U$29758 ( \30101 , \30100 , \29527 );
xor \U$29759 ( \30102 , \30099 , \30101 );
xnor \U$29760 ( \30103 , \28979 , \29006 );
not \U$29761 ( \30104 , \30103 );
not \U$29762 ( \30105 , \28955 );
and \U$29763 ( \30106 , \30104 , \30105 );
and \U$29764 ( \30107 , \30103 , \28955 );
nor \U$29765 ( \30108 , \30106 , \30107 );
xor \U$29766 ( \30109 , \30102 , \30108 );
not \U$29767 ( \30110 , \30109 );
and \U$29768 ( \30111 , \30095 , \30110 );
and \U$29769 ( \30112 , \30094 , \30109 );
nor \U$29770 ( \30113 , \30111 , \30112 );
xor \U$29771 ( \30114 , \29553 , \29554 );
and \U$29772 ( \30115 , \30114 , \29559 );
and \U$29773 ( \30116 , \29553 , \29554 );
nor \U$29774 ( \30117 , \30115 , \30116 );
xnor \U$29775 ( \30118 , \30113 , \30117 );
or \U$29776 ( \30119 , \30083 , \30118 );
or \U$29777 ( \30120 , \30113 , \30117 );
nand \U$29778 ( \30121 , \30119 , \30120 );
or \U$29779 ( \30122 , \30109 , \30085 );
not \U$29780 ( \30123 , \30085 );
not \U$29781 ( \30124 , \30109 );
or \U$29782 ( \30125 , \30123 , \30124 );
nand \U$29783 ( \30126 , \30125 , \30090 );
nand \U$29784 ( \30127 , \30122 , \30126 );
xor \U$29785 ( \30128 , \29084 , \29095 );
not \U$29786 ( \30129 , \30128 );
xor \U$29787 ( \30130 , \30099 , \30101 );
and \U$29788 ( \30131 , \30130 , \30108 );
and \U$29789 ( \30132 , \30099 , \30101 );
or \U$29790 ( \30133 , \30131 , \30132 );
not \U$29791 ( \30134 , \30133 );
xor \U$29792 ( \30135 , \28918 , \28935 );
xor \U$29793 ( \30136 , \30135 , \29008 );
not \U$29794 ( \30137 , \30136 );
and \U$29795 ( \30138 , \30134 , \30137 );
and \U$29796 ( \30139 , \30133 , \30136 );
nor \U$29797 ( \30140 , \30138 , \30139 );
not \U$29798 ( \30141 , \30140 );
or \U$29799 ( \30142 , \30129 , \30141 );
or \U$29800 ( \30143 , \30140 , \30128 );
nand \U$29801 ( \30144 , \30142 , \30143 );
xor \U$29802 ( \30145 , \30127 , \30144 );
and \U$29803 ( \30146 , \30121 , \30145 );
and \U$29804 ( \30147 , \30127 , \30144 );
nor \U$29805 ( \30148 , \30146 , \30147 );
and \U$29806 ( \30149 , \30136 , \30128 );
not \U$29807 ( \30150 , \30136 );
not \U$29808 ( \30151 , \30128 );
and \U$29809 ( \30152 , \30150 , \30151 );
nor \U$29810 ( \30153 , \30152 , \30133 );
nor \U$29811 ( \30154 , \30149 , \30153 );
not \U$29812 ( \30155 , \29254 );
not \U$29813 ( \30156 , \29257 );
and \U$29814 ( \30157 , \30155 , \30156 );
and \U$29815 ( \30158 , \29254 , \29257 );
nor \U$29816 ( \30159 , \30157 , \30158 );
xnor \U$29817 ( \30160 , \30154 , \30159 );
or \U$29818 ( \30161 , \30148 , \30160 );
or \U$29819 ( \30162 , \30154 , \30159 );
nand \U$29820 ( \30163 , \30161 , \30162 );
and \U$29821 ( \30164 , \29260 , \30163 );
nor \U$29822 ( \30165 , \29259 , \30164 );
not \U$29823 ( \30166 , \29248 );
nand \U$29824 ( \30167 , \30166 , \29099 );
xor \U$29825 ( \30168 , \29217 , \29222 );
xor \U$29826 ( \30169 , \30168 , \29225 );
and \U$29827 ( \30170 , \29228 , \30169 );
xor \U$29828 ( \30171 , \29217 , \29222 );
xor \U$29829 ( \30172 , \30171 , \29225 );
and \U$29830 ( \30173 , \29242 , \30172 );
and \U$29831 ( \30174 , \29228 , \29242 );
or \U$29832 ( \30175 , \30170 , \30173 , \30174 );
xor \U$29833 ( \30176 , \28324 , \28331 );
xor \U$29834 ( \30177 , \30176 , \28339 );
xor \U$29835 ( \30178 , \28802 , \28807 );
xor \U$29836 ( \30179 , \30177 , \30178 );
xor \U$29837 ( \30180 , \30175 , \30179 );
xor \U$29838 ( \30181 , \29198 , \29200 );
and \U$29839 ( \30182 , \30181 , \29207 );
and \U$29840 ( \30183 , \29198 , \29200 );
or \U$29841 ( \30184 , \30182 , \30183 );
xor \U$29842 ( \30185 , \30180 , \30184 );
not \U$29843 ( \30186 , \29208 );
not \U$29844 ( \30187 , \29244 );
or \U$29845 ( \30188 , \30186 , \30187 );
or \U$29846 ( \30189 , \29244 , \29208 );
nand \U$29847 ( \30190 , \30189 , \29194 );
nand \U$29848 ( \30191 , \30188 , \30190 );
xnor \U$29849 ( \30192 , \30185 , \30191 );
not \U$29850 ( \30193 , \30192 );
xor \U$29851 ( \30194 , \28746 , \28765 );
xor \U$29852 ( \30195 , \30194 , \28791 );
xor \U$29853 ( \30196 , \29217 , \29222 );
and \U$29854 ( \30197 , \30196 , \29225 );
and \U$29855 ( \30198 , \29217 , \29222 );
or \U$29856 ( \30199 , \30197 , \30198 );
xor \U$29857 ( \30200 , \28349 , \28357 );
xor \U$29858 ( \30201 , \30200 , \28365 );
xor \U$29859 ( \30202 , \30199 , \30201 );
xor \U$29860 ( \30203 , \29232 , \29236 );
and \U$29861 ( \30204 , \30203 , \29241 );
and \U$29862 ( \30205 , \29232 , \29236 );
or \U$29863 ( \30206 , \30204 , \30205 );
xor \U$29864 ( \30207 , \30202 , \30206 );
xor \U$29865 ( \30208 , \30195 , \30207 );
not \U$29866 ( \30209 , \30208 );
and \U$29867 ( \30210 , \30193 , \30209 );
and \U$29868 ( \30211 , \30192 , \30208 );
nor \U$29869 ( \30212 , \30210 , \30211 );
xnor \U$29870 ( \30213 , \30167 , \30212 );
or \U$29871 ( \30214 , \30165 , \30213 );
or \U$29872 ( \30215 , \30167 , \30212 );
nand \U$29873 ( \30216 , \30214 , \30215 );
not \U$29874 ( \30217 , \30208 );
not \U$29875 ( \30218 , \30185 );
or \U$29876 ( \30219 , \30217 , \30218 );
or \U$29877 ( \30220 , \30185 , \30208 );
nand \U$29878 ( \30221 , \30220 , \30191 );
nand \U$29879 ( \30222 , \30219 , \30221 );
xor \U$29880 ( \30223 , \28831 , \28835 );
xor \U$29881 ( \30224 , \30199 , \30201 );
and \U$29882 ( \30225 , \30224 , \30206 );
and \U$29883 ( \30226 , \30199 , \30201 );
or \U$29884 ( \30227 , \30225 , \30226 );
xor \U$29885 ( \30228 , \30223 , \30227 );
xor \U$29886 ( \30229 , \28721 , \28794 );
xor \U$29887 ( \30230 , \30229 , \28812 );
xor \U$29888 ( \30231 , \30228 , \30230 );
and \U$29889 ( \30232 , \30195 , \30207 );
xor \U$29890 ( \30233 , \30231 , \30232 );
xor \U$29891 ( \30234 , \30175 , \30179 );
and \U$29892 ( \30235 , \30234 , \30184 );
and \U$29893 ( \30236 , \30175 , \30179 );
or \U$29894 ( \30237 , \30235 , \30236 );
xor \U$29895 ( \30238 , \30233 , \30237 );
xor \U$29896 ( \30239 , \30222 , \30238 );
and \U$29897 ( \30240 , \30216 , \30239 );
and \U$29898 ( \30241 , \30222 , \30238 );
nor \U$29899 ( \30242 , \30240 , \30241 );
xor \U$29900 ( \30243 , \30231 , \30232 );
and \U$29901 ( \30244 , \30243 , \30237 );
and \U$29902 ( \30245 , \30231 , \30232 );
nor \U$29903 ( \30246 , \30244 , \30245 );
xor \U$29904 ( \30247 , \30223 , \30227 );
and \U$29905 ( \30248 , \30247 , \30230 );
and \U$29906 ( \30249 , \30223 , \30227 );
or \U$29907 ( \30250 , \30248 , \30249 );
not \U$29908 ( \30251 , \30250 );
not \U$29909 ( \30252 , \28836 );
not \U$29910 ( \30253 , \28815 );
or \U$29911 ( \30254 , \30252 , \30253 );
or \U$29912 ( \30255 , \28815 , \28836 );
nand \U$29913 ( \30256 , \30254 , \30255 );
not \U$29914 ( \30257 , \30256 );
not \U$29915 ( \30258 , \28825 );
and \U$29916 ( \30259 , \30257 , \30258 );
and \U$29917 ( \30260 , \30256 , \28825 );
nor \U$29918 ( \30261 , \30259 , \30260 );
not \U$29919 ( \30262 , \30261 );
and \U$29920 ( \30263 , \30251 , \30262 );
and \U$29921 ( \30264 , \30250 , \30261 );
nor \U$29922 ( \30265 , \30263 , \30264 );
not \U$29923 ( \30266 , \28717 );
not \U$29924 ( \30267 , \28714 );
and \U$29925 ( \30268 , \30266 , \30267 );
and \U$29926 ( \30269 , \28717 , \28714 );
nor \U$29927 ( \30270 , \30268 , \30269 );
xnor \U$29928 ( \30271 , \30265 , \30270 );
xnor \U$29929 ( \30272 , \30246 , \30271 );
or \U$29930 ( \30273 , \30242 , \30272 );
or \U$29931 ( \30274 , \30246 , \30271 );
nand \U$29932 ( \30275 , \30273 , \30274 );
or \U$29933 ( \30276 , \30261 , \30270 );
not \U$29934 ( \30277 , \30270 );
not \U$29935 ( \30278 , \30261 );
or \U$29936 ( \30279 , \30277 , \30278 );
nand \U$29937 ( \30280 , \30279 , \30250 );
nand \U$29938 ( \30281 , \30276 , \30280 );
xor \U$29939 ( \30282 , \28712 , \28718 );
xor \U$29940 ( \30283 , \30282 , \28838 );
xor \U$29941 ( \30284 , \30281 , \30283 );
and \U$29942 ( \30285 , \30275 , \30284 );
and \U$29943 ( \30286 , \30281 , \30283 );
nor \U$29944 ( \30287 , \30285 , \30286 );
or \U$29945 ( \30288 , \28843 , \30287 );
nand \U$29946 ( \30289 , \28842 , \30288 );
not \U$29947 ( \30290 , \28704 );
or \U$29948 ( \30291 , \30290 , \28676 );
not \U$29949 ( \30292 , \28676 );
not \U$29950 ( \30293 , \30290 );
or \U$29951 ( \30294 , \30292 , \30293 );
nand \U$29952 ( \30295 , \30294 , \28650 );
nand \U$29953 ( \30296 , \30291 , \30295 );
xor \U$29954 ( \30297 , \28173 , \28192 );
xor \U$29955 ( \30298 , \30297 , \28218 );
and \U$29956 ( \30299 , \28697 , \30298 );
xor \U$29957 ( \30300 , \28173 , \28192 );
xor \U$29958 ( \30301 , \30300 , \28218 );
and \U$29959 ( \30302 , \28701 , \30301 );
and \U$29960 ( \30303 , \28697 , \28701 );
or \U$29961 ( \30304 , \30299 , \30302 , \30303 );
or \U$29962 ( \30305 , \28665 , \28672 );
not \U$29963 ( \30306 , \28672 );
not \U$29964 ( \30307 , \28665 );
or \U$29965 ( \30308 , \30306 , \30307 );
nand \U$29966 ( \30309 , \30308 , \28655 );
nand \U$29967 ( \30310 , \30305 , \30309 );
xor \U$29968 ( \30311 , \30304 , \30310 );
xor \U$29969 ( \30312 , \28028 , \28029 );
xor \U$29970 ( \30313 , \30312 , \28032 );
xor \U$29971 ( \30314 , \28270 , \28277 );
xor \U$29972 ( \30315 , \30313 , \30314 );
xor \U$29973 ( \30316 , \30311 , \30315 );
xor \U$29974 ( \30317 , \28221 , \28226 );
xor \U$29975 ( \30318 , \30317 , \28262 );
xor \U$29976 ( \30319 , \30316 , \30318 );
xor \U$29977 ( \30320 , \28689 , \28693 );
and \U$29978 ( \30321 , \30320 , \28703 );
and \U$29979 ( \30322 , \28689 , \28693 );
or \U$29980 ( \30323 , \30321 , \30322 );
xor \U$29981 ( \30324 , \30319 , \30323 );
xor \U$29982 ( \30325 , \30296 , \30324 );
and \U$29983 ( \30326 , \30289 , \30325 );
and \U$29984 ( \30327 , \30296 , \30324 );
nor \U$29985 ( \30328 , \30326 , \30327 );
xor \U$29986 ( \30329 , \30316 , \30318 );
and \U$29987 ( \30330 , \30329 , \30323 );
and \U$29988 ( \30331 , \30316 , \30318 );
nor \U$29989 ( \30332 , \30330 , \30331 );
xor \U$29990 ( \30333 , \30304 , \30310 );
and \U$29991 ( \30334 , \30333 , \30315 );
and \U$29992 ( \30335 , \30304 , \30310 );
nor \U$29993 ( \30336 , \30334 , \30335 );
not \U$29994 ( \30337 , \30336 );
xor \U$29995 ( \30338 , \28265 , \28267 );
xor \U$29996 ( \30339 , \30338 , \28282 );
not \U$29997 ( \30340 , \30339 );
or \U$29998 ( \30341 , \30337 , \30340 );
or \U$29999 ( \30342 , \30339 , \30336 );
nand \U$30000 ( \30343 , \30341 , \30342 );
not \U$30001 ( \30344 , \30343 );
not \U$30002 ( \30345 , \28146 );
not \U$30003 ( \30346 , \28143 );
and \U$30004 ( \30347 , \30345 , \30346 );
and \U$30005 ( \30348 , \28146 , \28143 );
nor \U$30006 ( \30349 , \30347 , \30348 );
not \U$30007 ( \30350 , \30349 );
and \U$30008 ( \30351 , \30344 , \30350 );
and \U$30009 ( \30352 , \30343 , \30349 );
nor \U$30010 ( \30353 , \30351 , \30352 );
xnor \U$30011 ( \30354 , \30332 , \30353 );
or \U$30012 ( \30355 , \30328 , \30354 );
or \U$30013 ( \30356 , \30332 , \30353 );
nand \U$30014 ( \30357 , \30355 , \30356 );
not \U$30015 ( \30358 , \30339 );
or \U$30016 ( \30359 , \30358 , \30349 );
and \U$30017 ( \30360 , \30358 , \30349 );
nor \U$30018 ( \30361 , \30360 , \30336 );
not \U$30019 ( \30362 , \30361 );
nand \U$30020 ( \30363 , \30359 , \30362 );
not \U$30021 ( \30364 , \28303 );
not \U$30022 ( \30365 , \28314 );
or \U$30023 ( \30366 , \30364 , \30365 );
or \U$30024 ( \30367 , \28314 , \28303 );
nand \U$30025 ( \30368 , \30366 , \30367 );
xor \U$30026 ( \30369 , \30363 , \30368 );
and \U$30027 ( \30370 , \30357 , \30369 );
and \U$30028 ( \30371 , \30363 , \30368 );
nor \U$30029 ( \30372 , \30370 , \30371 );
or \U$30030 ( \30373 , \28317 , \30372 );
nand \U$30031 ( \30374 , \28316 , \30373 );
not \U$30032 ( \30375 , \28137 );
nor \U$30033 ( \30376 , \30375 , \28289 );
xor \U$30034 ( \30377 , \27765 , \27767 );
xor \U$30035 ( \30378 , \27947 , \27949 );
xor \U$30036 ( \30379 , \30378 , \27952 );
and \U$30037 ( \30380 , \28133 , \30379 );
xor \U$30038 ( \30381 , \27947 , \27949 );
xor \U$30039 ( \30382 , \30381 , \27952 );
and \U$30040 ( \30383 , \28135 , \30382 );
and \U$30041 ( \30384 , \28133 , \28135 );
or \U$30042 ( \30385 , \30380 , \30383 , \30384 );
xor \U$30043 ( \30386 , \30377 , \30385 );
xor \U$30044 ( \30387 , \27942 , \27944 );
xor \U$30045 ( \30388 , \30387 , \27955 );
xor \U$30046 ( \30389 , \30386 , \30388 );
xor \U$30047 ( \30390 , \30376 , \30389 );
and \U$30048 ( \30391 , \30374 , \30390 );
and \U$30049 ( \30392 , \30376 , \30389 );
nor \U$30050 ( \30393 , \30391 , \30392 );
xnor \U$30051 ( \30394 , \27768 , \27958 );
not \U$30052 ( \30395 , \30394 );
not \U$30053 ( \30396 , \27771 );
and \U$30054 ( \30397 , \30395 , \30396 );
and \U$30055 ( \30398 , \30394 , \27771 );
nor \U$30056 ( \30399 , \30397 , \30398 );
xor \U$30057 ( \30400 , \30377 , \30385 );
and \U$30058 ( \30401 , \30400 , \30388 );
and \U$30059 ( \30402 , \30377 , \30385 );
nor \U$30060 ( \30403 , \30401 , \30402 );
xnor \U$30061 ( \30404 , \30399 , \30403 );
or \U$30062 ( \30405 , \30393 , \30404 );
or \U$30063 ( \30406 , \30403 , \30399 );
nand \U$30064 ( \30407 , \30405 , \30406 );
and \U$30065 ( \30408 , \27962 , \30407 );
nor \U$30066 ( \30409 , \27961 , \30408 );
xor \U$30067 ( \30410 , \27589 , \27591 );
and \U$30068 ( \30411 , \30410 , \27762 );
and \U$30069 ( \30412 , \27589 , \27591 );
nor \U$30070 ( \30413 , \30411 , \30412 );
not \U$30071 ( \30414 , \27368 );
not \U$30072 ( \30415 , \27580 );
not \U$30073 ( \30416 , \27382 );
or \U$30074 ( \30417 , \30415 , \30416 );
or \U$30075 ( \30418 , \27382 , \27580 );
nand \U$30076 ( \30419 , \30417 , \30418 );
not \U$30077 ( \30420 , \30419 );
and \U$30078 ( \30421 , \30414 , \30420 );
and \U$30079 ( \30422 , \27368 , \30419 );
nor \U$30080 ( \30423 , \30421 , \30422 );
xnor \U$30081 ( \30424 , \30413 , \30423 );
or \U$30082 ( \30425 , \30409 , \30424 );
or \U$30083 ( \30426 , \30413 , \30423 );
nand \U$30084 ( \30427 , \30425 , \30426 );
and \U$30085 ( \30428 , \27584 , \30427 );
nor \U$30086 ( \30429 , \27583 , \30428 );
or \U$30087 ( \30430 , \27360 , \30429 );
nand \U$30088 ( \30431 , \27359 , \30430 );
or \U$30089 ( \30432 , \27174 , \26546 );
not \U$30090 ( \30433 , \26546 );
not \U$30091 ( \30434 , \27174 );
or \U$30092 ( \30435 , \30433 , \30434 );
nand \U$30093 ( \30436 , \30435 , \26939 );
nand \U$30094 ( \30437 , \30432 , \30436 );
xor \U$30095 ( \30438 , \26980 , \26984 );
and \U$30096 ( \30439 , \30438 , \26989 );
and \U$30097 ( \30440 , \26980 , \26984 );
nor \U$30098 ( \30441 , \30439 , \30440 );
xor \U$30099 ( \30442 , \27085 , \27089 );
and \U$30100 ( \30443 , \30442 , \27094 );
and \U$30101 ( \30444 , \27085 , \27089 );
nor \U$30102 ( \30445 , \30443 , \30444 );
xor \U$30103 ( \30446 , \30441 , \30445 );
not \U$30104 ( \30447 , \27077 );
not \U$30105 ( \30448 , \27032 );
or \U$30106 ( \30449 , \30447 , \30448 );
or \U$30107 ( \30450 , \27032 , \27077 );
nand \U$30108 ( \30451 , \30450 , \27055 );
nand \U$30109 ( \30452 , \30449 , \30451 );
xor \U$30110 ( \30453 , \30446 , \30452 );
not \U$30111 ( \30454 , \30453 );
xor \U$30112 ( \30455 , \26994 , \27002 );
and \U$30113 ( \30456 , \30455 , \27007 );
and \U$30114 ( \30457 , \26994 , \27002 );
nor \U$30115 ( \30458 , \30456 , \30457 );
not \U$30116 ( \30459 , \30458 );
xor \U$30117 ( \30460 , \27081 , \27095 );
and \U$30118 ( \30461 , \30460 , \27168 );
and \U$30119 ( \30462 , \27081 , \27095 );
or \U$30120 ( \30463 , \30461 , \30462 );
not \U$30121 ( \30464 , \30463 );
or \U$30122 ( \30465 , \30459 , \30464 );
or \U$30123 ( \30466 , \30463 , \30458 );
nand \U$30124 ( \30467 , \30465 , \30466 );
not \U$30125 ( \30468 , \30467 );
xor \U$30126 ( \30469 , \27039 , \27046 );
and \U$30127 ( \30470 , \30469 , \27054 );
and \U$30128 ( \30471 , \27039 , \27046 );
or \U$30129 ( \30472 , \30470 , \30471 );
not \U$30130 ( \30473 , \30472 );
xor \U$30131 ( \30474 , \27016 , \27023 );
and \U$30132 ( \30475 , \30474 , \27031 );
and \U$30133 ( \30476 , \27016 , \27023 );
nor \U$30134 ( \30477 , \30475 , \30476 );
not \U$30135 ( \30478 , \30477 );
or \U$30136 ( \30479 , \30473 , \30478 );
or \U$30137 ( \30480 , \30477 , \30472 );
nand \U$30138 ( \30481 , \30479 , \30480 );
not \U$30139 ( \30482 , \30481 );
not \U$30140 ( \30483 , \27064 );
nand \U$30141 ( \30484 , \30483 , \27073 );
not \U$30142 ( \30485 , \30484 );
and \U$30143 ( \30486 , \30482 , \30485 );
and \U$30144 ( \30487 , \30481 , \30484 );
nor \U$30145 ( \30488 , \30486 , \30487 );
xor \U$30146 ( \30489 , \27126 , \27134 );
and \U$30147 ( \30490 , \30489 , \27142 );
and \U$30148 ( \30491 , \27126 , \27134 );
or \U$30149 ( \30492 , \30490 , \30491 );
xor \U$30150 ( \30493 , \27103 , \27110 );
and \U$30151 ( \30494 , \30493 , \27118 );
and \U$30152 ( \30495 , \27103 , \27110 );
or \U$30153 ( \30496 , \30494 , \30495 );
xor \U$30154 ( \30497 , \30492 , \30496 );
xor \U$30155 ( \30498 , \27151 , \27158 );
and \U$30156 ( \30499 , \30498 , \27166 );
and \U$30157 ( \30500 , \27151 , \27158 );
or \U$30158 ( \30501 , \30499 , \30500 );
xor \U$30159 ( \30502 , \30497 , \30501 );
xor \U$30160 ( \30503 , \30488 , \30502 );
not \U$30161 ( \30504 , \3412 );
nand \U$30162 ( \30505 , RI9870420_85, \3681 );
not \U$30163 ( \30506 , \30505 );
and \U$30164 ( \30507 , \30504 , \30506 );
and \U$30165 ( \30508 , \3412 , \30505 );
nor \U$30166 ( \30509 , \30507 , \30508 );
not \U$30167 ( \30510 , \30509 );
and \U$30168 ( \30511 , \7079 , RI986fca0_69);
and \U$30169 ( \30512 , RI986ff70_75, \7077 );
nor \U$30170 ( \30513 , \30511 , \30512 );
and \U$30171 ( \30514 , \30513 , \6710 );
not \U$30172 ( \30515 , \30513 );
and \U$30173 ( \30516 , \30515 , \6709 );
nor \U$30174 ( \30517 , \30514 , \30516 );
and \U$30175 ( \30518 , \5881 , RI98707e0_93);
and \U$30176 ( \30519 , RI986fac0_65, \5879 );
nor \U$30177 ( \30520 , \30518 , \30519 );
and \U$30178 ( \30521 , \30520 , \5594 );
not \U$30179 ( \30522 , \30520 );
and \U$30180 ( \30523 , \30522 , \5885 );
nor \U$30181 ( \30524 , \30521 , \30523 );
xor \U$30182 ( \30525 , \30517 , \30524 );
and \U$30183 ( \30526 , \6453 , RI986fbb0_67);
and \U$30184 ( \30527 , RI986fd90_71, \6451 );
nor \U$30185 ( \30528 , \30526 , \30527 );
and \U$30186 ( \30529 , \30528 , \6190 );
not \U$30187 ( \30530 , \30528 );
and \U$30188 ( \30531 , \30530 , \6180 );
nor \U$30189 ( \30532 , \30529 , \30531 );
xor \U$30190 ( \30533 , \30525 , \30532 );
not \U$30191 ( \30534 , \30533 );
or \U$30192 ( \30535 , \30510 , \30534 );
or \U$30193 ( \30536 , \30533 , \30509 );
nand \U$30194 ( \30537 , \30535 , \30536 );
not \U$30195 ( \30538 , \30537 );
and \U$30196 ( \30539 , \4710 , RI9870240_81);
and \U$30197 ( \30540 , RI98706f0_91, \4708 );
nor \U$30198 ( \30541 , \30539 , \30540 );
not \U$30199 ( \30542 , \30541 );
not \U$30200 ( \30543 , \4519 );
and \U$30201 ( \30544 , \30542 , \30543 );
and \U$30202 ( \30545 , \30541 , \4521 );
nor \U$30203 ( \30546 , \30544 , \30545 );
and \U$30204 ( \30547 , \4203 , RI9870510_87);
and \U$30205 ( \30548 , RI9870330_83, \4201 );
nor \U$30206 ( \30549 , \30547 , \30548 );
and \U$30207 ( \30550 , \30549 , \3923 );
not \U$30208 ( \30551 , \30549 );
and \U$30209 ( \30552 , \30551 , \4207 );
nor \U$30210 ( \30553 , \30550 , \30552 );
xor \U$30211 ( \30554 , \30546 , \30553 );
and \U$30212 ( \30555 , \5318 , RI9870600_89);
and \U$30213 ( \30556 , RI98708d0_95, \5316 );
nor \U$30214 ( \30557 , \30555 , \30556 );
and \U$30215 ( \30558 , \30557 , \5322 );
not \U$30216 ( \30559 , \30557 );
and \U$30217 ( \30560 , \30559 , \5052 );
nor \U$30218 ( \30561 , \30558 , \30560 );
xor \U$30219 ( \30562 , \30554 , \30561 );
not \U$30220 ( \30563 , \30562 );
and \U$30221 ( \30564 , \30538 , \30563 );
and \U$30222 ( \30565 , \30537 , \30562 );
nor \U$30223 ( \30566 , \30564 , \30565 );
xor \U$30224 ( \30567 , \30503 , \30566 );
not \U$30225 ( \30568 , \30567 );
and \U$30226 ( \30569 , \30468 , \30568 );
and \U$30227 ( \30570 , \30467 , \30567 );
nor \U$30228 ( \30571 , \30569 , \30570 );
not \U$30229 ( \30572 , \30571 );
or \U$30230 ( \30573 , \30454 , \30572 );
or \U$30231 ( \30574 , \30571 , \30453 );
nand \U$30232 ( \30575 , \30573 , \30574 );
or \U$30233 ( \30576 , \27170 , \26971 );
not \U$30234 ( \30577 , \26971 );
not \U$30235 ( \30578 , \27170 );
or \U$30236 ( \30579 , \30577 , \30578 );
nand \U$30237 ( \30580 , \30579 , \26964 );
nand \U$30238 ( \30581 , \30576 , \30580 );
xor \U$30239 ( \30582 , \30575 , \30581 );
not \U$30240 ( \30583 , \26217 );
or \U$30241 ( \30584 , \30583 , \26542 );
and \U$30242 ( \30585 , \30583 , \26542 );
nor \U$30243 ( \30586 , \30585 , \26442 );
not \U$30244 ( \30587 , \30586 );
nand \U$30245 ( \30588 , \30584 , \30587 );
xor \U$30246 ( \30589 , \27119 , \27143 );
and \U$30247 ( \30590 , \30589 , \27167 );
and \U$30248 ( \30591 , \27119 , \27143 );
nor \U$30249 ( \30592 , \30590 , \30591 );
not \U$30250 ( \30593 , RI9873558_190);
and \U$30251 ( \30594 , \15780 , RI986e9e0_29);
and \U$30252 ( \30595 , RI9873648_192, RI986e8f0_27);
nor \U$30253 ( \30596 , \30594 , \30595 );
not \U$30254 ( \30597 , \30596 );
or \U$30255 ( \30598 , \30593 , \30597 );
or \U$30256 ( \30599 , \30596 , RI9873558_190);
nand \U$30257 ( \30600 , \30598 , \30599 );
xor \U$30258 ( \30601 , \30600 , \3918 );
and \U$30259 ( \30602 , \14937 , RI98715f0_123);
and \U$30260 ( \30603 , RI986ead0_31, \14935 );
nor \U$30261 ( \30604 , \30602 , \30603 );
and \U$30262 ( \30605 , \30604 , \14539 );
not \U$30263 ( \30606 , \30604 );
and \U$30264 ( \30607 , \30606 , \14538 );
nor \U$30265 ( \30608 , \30605 , \30607 );
xor \U$30266 ( \30609 , \30601 , \30608 );
xor \U$30267 ( \30610 , \30592 , \30609 );
and \U$30268 ( \30611 , \7729 , RI986fe80_73);
and \U$30269 ( \30612 , RI9870060_77, \7727 );
nor \U$30270 ( \30613 , \30611 , \30612 );
and \U$30271 ( \30614 , \30613 , \7733 );
not \U$30272 ( \30615 , \30613 );
and \U$30273 ( \30616 , \30615 , \7480 );
nor \U$30274 ( \30617 , \30614 , \30616 );
not \U$30275 ( \30618 , \30617 );
and \U$30276 ( \30619 , \8486 , RI9870150_79);
and \U$30277 ( \30620 , RI9870f60_109, \8484 );
nor \U$30278 ( \30621 , \30619 , \30620 );
and \U$30279 ( \30622 , \30621 , \8051 );
not \U$30280 ( \30623 , \30621 );
and \U$30281 ( \30624 , \30623 , \8050 );
nor \U$30282 ( \30625 , \30622 , \30624 );
and \U$30283 ( \30626 , \9237 , RI9870ab0_99);
and \U$30284 ( \30627 , RI9870d80_105, \9235 );
nor \U$30285 ( \30628 , \30626 , \30627 );
and \U$30286 ( \30629 , \30628 , \8836 );
not \U$30287 ( \30630 , \30628 );
and \U$30288 ( \30631 , \30630 , \9241 );
nor \U$30289 ( \30632 , \30629 , \30631 );
xor \U$30290 ( \30633 , \30625 , \30632 );
not \U$30291 ( \30634 , \30633 );
or \U$30292 ( \30635 , \30618 , \30634 );
or \U$30293 ( \30636 , \30633 , \30617 );
nand \U$30294 ( \30637 , \30635 , \30636 );
and \U$30295 ( \30638 , \11696 , RI9870c90_103);
and \U$30296 ( \30639 , RI9871230_115, \11694 );
nor \U$30297 ( \30640 , \30638 , \30639 );
and \U$30298 ( \30641 , \30640 , \10965 );
not \U$30299 ( \30642 , \30640 );
and \U$30300 ( \30643 , \30642 , \11702 );
nor \U$30301 ( \30644 , \30641 , \30643 );
and \U$30302 ( \30645 , \9505 , RI98709c0_97);
and \U$30303 ( \30646 , RI9870e70_107, \9503 );
nor \U$30304 ( \30647 , \30645 , \30646 );
and \U$30305 ( \30648 , \30647 , \9510 );
not \U$30306 ( \30649 , \30647 );
and \U$30307 ( \30650 , \30649 , \9513 );
nor \U$30308 ( \30651 , \30648 , \30650 );
xor \U$30309 ( \30652 , \30644 , \30651 );
and \U$30310 ( \30653 , \10424 , RI9870ba0_101);
and \U$30311 ( \30654 , RI9871050_111, \10422 );
nor \U$30312 ( \30655 , \30653 , \30654 );
and \U$30313 ( \30656 , \30655 , \9840 );
not \U$30314 ( \30657 , \30655 );
and \U$30315 ( \30658 , \30657 , \10428 );
nor \U$30316 ( \30659 , \30656 , \30658 );
xor \U$30317 ( \30660 , \30652 , \30659 );
xor \U$30318 ( \30661 , \30637 , \30660 );
and \U$30319 ( \30662 , \12293 , RI9871140_113);
and \U$30320 ( \30663 , RI9871320_117, \12291 );
nor \U$30321 ( \30664 , \30662 , \30663 );
and \U$30322 ( \30665 , \30664 , \11687 );
not \U$30323 ( \30666 , \30664 );
and \U$30324 ( \30667 , \30666 , \11686 );
nor \U$30325 ( \30668 , \30665 , \30667 );
and \U$30326 ( \30669 , \13045 , RI9871410_119);
and \U$30327 ( \30670 , RI98716e0_125, \13043 );
nor \U$30328 ( \30671 , \30669 , \30670 );
and \U$30329 ( \30672 , \30671 , \13047 );
not \U$30330 ( \30673 , \30671 );
and \U$30331 ( \30674 , \30673 , \12619 );
nor \U$30332 ( \30675 , \30672 , \30674 );
xor \U$30333 ( \30676 , \30668 , \30675 );
and \U$30334 ( \30677 , \13882 , RI98717d0_127);
and \U$30335 ( \30678 , RI9871500_121, \13880 );
nor \U$30336 ( \30679 , \30677 , \30678 );
and \U$30337 ( \30680 , \30679 , \13358 );
not \U$30338 ( \30681 , \30679 );
and \U$30339 ( \30682 , \30681 , \13359 );
nor \U$30340 ( \30683 , \30680 , \30682 );
xor \U$30341 ( \30684 , \30676 , \30683 );
xor \U$30342 ( \30685 , \30661 , \30684 );
xor \U$30343 ( \30686 , \30610 , \30685 );
xor \U$30344 ( \30687 , \30588 , \30686 );
xor \U$30345 ( \30688 , \26990 , \27008 );
and \U$30346 ( \30689 , \30688 , \27169 );
and \U$30347 ( \30690 , \26990 , \27008 );
nor \U$30348 ( \30691 , \30689 , \30690 );
xor \U$30349 ( \30692 , \30687 , \30691 );
xor \U$30350 ( \30693 , \30582 , \30692 );
xor \U$30351 ( \30694 , \30437 , \30693 );
and \U$30352 ( \30695 , \30431 , \30694 );
and \U$30353 ( \30696 , \30437 , \30693 );
nor \U$30354 ( \30697 , \30695 , \30696 );
xor \U$30355 ( \30698 , \30588 , \30686 );
and \U$30356 ( \30699 , \30698 , \30691 );
and \U$30357 ( \30700 , \30588 , \30686 );
or \U$30358 ( \30701 , \30699 , \30700 );
not \U$30359 ( \30702 , \30701 );
not \U$30360 ( \30703 , \30571 );
nand \U$30361 ( \30704 , \30703 , \30453 );
not \U$30362 ( \30705 , \30704 );
and \U$30363 ( \30706 , \30702 , \30705 );
and \U$30364 ( \30707 , \30701 , \30704 );
nor \U$30365 ( \30708 , \30706 , \30707 );
not \U$30366 ( \30709 , \30708 );
xor \U$30367 ( \30710 , \30488 , \30502 );
and \U$30368 ( \30711 , \30710 , \30566 );
and \U$30369 ( \30712 , \30488 , \30502 );
nor \U$30370 ( \30713 , \30711 , \30712 );
xor \U$30371 ( \30714 , \30441 , \30445 );
and \U$30372 ( \30715 , \30714 , \30452 );
and \U$30373 ( \30716 , \30441 , \30445 );
or \U$30374 ( \30717 , \30715 , \30716 );
xor \U$30375 ( \30718 , \30713 , \30717 );
xor \U$30376 ( \30719 , \30592 , \30609 );
and \U$30377 ( \30720 , \30719 , \30685 );
and \U$30378 ( \30721 , \30592 , \30609 );
or \U$30379 ( \30722 , \30720 , \30721 );
xor \U$30380 ( \30723 , \30718 , \30722 );
or \U$30381 ( \30724 , \30567 , \30463 );
not \U$30382 ( \30725 , \30463 );
not \U$30383 ( \30726 , \30567 );
or \U$30384 ( \30727 , \30725 , \30726 );
nand \U$30385 ( \30728 , \30727 , \30458 );
nand \U$30386 ( \30729 , \30724 , \30728 );
xor \U$30387 ( \30730 , \30492 , \30496 );
and \U$30388 ( \30731 , \30730 , \30501 );
and \U$30389 ( \30732 , \30492 , \30496 );
nor \U$30390 ( \30733 , \30731 , \30732 );
or \U$30391 ( \30734 , \30477 , \30484 );
not \U$30392 ( \30735 , \30484 );
not \U$30393 ( \30736 , \30477 );
or \U$30394 ( \30737 , \30735 , \30736 );
nand \U$30395 ( \30738 , \30737 , \30472 );
nand \U$30396 ( \30739 , \30734 , \30738 );
xor \U$30397 ( \30740 , \30733 , \30739 );
or \U$30398 ( \30741 , \30562 , \30509 );
not \U$30399 ( \30742 , \30509 );
not \U$30400 ( \30743 , \30562 );
or \U$30401 ( \30744 , \30742 , \30743 );
nand \U$30402 ( \30745 , \30744 , \30533 );
nand \U$30403 ( \30746 , \30741 , \30745 );
xor \U$30404 ( \30747 , \30740 , \30746 );
xor \U$30405 ( \30748 , \30668 , \30675 );
and \U$30406 ( \30749 , \30748 , \30683 );
and \U$30407 ( \30750 , \30668 , \30675 );
or \U$30408 ( \30751 , \30749 , \30750 );
xor \U$30409 ( \30752 , \30600 , \3918 );
and \U$30410 ( \30753 , \30752 , \30608 );
and \U$30411 ( \30754 , \30600 , \3918 );
or \U$30412 ( \30755 , \30753 , \30754 );
xor \U$30413 ( \30756 , \30751 , \30755 );
xor \U$30414 ( \30757 , \30644 , \30651 );
and \U$30415 ( \30758 , \30757 , \30659 );
and \U$30416 ( \30759 , \30644 , \30651 );
or \U$30417 ( \30760 , \30758 , \30759 );
xor \U$30418 ( \30761 , \30756 , \30760 );
not \U$30419 ( \30762 , \30761 );
xor \U$30420 ( \30763 , \30517 , \30524 );
and \U$30421 ( \30764 , \30763 , \30532 );
and \U$30422 ( \30765 , \30517 , \30524 );
or \U$30423 ( \30766 , \30764 , \30765 );
not \U$30424 ( \30767 , \30766 );
not \U$30425 ( \30768 , \30617 );
not \U$30426 ( \30769 , \30625 );
and \U$30427 ( \30770 , \30768 , \30769 );
and \U$30428 ( \30771 , \30625 , \30617 );
nor \U$30429 ( \30772 , \30771 , \30632 );
nor \U$30430 ( \30773 , \30770 , \30772 );
not \U$30431 ( \30774 , \30773 );
or \U$30432 ( \30775 , \30767 , \30774 );
or \U$30433 ( \30776 , \30773 , \30766 );
nand \U$30434 ( \30777 , \30775 , \30776 );
not \U$30435 ( \30778 , \30777 );
xor \U$30436 ( \30779 , \30546 , \30553 );
and \U$30437 ( \30780 , \30779 , \30561 );
and \U$30438 ( \30781 , \30546 , \30553 );
or \U$30439 ( \30782 , \30780 , \30781 );
not \U$30440 ( \30783 , \30782 );
and \U$30441 ( \30784 , \30778 , \30783 );
and \U$30442 ( \30785 , \30777 , \30782 );
nor \U$30443 ( \30786 , \30784 , \30785 );
not \U$30444 ( \30787 , \30786 );
or \U$30445 ( \30788 , \30762 , \30787 );
or \U$30446 ( \30789 , \30786 , \30761 );
nand \U$30447 ( \30790 , \30788 , \30789 );
xor \U$30448 ( \30791 , \30747 , \30790 );
and \U$30449 ( \30792 , \6453 , RI986fd90_71);
and \U$30450 ( \30793 , RI986fca0_69, \6451 );
nor \U$30451 ( \30794 , \30792 , \30793 );
and \U$30452 ( \30795 , \30794 , \6190 );
not \U$30453 ( \30796 , \30794 );
and \U$30454 ( \30797 , \30796 , \6705 );
nor \U$30455 ( \30798 , \30795 , \30797 );
and \U$30456 ( \30799 , \5318 , RI98708d0_95);
and \U$30457 ( \30800 , RI98707e0_93, \5316 );
nor \U$30458 ( \30801 , \30799 , \30800 );
and \U$30459 ( \30802 , \30801 , \5052 );
not \U$30460 ( \30803 , \30801 );
and \U$30461 ( \30804 , \30803 , \5322 );
nor \U$30462 ( \30805 , \30802 , \30804 );
xor \U$30463 ( \30806 , \30798 , \30805 );
and \U$30464 ( \30807 , \5881 , RI986fac0_65);
and \U$30465 ( \30808 , RI986fbb0_67, \5879 );
nor \U$30466 ( \30809 , \30807 , \30808 );
and \U$30467 ( \30810 , \30809 , \5594 );
not \U$30468 ( \30811 , \30809 );
and \U$30469 ( \30812 , \30811 , \5885 );
nor \U$30470 ( \30813 , \30810 , \30812 );
xor \U$30471 ( \30814 , \30806 , \30813 );
and \U$30472 ( \30815 , \4203 , RI9870330_83);
and \U$30473 ( \30816 , RI9870240_81, \4201 );
nor \U$30474 ( \30817 , \30815 , \30816 );
and \U$30475 ( \30818 , \30817 , \4207 );
not \U$30476 ( \30819 , \30817 );
and \U$30477 ( \30820 , \30819 , \3922 );
nor \U$30478 ( \30821 , \30818 , \30820 );
not \U$30479 ( \30822 , \3412 );
and \U$30480 ( \30823 , \3683 , RI9870420_85);
and \U$30481 ( \30824 , RI9870510_87, \3681 );
nor \U$30482 ( \30825 , \30823 , \30824 );
not \U$30483 ( \30826 , \30825 );
or \U$30484 ( \30827 , \30822 , \30826 );
or \U$30485 ( \30828 , \30825 , \3412 );
nand \U$30486 ( \30829 , \30827 , \30828 );
xor \U$30487 ( \30830 , \30821 , \30829 );
not \U$30488 ( \30831 , \4519 );
and \U$30489 ( \30832 , \4710 , RI98706f0_91);
and \U$30490 ( \30833 , RI9870600_89, \4708 );
nor \U$30491 ( \30834 , \30832 , \30833 );
not \U$30492 ( \30835 , \30834 );
or \U$30493 ( \30836 , \30831 , \30835 );
or \U$30494 ( \30837 , \30834 , \4521 );
nand \U$30495 ( \30838 , \30836 , \30837 );
xor \U$30496 ( \30839 , \30830 , \30838 );
xor \U$30497 ( \30840 , \30814 , \30839 );
and \U$30498 ( \30841 , \8486 , RI9870f60_109);
and \U$30499 ( \30842 , RI9870ab0_99, \8484 );
nor \U$30500 ( \30843 , \30841 , \30842 );
and \U$30501 ( \30844 , \30843 , \8050 );
not \U$30502 ( \30845 , \30843 );
and \U$30503 ( \30846 , \30845 , \8051 );
nor \U$30504 ( \30847 , \30844 , \30846 );
and \U$30505 ( \30848 , \7079 , RI986ff70_75);
and \U$30506 ( \30849 , RI986fe80_73, \7077 );
nor \U$30507 ( \30850 , \30848 , \30849 );
and \U$30508 ( \30851 , \30850 , \6710 );
not \U$30509 ( \30852 , \30850 );
and \U$30510 ( \30853 , \30852 , \6709 );
nor \U$30511 ( \30854 , \30851 , \30853 );
xor \U$30512 ( \30855 , \30847 , \30854 );
and \U$30513 ( \30856 , \7729 , RI9870060_77);
and \U$30514 ( \30857 , RI9870150_79, \7727 );
nor \U$30515 ( \30858 , \30856 , \30857 );
and \U$30516 ( \30859 , \30858 , \7480 );
not \U$30517 ( \30860 , \30858 );
and \U$30518 ( \30861 , \30860 , \7733 );
nor \U$30519 ( \30862 , \30859 , \30861 );
xor \U$30520 ( \30863 , \30855 , \30862 );
xor \U$30521 ( \30864 , \30840 , \30863 );
xor \U$30522 ( \30865 , \30637 , \30660 );
and \U$30523 ( \30866 , \30865 , \30684 );
and \U$30524 ( \30867 , \30637 , \30660 );
or \U$30525 ( \30868 , \30866 , \30867 );
and \U$30526 ( \30869 , \9505 , RI9870e70_107);
and \U$30527 ( \30870 , RI9870ba0_101, \9503 );
nor \U$30528 ( \30871 , \30869 , \30870 );
and \U$30529 ( \30872 , \30871 , \9510 );
not \U$30530 ( \30873 , \30871 );
and \U$30531 ( \30874 , \30873 , \9513 );
nor \U$30532 ( \30875 , \30872 , \30874 );
and \U$30533 ( \30876 , \9237 , RI9870d80_105);
and \U$30534 ( \30877 , RI98709c0_97, \9235 );
nor \U$30535 ( \30878 , \30876 , \30877 );
and \U$30536 ( \30879 , \30878 , \9241 );
not \U$30537 ( \30880 , \30878 );
and \U$30538 ( \30881 , \30880 , \8836 );
nor \U$30539 ( \30882 , \30879 , \30881 );
xor \U$30540 ( \30883 , \30875 , \30882 );
and \U$30541 ( \30884 , \10424 , RI9871050_111);
and \U$30542 ( \30885 , RI9870c90_103, \10422 );
nor \U$30543 ( \30886 , \30884 , \30885 );
and \U$30544 ( \30887 , \30886 , \9840 );
not \U$30545 ( \30888 , \30886 );
and \U$30546 ( \30889 , \30888 , \10428 );
nor \U$30547 ( \30890 , \30887 , \30889 );
xor \U$30548 ( \30891 , \30883 , \30890 );
and \U$30549 ( \30892 , \14937 , RI986ead0_31);
and \U$30550 ( \30893 , RI986e9e0_29, \14935 );
nor \U$30551 ( \30894 , \30892 , \30893 );
and \U$30552 ( \30895 , \30894 , \14539 );
not \U$30553 ( \30896 , \30894 );
and \U$30554 ( \30897 , \30896 , \14538 );
nor \U$30555 ( \30898 , \30895 , \30897 );
not \U$30556 ( \30899 , RI9873558_190);
and \U$30557 ( \30900 , \15780 , RI986e8f0_27);
and \U$30558 ( \30901 , RI9873648_192, RI986e800_25);
nor \U$30559 ( \30902 , \30900 , \30901 );
not \U$30560 ( \30903 , \30902 );
or \U$30561 ( \30904 , \30899 , \30903 );
or \U$30562 ( \30905 , \30902 , RI9873558_190);
nand \U$30563 ( \30906 , \30904 , \30905 );
xor \U$30564 ( \30907 , \30898 , \30906 );
and \U$30565 ( \30908 , \13882 , RI9871500_121);
and \U$30566 ( \30909 , RI98715f0_123, \13880 );
nor \U$30567 ( \30910 , \30908 , \30909 );
and \U$30568 ( \30911 , \30910 , \13358 );
not \U$30569 ( \30912 , \30910 );
and \U$30570 ( \30913 , \30912 , \13359 );
nor \U$30571 ( \30914 , \30911 , \30913 );
xor \U$30572 ( \30915 , \30907 , \30914 );
and \U$30573 ( \30916 , \12293 , RI9871320_117);
and \U$30574 ( \30917 , RI9871410_119, \12291 );
nor \U$30575 ( \30918 , \30916 , \30917 );
and \U$30576 ( \30919 , \30918 , \11687 );
not \U$30577 ( \30920 , \30918 );
and \U$30578 ( \30921 , \30920 , \11686 );
nor \U$30579 ( \30922 , \30919 , \30921 );
and \U$30580 ( \30923 , \11696 , RI9871230_115);
and \U$30581 ( \30924 , RI9871140_113, \11694 );
nor \U$30582 ( \30925 , \30923 , \30924 );
and \U$30583 ( \30926 , \30925 , \10965 );
not \U$30584 ( \30927 , \30925 );
and \U$30585 ( \30928 , \30927 , \11702 );
nor \U$30586 ( \30929 , \30926 , \30928 );
xor \U$30587 ( \30930 , \30922 , \30929 );
and \U$30588 ( \30931 , \13045 , RI98716e0_125);
and \U$30589 ( \30932 , RI98717d0_127, \13043 );
nor \U$30590 ( \30933 , \30931 , \30932 );
and \U$30591 ( \30934 , \30933 , \13047 );
not \U$30592 ( \30935 , \30933 );
and \U$30593 ( \30936 , \30935 , \12619 );
nor \U$30594 ( \30937 , \30934 , \30936 );
xor \U$30595 ( \30938 , \30930 , \30937 );
xor \U$30596 ( \30939 , \30915 , \30938 );
xor \U$30597 ( \30940 , \30891 , \30939 );
xor \U$30598 ( \30941 , \30868 , \30940 );
xor \U$30599 ( \30942 , \30864 , \30941 );
xor \U$30600 ( \30943 , \30791 , \30942 );
xor \U$30601 ( \30944 , \30729 , \30943 );
xor \U$30602 ( \30945 , \30723 , \30944 );
not \U$30603 ( \30946 , \30945 );
and \U$30604 ( \30947 , \30709 , \30946 );
and \U$30605 ( \30948 , \30708 , \30945 );
nor \U$30606 ( \30949 , \30947 , \30948 );
xor \U$30607 ( \30950 , \30575 , \30581 );
and \U$30608 ( \30951 , \30950 , \30692 );
and \U$30609 ( \30952 , \30575 , \30581 );
nor \U$30610 ( \30953 , \30951 , \30952 );
xnor \U$30611 ( \30954 , \30949 , \30953 );
or \U$30612 ( \30955 , \30697 , \30954 );
or \U$30613 ( \30956 , \30949 , \30953 );
nand \U$30614 ( \30957 , \30955 , \30956 );
not \U$30615 ( \30958 , \30945 );
or \U$30616 ( \30959 , \30958 , \30704 );
not \U$30617 ( \30960 , \30704 );
not \U$30618 ( \30961 , \30958 );
or \U$30619 ( \30962 , \30960 , \30961 );
nand \U$30620 ( \30963 , \30962 , \30701 );
nand \U$30621 ( \30964 , \30959 , \30963 );
xor \U$30622 ( \30965 , \30713 , \30717 );
and \U$30623 ( \30966 , \30965 , \30722 );
and \U$30624 ( \30967 , \30713 , \30717 );
or \U$30625 ( \30968 , \30966 , \30967 );
xor \U$30626 ( \30969 , \30747 , \30790 );
and \U$30627 ( \30970 , \30969 , \30942 );
and \U$30628 ( \30971 , \30747 , \30790 );
or \U$30629 ( \30972 , \30970 , \30971 );
xor \U$30630 ( \30973 , \30968 , \30972 );
xor \U$30631 ( \30974 , \30798 , \30805 );
and \U$30632 ( \30975 , \30974 , \30813 );
and \U$30633 ( \30976 , \30798 , \30805 );
or \U$30634 ( \30977 , \30975 , \30976 );
xor \U$30635 ( \30978 , \30821 , \30829 );
and \U$30636 ( \30979 , \30978 , \30838 );
and \U$30637 ( \30980 , \30821 , \30829 );
or \U$30638 ( \30981 , \30979 , \30980 );
xor \U$30639 ( \30982 , \30977 , \30981 );
xor \U$30640 ( \30983 , \30847 , \30854 );
and \U$30641 ( \30984 , \30983 , \30862 );
and \U$30642 ( \30985 , \30847 , \30854 );
or \U$30643 ( \30986 , \30984 , \30985 );
xor \U$30644 ( \30987 , \30982 , \30986 );
nand \U$30645 ( \30988 , RI9870420_85, \3252 );
not \U$30646 ( \30989 , \30988 );
not \U$30647 ( \30990 , \2935 );
or \U$30648 ( \30991 , \30989 , \30990 );
or \U$30649 ( \30992 , \2935 , \30988 );
nand \U$30650 ( \30993 , \30991 , \30992 );
not \U$30651 ( \30994 , \3918 );
and \U$30652 ( \30995 , \3683 , RI9870510_87);
and \U$30653 ( \30996 , RI9870330_83, \3681 );
nor \U$30654 ( \30997 , \30995 , \30996 );
not \U$30655 ( \30998 , \30997 );
or \U$30656 ( \30999 , \30994 , \30998 );
or \U$30657 ( \31000 , \30997 , \3918 );
nand \U$30658 ( \31001 , \30999 , \31000 );
xor \U$30659 ( \31002 , \30993 , \31001 );
and \U$30660 ( \31003 , \4203 , RI9870240_81);
and \U$30661 ( \31004 , RI98706f0_91, \4201 );
nor \U$30662 ( \31005 , \31003 , \31004 );
and \U$30663 ( \31006 , \31005 , \3923 );
not \U$30664 ( \31007 , \31005 );
and \U$30665 ( \31008 , \31007 , \4207 );
nor \U$30666 ( \31009 , \31006 , \31008 );
not \U$30667 ( \31010 , \31009 );
and \U$30668 ( \31011 , \4710 , RI9870600_89);
and \U$30669 ( \31012 , RI98708d0_95, \4708 );
nor \U$30670 ( \31013 , \31011 , \31012 );
not \U$30671 ( \31014 , \31013 );
not \U$30672 ( \31015 , \4521 );
and \U$30673 ( \31016 , \31014 , \31015 );
and \U$30674 ( \31017 , \31013 , \4521 );
nor \U$30675 ( \31018 , \31016 , \31017 );
and \U$30676 ( \31019 , \5318 , RI98707e0_93);
and \U$30677 ( \31020 , RI986fac0_65, \5316 );
nor \U$30678 ( \31021 , \31019 , \31020 );
and \U$30679 ( \31022 , \31021 , \5322 );
not \U$30680 ( \31023 , \31021 );
and \U$30681 ( \31024 , \31023 , \5052 );
nor \U$30682 ( \31025 , \31022 , \31024 );
xor \U$30683 ( \31026 , \31018 , \31025 );
not \U$30684 ( \31027 , \31026 );
or \U$30685 ( \31028 , \31010 , \31027 );
or \U$30686 ( \31029 , \31026 , \31009 );
nand \U$30687 ( \31030 , \31028 , \31029 );
xor \U$30688 ( \31031 , \31002 , \31030 );
xor \U$30689 ( \31032 , \30987 , \31031 );
xor \U$30690 ( \31033 , \30922 , \30929 );
and \U$30691 ( \31034 , \31033 , \30937 );
and \U$30692 ( \31035 , \30922 , \30929 );
or \U$30693 ( \31036 , \31034 , \31035 );
xor \U$30694 ( \31037 , \30898 , \30906 );
and \U$30695 ( \31038 , \31037 , \30914 );
and \U$30696 ( \31039 , \30898 , \30906 );
or \U$30697 ( \31040 , \31038 , \31039 );
xor \U$30698 ( \31041 , \31036 , \31040 );
xor \U$30699 ( \31042 , \30875 , \30882 );
and \U$30700 ( \31043 , \31042 , \30890 );
and \U$30701 ( \31044 , \30875 , \30882 );
or \U$30702 ( \31045 , \31043 , \31044 );
xor \U$30703 ( \31046 , \31041 , \31045 );
xor \U$30704 ( \31047 , \31032 , \31046 );
or \U$30705 ( \31048 , \30782 , \30773 );
not \U$30706 ( \31049 , \30782 );
not \U$30707 ( \31050 , \30773 );
or \U$30708 ( \31051 , \31049 , \31050 );
nand \U$30709 ( \31052 , \31051 , \30766 );
nand \U$30710 ( \31053 , \31048 , \31052 );
xor \U$30711 ( \31054 , \30751 , \30755 );
and \U$30712 ( \31055 , \31054 , \30760 );
and \U$30713 ( \31056 , \30751 , \30755 );
or \U$30714 ( \31057 , \31055 , \31056 );
xor \U$30715 ( \31058 , \31053 , \31057 );
xor \U$30716 ( \31059 , \30814 , \30839 );
and \U$30717 ( \31060 , \31059 , \30863 );
and \U$30718 ( \31061 , \30814 , \30839 );
or \U$30719 ( \31062 , \31060 , \31061 );
xor \U$30720 ( \31063 , \31058 , \31062 );
xor \U$30721 ( \31064 , \30875 , \30882 );
xor \U$30722 ( \31065 , \31064 , \30890 );
and \U$30723 ( \31066 , \30915 , \31065 );
xor \U$30724 ( \31067 , \30875 , \30882 );
xor \U$30725 ( \31068 , \31067 , \30890 );
and \U$30726 ( \31069 , \30938 , \31068 );
and \U$30727 ( \31070 , \30915 , \30938 );
or \U$30728 ( \31071 , \31066 , \31069 , \31070 );
and \U$30729 ( \31072 , \13045 , RI98717d0_127);
and \U$30730 ( \31073 , RI9871500_121, \13043 );
nor \U$30731 ( \31074 , \31072 , \31073 );
and \U$30732 ( \31075 , \31074 , \12619 );
not \U$30733 ( \31076 , \31074 );
and \U$30734 ( \31077 , \31076 , \13047 );
nor \U$30735 ( \31078 , \31075 , \31077 );
not \U$30736 ( \31079 , \31078 );
and \U$30737 ( \31080 , \13882 , RI98715f0_123);
and \U$30738 ( \31081 , RI986ead0_31, \13880 );
nor \U$30739 ( \31082 , \31080 , \31081 );
and \U$30740 ( \31083 , \31082 , \13358 );
not \U$30741 ( \31084 , \31082 );
and \U$30742 ( \31085 , \31084 , \13359 );
nor \U$30743 ( \31086 , \31083 , \31085 );
not \U$30744 ( \31087 , \31086 );
or \U$30745 ( \31088 , \31079 , \31087 );
or \U$30746 ( \31089 , \31078 , \31086 );
nand \U$30747 ( \31090 , \31088 , \31089 );
not \U$30748 ( \31091 , \31090 );
and \U$30749 ( \31092 , \12293 , RI9871410_119);
and \U$30750 ( \31093 , RI98716e0_125, \12291 );
nor \U$30751 ( \31094 , \31092 , \31093 );
and \U$30752 ( \31095 , \31094 , \11686 );
not \U$30753 ( \31096 , \31094 );
and \U$30754 ( \31097 , \31096 , \11687 );
nor \U$30755 ( \31098 , \31095 , \31097 );
not \U$30756 ( \31099 , \31098 );
and \U$30757 ( \31100 , \31091 , \31099 );
and \U$30758 ( \31101 , \31090 , \31098 );
nor \U$30759 ( \31102 , \31100 , \31101 );
not \U$30760 ( \31103 , \31102 );
not \U$30761 ( \31104 , RI9873558_190);
and \U$30762 ( \31105 , \15780 , RI986e800_25);
and \U$30763 ( \31106 , RI9873648_192, RI986ee90_39);
nor \U$30764 ( \31107 , \31105 , \31106 );
not \U$30765 ( \31108 , \31107 );
or \U$30766 ( \31109 , \31104 , \31108 );
or \U$30767 ( \31110 , \31107 , RI9873558_190);
nand \U$30768 ( \31111 , \31109 , \31110 );
xor \U$30769 ( \31112 , \31111 , \3406 );
and \U$30770 ( \31113 , \14937 , RI986e9e0_29);
and \U$30771 ( \31114 , RI986e8f0_27, \14935 );
nor \U$30772 ( \31115 , \31113 , \31114 );
and \U$30773 ( \31116 , \31115 , \14539 );
not \U$30774 ( \31117 , \31115 );
and \U$30775 ( \31118 , \31117 , \14538 );
nor \U$30776 ( \31119 , \31116 , \31118 );
xor \U$30777 ( \31120 , \31112 , \31119 );
not \U$30778 ( \31121 , \31120 );
or \U$30779 ( \31122 , \31103 , \31121 );
or \U$30780 ( \31123 , \31120 , \31102 );
nand \U$30781 ( \31124 , \31122 , \31123 );
xor \U$30782 ( \31125 , \31071 , \31124 );
and \U$30783 ( \31126 , \5881 , RI986fbb0_67);
and \U$30784 ( \31127 , RI986fd90_71, \5879 );
nor \U$30785 ( \31128 , \31126 , \31127 );
and \U$30786 ( \31129 , \31128 , \5885 );
not \U$30787 ( \31130 , \31128 );
and \U$30788 ( \31131 , \31130 , \5594 );
nor \U$30789 ( \31132 , \31129 , \31131 );
and \U$30790 ( \31133 , \6453 , RI986fca0_69);
and \U$30791 ( \31134 , RI986ff70_75, \6451 );
nor \U$30792 ( \31135 , \31133 , \31134 );
and \U$30793 ( \31136 , \31135 , \6180 );
not \U$30794 ( \31137 , \31135 );
and \U$30795 ( \31138 , \31137 , \6190 );
nor \U$30796 ( \31139 , \31136 , \31138 );
xor \U$30797 ( \31140 , \31132 , \31139 );
and \U$30798 ( \31141 , \7079 , RI986fe80_73);
and \U$30799 ( \31142 , RI9870060_77, \7077 );
nor \U$30800 ( \31143 , \31141 , \31142 );
and \U$30801 ( \31144 , \31143 , \6709 );
not \U$30802 ( \31145 , \31143 );
and \U$30803 ( \31146 , \31145 , \6710 );
nor \U$30804 ( \31147 , \31144 , \31146 );
xor \U$30805 ( \31148 , \31140 , \31147 );
not \U$30806 ( \31149 , \31148 );
and \U$30807 ( \31150 , \7729 , RI9870150_79);
and \U$30808 ( \31151 , RI9870f60_109, \7727 );
nor \U$30809 ( \31152 , \31150 , \31151 );
and \U$30810 ( \31153 , \31152 , \7733 );
not \U$30811 ( \31154 , \31152 );
and \U$30812 ( \31155 , \31154 , \7480 );
nor \U$30813 ( \31156 , \31153 , \31155 );
and \U$30814 ( \31157 , \8486 , RI9870ab0_99);
and \U$30815 ( \31158 , RI9870d80_105, \8484 );
nor \U$30816 ( \31159 , \31157 , \31158 );
and \U$30817 ( \31160 , \31159 , \8051 );
not \U$30818 ( \31161 , \31159 );
and \U$30819 ( \31162 , \31161 , \8050 );
nor \U$30820 ( \31163 , \31160 , \31162 );
xor \U$30821 ( \31164 , \31156 , \31163 );
and \U$30822 ( \31165 , \9237 , RI98709c0_97);
and \U$30823 ( \31166 , RI9870e70_107, \9235 );
nor \U$30824 ( \31167 , \31165 , \31166 );
and \U$30825 ( \31168 , \31167 , \8836 );
not \U$30826 ( \31169 , \31167 );
and \U$30827 ( \31170 , \31169 , \9241 );
nor \U$30828 ( \31171 , \31168 , \31170 );
xor \U$30829 ( \31172 , \31164 , \31171 );
and \U$30830 ( \31173 , \10424 , RI9870c90_103);
and \U$30831 ( \31174 , RI9871230_115, \10422 );
nor \U$30832 ( \31175 , \31173 , \31174 );
and \U$30833 ( \31176 , \31175 , \10428 );
not \U$30834 ( \31177 , \31175 );
and \U$30835 ( \31178 , \31177 , \9840 );
nor \U$30836 ( \31179 , \31176 , \31178 );
and \U$30837 ( \31180 , \11696 , RI9871140_113);
and \U$30838 ( \31181 , RI9871320_117, \11694 );
nor \U$30839 ( \31182 , \31180 , \31181 );
and \U$30840 ( \31183 , \31182 , \11702 );
not \U$30841 ( \31184 , \31182 );
and \U$30842 ( \31185 , \31184 , \10965 );
nor \U$30843 ( \31186 , \31183 , \31185 );
xor \U$30844 ( \31187 , \31179 , \31186 );
and \U$30845 ( \31188 , \9505 , RI9870ba0_101);
and \U$30846 ( \31189 , RI9871050_111, \9503 );
nor \U$30847 ( \31190 , \31188 , \31189 );
and \U$30848 ( \31191 , \31190 , \9513 );
not \U$30849 ( \31192 , \31190 );
and \U$30850 ( \31193 , \31192 , \9510 );
nor \U$30851 ( \31194 , \31191 , \31193 );
xor \U$30852 ( \31195 , \31187 , \31194 );
xor \U$30853 ( \31196 , \31172 , \31195 );
not \U$30854 ( \31197 , \31196 );
or \U$30855 ( \31198 , \31149 , \31197 );
or \U$30856 ( \31199 , \31196 , \31148 );
nand \U$30857 ( \31200 , \31198 , \31199 );
xor \U$30858 ( \31201 , \31125 , \31200 );
xor \U$30859 ( \31202 , \31063 , \31201 );
xor \U$30860 ( \31203 , \31047 , \31202 );
xor \U$30861 ( \31204 , \30973 , \31203 );
not \U$30862 ( \31205 , \30786 );
nand \U$30863 ( \31206 , \31205 , \30761 );
not \U$30864 ( \31207 , \31206 );
xor \U$30865 ( \31208 , \30733 , \30739 );
and \U$30866 ( \31209 , \31208 , \30746 );
and \U$30867 ( \31210 , \30733 , \30739 );
nor \U$30868 ( \31211 , \31209 , \31210 );
not \U$30869 ( \31212 , \31211 );
xor \U$30870 ( \31213 , \30814 , \30839 );
xor \U$30871 ( \31214 , \31213 , \30863 );
and \U$30872 ( \31215 , \30868 , \31214 );
xor \U$30873 ( \31216 , \30814 , \30839 );
xor \U$30874 ( \31217 , \31216 , \30863 );
and \U$30875 ( \31218 , \30940 , \31217 );
and \U$30876 ( \31219 , \30868 , \30940 );
or \U$30877 ( \31220 , \31215 , \31218 , \31219 );
not \U$30878 ( \31221 , \31220 );
or \U$30879 ( \31222 , \31212 , \31221 );
or \U$30880 ( \31223 , \31220 , \31211 );
nand \U$30881 ( \31224 , \31222 , \31223 );
not \U$30882 ( \31225 , \31224 );
or \U$30883 ( \31226 , \31207 , \31225 );
or \U$30884 ( \31227 , \31224 , \31206 );
nand \U$30885 ( \31228 , \31226 , \31227 );
xor \U$30886 ( \31229 , \31204 , \31228 );
xor \U$30887 ( \31230 , \30713 , \30717 );
xor \U$30888 ( \31231 , \31230 , \30722 );
and \U$30889 ( \31232 , \30729 , \31231 );
xor \U$30890 ( \31233 , \30713 , \30717 );
xor \U$30891 ( \31234 , \31233 , \30722 );
and \U$30892 ( \31235 , \30943 , \31234 );
and \U$30893 ( \31236 , \30729 , \30943 );
or \U$30894 ( \31237 , \31232 , \31235 , \31236 );
xor \U$30895 ( \31238 , \31229 , \31237 );
xor \U$30896 ( \31239 , \30964 , \31238 );
and \U$30897 ( \31240 , \30957 , \31239 );
and \U$30898 ( \31241 , \30964 , \31238 );
nor \U$30899 ( \31242 , \31240 , \31241 );
xor \U$30900 ( \31243 , \31204 , \31228 );
and \U$30901 ( \31244 , \31243 , \31237 );
and \U$30902 ( \31245 , \31204 , \31228 );
nor \U$30903 ( \31246 , \31244 , \31245 );
xor \U$30904 ( \31247 , \30968 , \30972 );
and \U$30905 ( \31248 , \31247 , \31203 );
and \U$30906 ( \31249 , \30968 , \30972 );
or \U$30907 ( \31250 , \31248 , \31249 );
xor \U$30908 ( \31251 , \31036 , \31040 );
and \U$30909 ( \31252 , \31251 , \31045 );
and \U$30910 ( \31253 , \31036 , \31040 );
nor \U$30911 ( \31254 , \31252 , \31253 );
xor \U$30912 ( \31255 , \30993 , \31001 );
and \U$30913 ( \31256 , \31255 , \31030 );
and \U$30914 ( \31257 , \30993 , \31001 );
nor \U$30915 ( \31258 , \31256 , \31257 );
xor \U$30916 ( \31259 , \31254 , \31258 );
xor \U$30917 ( \31260 , \30977 , \30981 );
and \U$30918 ( \31261 , \31260 , \30986 );
and \U$30919 ( \31262 , \30977 , \30981 );
nor \U$30920 ( \31263 , \31261 , \31262 );
xor \U$30921 ( \31264 , \31259 , \31263 );
not \U$30922 ( \31265 , \31264 );
not \U$30923 ( \31266 , \31206 );
and \U$30924 ( \31267 , \31220 , \31266 );
not \U$30925 ( \31268 , \31220 );
not \U$30926 ( \31269 , \31266 );
and \U$30927 ( \31270 , \31268 , \31269 );
nor \U$30928 ( \31271 , \31270 , \31211 );
nor \U$30929 ( \31272 , \31267 , \31271 );
xor \U$30930 ( \31273 , \30987 , \31031 );
xor \U$30931 ( \31274 , \31273 , \31046 );
and \U$30932 ( \31275 , \31063 , \31274 );
xor \U$30933 ( \31276 , \30987 , \31031 );
xor \U$30934 ( \31277 , \31276 , \31046 );
and \U$30935 ( \31278 , \31201 , \31277 );
and \U$30936 ( \31279 , \31063 , \31201 );
or \U$30937 ( \31280 , \31275 , \31278 , \31279 );
not \U$30938 ( \31281 , \31280 );
xor \U$30939 ( \31282 , \31272 , \31281 );
not \U$30940 ( \31283 , \31282 );
or \U$30941 ( \31284 , \31265 , \31283 );
or \U$30942 ( \31285 , \31282 , \31264 );
nand \U$30943 ( \31286 , \31284 , \31285 );
xnor \U$30944 ( \31287 , \31250 , \31286 );
not \U$30945 ( \31288 , \31287 );
xor \U$30946 ( \31289 , \30987 , \31031 );
and \U$30947 ( \31290 , \31289 , \31046 );
and \U$30948 ( \31291 , \30987 , \31031 );
or \U$30949 ( \31292 , \31290 , \31291 );
xor \U$30950 ( \31293 , \31053 , \31057 );
and \U$30951 ( \31294 , \31293 , \31062 );
and \U$30952 ( \31295 , \31053 , \31057 );
or \U$30953 ( \31296 , \31294 , \31295 );
xor \U$30954 ( \31297 , \31292 , \31296 );
xor \U$30955 ( \31298 , \31071 , \31124 );
and \U$30956 ( \31299 , \31298 , \31200 );
and \U$30957 ( \31300 , \31071 , \31124 );
or \U$30958 ( \31301 , \31299 , \31300 );
xor \U$30959 ( \31302 , \31297 , \31301 );
not \U$30960 ( \31303 , \31302 );
or \U$30961 ( \31304 , \31098 , \31078 );
not \U$30962 ( \31305 , \31078 );
not \U$30963 ( \31306 , \31098 );
or \U$30964 ( \31307 , \31305 , \31306 );
nand \U$30965 ( \31308 , \31307 , \31086 );
nand \U$30966 ( \31309 , \31304 , \31308 );
xor \U$30967 ( \31310 , \31179 , \31186 );
and \U$30968 ( \31311 , \31310 , \31194 );
and \U$30969 ( \31312 , \31179 , \31186 );
nor \U$30970 ( \31313 , \31311 , \31312 );
xnor \U$30971 ( \31314 , \31309 , \31313 );
not \U$30972 ( \31315 , \31314 );
xor \U$30973 ( \31316 , \31111 , \3406 );
and \U$30974 ( \31317 , \31316 , \31119 );
and \U$30975 ( \31318 , \31111 , \3406 );
or \U$30976 ( \31319 , \31317 , \31318 );
not \U$30977 ( \31320 , \31319 );
and \U$30978 ( \31321 , \31315 , \31320 );
and \U$30979 ( \31322 , \31314 , \31319 );
nor \U$30980 ( \31323 , \31321 , \31322 );
not \U$30981 ( \31324 , \31102 );
nand \U$30982 ( \31325 , \31324 , \31120 );
not \U$30983 ( \31326 , \25931 );
not \U$30984 ( \31327 , \25942 );
or \U$30985 ( \31328 , \31326 , \31327 );
or \U$30986 ( \31329 , \25942 , \25931 );
nand \U$30987 ( \31330 , \31328 , \31329 );
not \U$30988 ( \31331 , \31330 );
not \U$30989 ( \31332 , \25923 );
and \U$30990 ( \31333 , \31331 , \31332 );
and \U$30991 ( \31334 , \31330 , \25923 );
nor \U$30992 ( \31335 , \31333 , \31334 );
xor \U$30993 ( \31336 , \31325 , \31335 );
not \U$30994 ( \31337 , \31148 );
not \U$30995 ( \31338 , \31195 );
and \U$30996 ( \31339 , \31337 , \31338 );
and \U$30997 ( \31340 , \31195 , \31148 );
nor \U$30998 ( \31341 , \31340 , \31172 );
nor \U$30999 ( \31342 , \31339 , \31341 );
xor \U$31000 ( \31343 , \31336 , \31342 );
xnor \U$31001 ( \31344 , \31323 , \31343 );
not \U$31002 ( \31345 , \31344 );
and \U$31003 ( \31346 , \3254 , RI9870420_85);
and \U$31004 ( \31347 , RI9870510_87, \3252 );
nor \U$31005 ( \31348 , \31346 , \31347 );
not \U$31006 ( \31349 , \31348 );
not \U$31007 ( \31350 , \3406 );
and \U$31008 ( \31351 , \31349 , \31350 );
and \U$31009 ( \31352 , \31348 , \2935 );
nor \U$31010 ( \31353 , \31351 , \31352 );
not \U$31011 ( \31354 , \31353 );
xor \U$31012 ( \31355 , \25841 , \25849 );
xor \U$31013 ( \31356 , \31355 , \25857 );
not \U$31014 ( \31357 , \31356 );
or \U$31015 ( \31358 , \31354 , \31357 );
or \U$31016 ( \31359 , \31356 , \31353 );
nand \U$31017 ( \31360 , \31358 , \31359 );
not \U$31018 ( \31361 , \31360 );
not \U$31019 ( \31362 , \25875 );
not \U$31020 ( \31363 , \25886 );
or \U$31021 ( \31364 , \31362 , \31363 );
or \U$31022 ( \31365 , \25875 , \25886 );
nand \U$31023 ( \31366 , \31364 , \31365 );
not \U$31024 ( \31367 , \31366 );
not \U$31025 ( \31368 , \25868 );
and \U$31026 ( \31369 , \31367 , \31368 );
and \U$31027 ( \31370 , \31366 , \25868 );
nor \U$31028 ( \31371 , \31369 , \31370 );
not \U$31029 ( \31372 , \31371 );
and \U$31030 ( \31373 , \31361 , \31372 );
and \U$31031 ( \31374 , \31360 , \31371 );
nor \U$31032 ( \31375 , \31373 , \31374 );
not \U$31033 ( \31376 , \31375 );
not \U$31034 ( \31377 , \31009 );
not \U$31035 ( \31378 , \31018 );
and \U$31036 ( \31379 , \31377 , \31378 );
and \U$31037 ( \31380 , \31018 , \31009 );
nor \U$31038 ( \31381 , \31380 , \31025 );
nor \U$31039 ( \31382 , \31379 , \31381 );
xor \U$31040 ( \31383 , \31156 , \31163 );
and \U$31041 ( \31384 , \31383 , \31171 );
and \U$31042 ( \31385 , \31156 , \31163 );
or \U$31043 ( \31386 , \31384 , \31385 );
xor \U$31044 ( \31387 , \31382 , \31386 );
xor \U$31045 ( \31388 , \31132 , \31139 );
and \U$31046 ( \31389 , \31388 , \31147 );
and \U$31047 ( \31390 , \31132 , \31139 );
or \U$31048 ( \31391 , \31389 , \31390 );
xor \U$31049 ( \31392 , \31387 , \31391 );
not \U$31050 ( \31393 , \25820 );
not \U$31051 ( \31394 , \25831 );
or \U$31052 ( \31395 , \31393 , \31394 );
or \U$31053 ( \31396 , \25820 , \25831 );
nand \U$31054 ( \31397 , \31395 , \31396 );
not \U$31055 ( \31398 , \31397 );
not \U$31056 ( \31399 , \25813 );
and \U$31057 ( \31400 , \31398 , \31399 );
and \U$31058 ( \31401 , \31397 , \25813 );
nor \U$31059 ( \31402 , \31400 , \31401 );
xor \U$31060 ( \31403 , \25898 , \25905 );
xor \U$31061 ( \31404 , \31403 , \25913 );
xor \U$31062 ( \31405 , \31402 , \31404 );
not \U$31063 ( \31406 , \25959 );
not \U$31064 ( \31407 , \25970 );
or \U$31065 ( \31408 , \31406 , \31407 );
or \U$31066 ( \31409 , \25959 , \25970 );
nand \U$31067 ( \31410 , \31408 , \31409 );
not \U$31068 ( \31411 , \31410 );
not \U$31069 ( \31412 , \25952 );
and \U$31070 ( \31413 , \31411 , \31412 );
and \U$31071 ( \31414 , \31410 , \25952 );
nor \U$31072 ( \31415 , \31413 , \31414 );
xor \U$31073 ( \31416 , \31405 , \31415 );
xor \U$31074 ( \31417 , \31392 , \31416 );
not \U$31075 ( \31418 , \31417 );
or \U$31076 ( \31419 , \31376 , \31418 );
or \U$31077 ( \31420 , \31417 , \31375 );
nand \U$31078 ( \31421 , \31419 , \31420 );
not \U$31079 ( \31422 , \31421 );
and \U$31080 ( \31423 , \31345 , \31422 );
and \U$31081 ( \31424 , \31344 , \31421 );
nor \U$31082 ( \31425 , \31423 , \31424 );
not \U$31083 ( \31426 , \31425 );
or \U$31084 ( \31427 , \31303 , \31426 );
or \U$31085 ( \31428 , \31425 , \31302 );
nand \U$31086 ( \31429 , \31427 , \31428 );
not \U$31087 ( \31430 , \31429 );
and \U$31088 ( \31431 , \31288 , \31430 );
and \U$31089 ( \31432 , \31287 , \31429 );
nor \U$31090 ( \31433 , \31431 , \31432 );
xnor \U$31091 ( \31434 , \31246 , \31433 );
or \U$31092 ( \31435 , \31242 , \31434 );
or \U$31093 ( \31436 , \31246 , \31433 );
nand \U$31094 ( \31437 , \31435 , \31436 );
not \U$31095 ( \31438 , \31429 );
not \U$31096 ( \31439 , \31286 );
or \U$31097 ( \31440 , \31438 , \31439 );
or \U$31098 ( \31441 , \31286 , \31429 );
nand \U$31099 ( \31442 , \31441 , \31250 );
nand \U$31100 ( \31443 , \31440 , \31442 );
or \U$31101 ( \31444 , \31343 , \31323 );
not \U$31102 ( \31445 , \31323 );
not \U$31103 ( \31446 , \31343 );
or \U$31104 ( \31447 , \31445 , \31446 );
nand \U$31105 ( \31448 , \31447 , \31421 );
nand \U$31106 ( \31449 , \31444 , \31448 );
xor \U$31107 ( \31450 , \31292 , \31296 );
and \U$31108 ( \31451 , \31450 , \31301 );
and \U$31109 ( \31452 , \31292 , \31296 );
or \U$31110 ( \31453 , \31451 , \31452 );
xor \U$31111 ( \31454 , \31449 , \31453 );
xor \U$31112 ( \31455 , \31402 , \31404 );
and \U$31113 ( \31456 , \31455 , \31415 );
and \U$31114 ( \31457 , \31402 , \31404 );
nor \U$31115 ( \31458 , \31456 , \31457 );
xor \U$31116 ( \31459 , \25724 , \2263 );
xor \U$31117 ( \31460 , \31459 , \25732 );
xor \U$31118 ( \31461 , \31458 , \31460 );
xor \U$31119 ( \31462 , \26052 , \26058 );
xor \U$31120 ( \31463 , \31462 , \26065 );
xor \U$31121 ( \31464 , \31461 , \31463 );
xor \U$31122 ( \31465 , \31382 , \31386 );
and \U$31123 ( \31466 , \31465 , \31391 );
and \U$31124 ( \31467 , \31382 , \31386 );
nor \U$31125 ( \31468 , \31466 , \31467 );
not \U$31126 ( \31469 , \31319 );
not \U$31127 ( \31470 , \31313 );
or \U$31128 ( \31471 , \31469 , \31470 );
or \U$31129 ( \31472 , \31313 , \31319 );
nand \U$31130 ( \31473 , \31472 , \31309 );
nand \U$31131 ( \31474 , \31471 , \31473 );
xor \U$31132 ( \31475 , \31468 , \31474 );
or \U$31133 ( \31476 , \31371 , \31353 );
not \U$31134 ( \31477 , \31353 );
not \U$31135 ( \31478 , \31371 );
or \U$31136 ( \31479 , \31477 , \31478 );
nand \U$31137 ( \31480 , \31479 , \31356 );
nand \U$31138 ( \31481 , \31476 , \31480 );
xor \U$31139 ( \31482 , \31475 , \31481 );
xor \U$31140 ( \31483 , \25833 , \25860 );
xor \U$31141 ( \31484 , \31483 , \25888 );
xor \U$31142 ( \31485 , \25916 , \25944 );
xor \U$31143 ( \31486 , \31485 , \25972 );
xor \U$31144 ( \31487 , \25982 , \25988 );
xor \U$31145 ( \31488 , \31487 , \25995 );
xor \U$31146 ( \31489 , \31486 , \31488 );
xor \U$31147 ( \31490 , \31484 , \31489 );
xor \U$31148 ( \31491 , \31482 , \31490 );
xor \U$31149 ( \31492 , \31464 , \31491 );
xor \U$31150 ( \31493 , \31454 , \31492 );
not \U$31151 ( \31494 , \31493 );
not \U$31152 ( \31495 , \31425 );
nand \U$31153 ( \31496 , \31495 , \31302 );
xor \U$31154 ( \31497 , \31254 , \31258 );
and \U$31155 ( \31498 , \31497 , \31263 );
and \U$31156 ( \31499 , \31254 , \31258 );
or \U$31157 ( \31500 , \31498 , \31499 );
xor \U$31158 ( \31501 , \31325 , \31335 );
and \U$31159 ( \31502 , \31501 , \31342 );
and \U$31160 ( \31503 , \31325 , \31335 );
or \U$31161 ( \31504 , \31502 , \31503 );
xor \U$31162 ( \31505 , \31500 , \31504 );
not \U$31163 ( \31506 , \31375 );
not \U$31164 ( \31507 , \31392 );
and \U$31165 ( \31508 , \31506 , \31507 );
and \U$31166 ( \31509 , \31375 , \31392 );
nor \U$31167 ( \31510 , \31509 , \31416 );
nor \U$31168 ( \31511 , \31508 , \31510 );
xor \U$31169 ( \31512 , \31505 , \31511 );
xor \U$31170 ( \31513 , \31496 , \31512 );
not \U$31171 ( \31514 , \31281 );
not \U$31172 ( \31515 , \31264 );
and \U$31173 ( \31516 , \31514 , \31515 );
and \U$31174 ( \31517 , \31281 , \31264 );
nor \U$31175 ( \31518 , \31517 , \31272 );
nor \U$31176 ( \31519 , \31516 , \31518 );
xor \U$31177 ( \31520 , \31513 , \31519 );
not \U$31178 ( \31521 , \31520 );
or \U$31179 ( \31522 , \31494 , \31521 );
or \U$31180 ( \31523 , \31520 , \31493 );
nand \U$31181 ( \31524 , \31522 , \31523 );
xor \U$31182 ( \31525 , \31443 , \31524 );
and \U$31183 ( \31526 , \31437 , \31525 );
and \U$31184 ( \31527 , \31443 , \31524 );
nor \U$31185 ( \31528 , \31526 , \31527 );
not \U$31186 ( \31529 , \31520 );
nand \U$31187 ( \31530 , \31529 , \31493 );
xor \U$31188 ( \31531 , \31449 , \31453 );
and \U$31189 ( \31532 , \31531 , \31492 );
and \U$31190 ( \31533 , \31449 , \31453 );
or \U$31191 ( \31534 , \31532 , \31533 );
xor \U$31192 ( \31535 , \25833 , \25860 );
xor \U$31193 ( \31536 , \31535 , \25888 );
and \U$31194 ( \31537 , \31486 , \31536 );
xor \U$31195 ( \31538 , \25833 , \25860 );
xor \U$31196 ( \31539 , \31538 , \25888 );
and \U$31197 ( \31540 , \31488 , \31539 );
and \U$31198 ( \31541 , \31486 , \31488 );
or \U$31199 ( \31542 , \31537 , \31540 , \31541 );
xor \U$31200 ( \31543 , \31468 , \31474 );
and \U$31201 ( \31544 , \31543 , \31481 );
and \U$31202 ( \31545 , \31468 , \31474 );
or \U$31203 ( \31546 , \31544 , \31545 );
xor \U$31204 ( \31547 , \31542 , \31546 );
xor \U$31205 ( \31548 , \31458 , \31460 );
and \U$31206 ( \31549 , \31548 , \31463 );
and \U$31207 ( \31550 , \31458 , \31460 );
or \U$31208 ( \31551 , \31549 , \31550 );
xor \U$31209 ( \31552 , \31547 , \31551 );
xor \U$31210 ( \31553 , \31534 , \31552 );
not \U$31211 ( \31554 , \26003 );
xor \U$31212 ( \31555 , \26019 , \26014 );
not \U$31213 ( \31556 , \31555 );
or \U$31214 ( \31557 , \31554 , \31556 );
or \U$31215 ( \31558 , \31555 , \26003 );
nand \U$31216 ( \31559 , \31557 , \31558 );
xor \U$31217 ( \31560 , \25891 , \25975 );
xor \U$31218 ( \31561 , \31560 , \25998 );
xor \U$31219 ( \31562 , \31559 , \31561 );
not \U$31220 ( \31563 , \26043 );
xor \U$31221 ( \31564 , \26068 , \26032 );
not \U$31222 ( \31565 , \31564 );
or \U$31223 ( \31566 , \31563 , \31565 );
or \U$31224 ( \31567 , \31564 , \26043 );
nand \U$31225 ( \31568 , \31566 , \31567 );
xor \U$31226 ( \31569 , \31562 , \31568 );
not \U$31227 ( \31570 , \31569 );
xor \U$31228 ( \31571 , \31458 , \31460 );
xor \U$31229 ( \31572 , \31571 , \31463 );
and \U$31230 ( \31573 , \31482 , \31572 );
xor \U$31231 ( \31574 , \31458 , \31460 );
xor \U$31232 ( \31575 , \31574 , \31463 );
and \U$31233 ( \31576 , \31490 , \31575 );
and \U$31234 ( \31577 , \31482 , \31490 );
or \U$31235 ( \31578 , \31573 , \31576 , \31577 );
not \U$31236 ( \31579 , \31578 );
xor \U$31237 ( \31580 , \31500 , \31504 );
and \U$31238 ( \31581 , \31580 , \31511 );
and \U$31239 ( \31582 , \31500 , \31504 );
or \U$31240 ( \31583 , \31581 , \31582 );
not \U$31241 ( \31584 , \31583 );
and \U$31242 ( \31585 , \31579 , \31584 );
and \U$31243 ( \31586 , \31578 , \31583 );
nor \U$31244 ( \31587 , \31585 , \31586 );
not \U$31245 ( \31588 , \31587 );
or \U$31246 ( \31589 , \31570 , \31588 );
or \U$31247 ( \31590 , \31587 , \31569 );
nand \U$31248 ( \31591 , \31589 , \31590 );
xor \U$31249 ( \31592 , \31553 , \31591 );
not \U$31250 ( \31593 , \31592 );
xor \U$31251 ( \31594 , \31496 , \31512 );
and \U$31252 ( \31595 , \31594 , \31519 );
and \U$31253 ( \31596 , \31496 , \31512 );
or \U$31254 ( \31597 , \31595 , \31596 );
not \U$31255 ( \31598 , \31597 );
and \U$31256 ( \31599 , \31593 , \31598 );
and \U$31257 ( \31600 , \31592 , \31597 );
nor \U$31258 ( \31601 , \31599 , \31600 );
xnor \U$31259 ( \31602 , \31530 , \31601 );
or \U$31260 ( \31603 , \31528 , \31602 );
or \U$31261 ( \31604 , \31530 , \31601 );
nand \U$31262 ( \31605 , \31603 , \31604 );
not \U$31263 ( \31606 , \31592 );
nor \U$31264 ( \31607 , \31606 , \31597 );
xor \U$31265 ( \31608 , \31534 , \31552 );
and \U$31266 ( \31609 , \31608 , \31591 );
and \U$31267 ( \31610 , \31534 , \31552 );
or \U$31268 ( \31611 , \31609 , \31610 );
not \U$31269 ( \31612 , \31611 );
xor \U$31270 ( \31613 , \31542 , \31546 );
and \U$31271 ( \31614 , \31613 , \31551 );
and \U$31272 ( \31615 , \31542 , \31546 );
or \U$31273 ( \31616 , \31614 , \31615 );
xor \U$31274 ( \31617 , \25504 , \25506 );
xor \U$31275 ( \31618 , \31617 , \25519 );
xor \U$31276 ( \31619 , \31616 , \31618 );
xor \U$31277 ( \31620 , \31559 , \31561 );
and \U$31278 ( \31621 , \31620 , \31568 );
and \U$31279 ( \31622 , \31559 , \31561 );
or \U$31280 ( \31623 , \31621 , \31622 );
xor \U$31281 ( \31624 , \31619 , \31623 );
not \U$31282 ( \31625 , \31624 );
and \U$31283 ( \31626 , \31569 , \31578 );
not \U$31284 ( \31627 , \31569 );
not \U$31285 ( \31628 , \31578 );
and \U$31286 ( \31629 , \31627 , \31628 );
nor \U$31287 ( \31630 , \31629 , \31583 );
nor \U$31288 ( \31631 , \31626 , \31630 );
not \U$31289 ( \31632 , \31631 );
or \U$31290 ( \31633 , \31625 , \31632 );
or \U$31291 ( \31634 , \31631 , \31624 );
nand \U$31292 ( \31635 , \31633 , \31634 );
not \U$31293 ( \31636 , \31635 );
not \U$31294 ( \31637 , \25654 );
not \U$31295 ( \31638 , \25737 );
or \U$31296 ( \31639 , \31637 , \31638 );
or \U$31297 ( \31640 , \25737 , \25654 );
nand \U$31298 ( \31641 , \31639 , \31640 );
not \U$31299 ( \31642 , \31641 );
not \U$31300 ( \31643 , \25608 );
and \U$31301 ( \31644 , \31642 , \31643 );
and \U$31302 ( \31645 , \31641 , \25608 );
nor \U$31303 ( \31646 , \31644 , \31645 );
xor \U$31304 ( \31647 , \26001 , \26021 );
xor \U$31305 ( \31648 , \31647 , \26070 );
xnor \U$31306 ( \31649 , \31646 , \31648 );
not \U$31307 ( \31650 , \31649 );
xor \U$31308 ( \31651 , \25273 , \25298 );
xor \U$31309 ( \31652 , \31651 , \25326 );
xor \U$31310 ( \31653 , \26075 , \26082 );
xor \U$31311 ( \31654 , \31652 , \31653 );
not \U$31312 ( \31655 , \31654 );
and \U$31313 ( \31656 , \31650 , \31655 );
and \U$31314 ( \31657 , \31649 , \31654 );
nor \U$31315 ( \31658 , \31656 , \31657 );
not \U$31316 ( \31659 , \31658 );
and \U$31317 ( \31660 , \31636 , \31659 );
and \U$31318 ( \31661 , \31635 , \31658 );
nor \U$31319 ( \31662 , \31660 , \31661 );
not \U$31320 ( \31663 , \31662 );
or \U$31321 ( \31664 , \31612 , \31663 );
or \U$31322 ( \31665 , \31662 , \31611 );
nand \U$31323 ( \31666 , \31664 , \31665 );
xor \U$31324 ( \31667 , \31607 , \31666 );
and \U$31325 ( \31668 , \31605 , \31667 );
and \U$31326 ( \31669 , \31607 , \31666 );
nor \U$31327 ( \31670 , \31668 , \31669 );
not \U$31328 ( \31671 , \31662 );
nand \U$31329 ( \31672 , \31671 , \31611 );
xor \U$31330 ( \31673 , \31616 , \31618 );
and \U$31331 ( \31674 , \31673 , \31623 );
and \U$31332 ( \31675 , \31616 , \31618 );
or \U$31333 ( \31676 , \31674 , \31675 );
xor \U$31334 ( \31677 , \25522 , \25739 );
xor \U$31335 ( \31678 , \31677 , \25754 );
xor \U$31336 ( \31679 , \31676 , \31678 );
or \U$31337 ( \31680 , \31648 , \31646 );
not \U$31338 ( \31681 , \31646 );
not \U$31339 ( \31682 , \31648 );
or \U$31340 ( \31683 , \31681 , \31682 );
nand \U$31341 ( \31684 , \31683 , \31654 );
nand \U$31342 ( \31685 , \31680 , \31684 );
xor \U$31343 ( \31686 , \31679 , \31685 );
or \U$31344 ( \31687 , \31658 , \31631 );
not \U$31345 ( \31688 , \31631 );
not \U$31346 ( \31689 , \31658 );
or \U$31347 ( \31690 , \31688 , \31689 );
nand \U$31348 ( \31691 , \31690 , \31624 );
nand \U$31349 ( \31692 , \31687 , \31691 );
xnor \U$31350 ( \31693 , \31686 , \31692 );
not \U$31351 ( \31694 , \31693 );
xor \U$31352 ( \31695 , \26073 , \26087 );
xor \U$31353 ( \31696 , \31695 , \26092 );
not \U$31354 ( \31697 , \31696 );
and \U$31355 ( \31698 , \31694 , \31697 );
and \U$31356 ( \31699 , \31693 , \31696 );
nor \U$31357 ( \31700 , \31698 , \31699 );
xnor \U$31358 ( \31701 , \31672 , \31700 );
or \U$31359 ( \31702 , \31670 , \31701 );
or \U$31360 ( \31703 , \31672 , \31700 );
nand \U$31361 ( \31704 , \31702 , \31703 );
xor \U$31362 ( \31705 , \31676 , \31678 );
and \U$31363 ( \31706 , \31705 , \31685 );
and \U$31364 ( \31707 , \31676 , \31678 );
or \U$31365 ( \31708 , \31706 , \31707 );
not \U$31366 ( \31709 , \31708 );
xnor \U$31367 ( \31710 , \26095 , \25803 );
not \U$31368 ( \31711 , \31710 );
not \U$31369 ( \31712 , \25800 );
and \U$31370 ( \31713 , \31711 , \31712 );
and \U$31371 ( \31714 , \31710 , \25800 );
nor \U$31372 ( \31715 , \31713 , \31714 );
not \U$31373 ( \31716 , \31715 );
or \U$31374 ( \31717 , \31709 , \31716 );
or \U$31375 ( \31718 , \31715 , \31708 );
nand \U$31376 ( \31719 , \31717 , \31718 );
not \U$31377 ( \31720 , \31696 );
not \U$31378 ( \31721 , \31686 );
or \U$31379 ( \31722 , \31720 , \31721 );
or \U$31380 ( \31723 , \31686 , \31696 );
nand \U$31381 ( \31724 , \31723 , \31692 );
nand \U$31382 ( \31725 , \31722 , \31724 );
xor \U$31383 ( \31726 , \31719 , \31725 );
and \U$31384 ( \31727 , \31704 , \31726 );
and \U$31385 ( \31728 , \31719 , \31725 );
nor \U$31386 ( \31729 , \31727 , \31728 );
not \U$31387 ( \31730 , \31715 );
nand \U$31388 ( \31731 , \31730 , \31708 );
xnor \U$31389 ( \31732 , \25793 , \26097 );
not \U$31390 ( \31733 , \31732 );
not \U$31391 ( \31734 , \25796 );
and \U$31392 ( \31735 , \31733 , \31734 );
and \U$31393 ( \31736 , \31732 , \25796 );
nor \U$31394 ( \31737 , \31735 , \31736 );
xnor \U$31395 ( \31738 , \31731 , \31737 );
or \U$31396 ( \31739 , \31729 , \31738 );
or \U$31397 ( \31740 , \31731 , \31737 );
nand \U$31398 ( \31741 , \31739 , \31740 );
and \U$31399 ( \31742 , \26101 , \31741 );
nor \U$31400 ( \31743 , \26100 , \31742 );
xnor \U$31401 ( \31744 , \25213 , \25476 );
not \U$31402 ( \31745 , \31744 );
not \U$31403 ( \31746 , \25216 );
and \U$31404 ( \31747 , \31745 , \31746 );
and \U$31405 ( \31748 , \31744 , \25216 );
nor \U$31406 ( \31749 , \31747 , \31748 );
xor \U$31407 ( \31750 , \25481 , \25483 );
and \U$31408 ( \31751 , \31750 , \25790 );
and \U$31409 ( \31752 , \25481 , \25483 );
nor \U$31410 ( \31753 , \31751 , \31752 );
xnor \U$31411 ( \31754 , \31749 , \31753 );
or \U$31412 ( \31755 , \31743 , \31754 );
or \U$31413 ( \31756 , \31749 , \31753 );
nand \U$31414 ( \31757 , \31755 , \31756 );
and \U$31415 ( \31758 , \25480 , \31757 );
nor \U$31416 ( \31759 , \25479 , \31758 );
xnor \U$31417 ( \31760 , \24927 , \24630 );
not \U$31418 ( \31761 , \31760 );
not \U$31419 ( \31762 , \24643 );
and \U$31420 ( \31763 , \31761 , \31762 );
and \U$31421 ( \31764 , \31760 , \24643 );
nor \U$31422 ( \31765 , \31763 , \31764 );
xor \U$31423 ( \31766 , \24942 , \25204 );
and \U$31424 ( \31767 , \31766 , \25207 );
and \U$31425 ( \31768 , \24942 , \25204 );
nor \U$31426 ( \31769 , \31767 , \31768 );
xnor \U$31427 ( \31770 , \31765 , \31769 );
or \U$31428 ( \31771 , \31759 , \31770 );
or \U$31429 ( \31772 , \31769 , \31765 );
nand \U$31430 ( \31773 , \31771 , \31772 );
and \U$31431 ( \31774 , \24941 , \31773 );
nor \U$31432 ( \31775 , \24940 , \31774 );
xor \U$31433 ( \31776 , \24931 , \24933 );
and \U$31434 ( \31777 , \31776 , \24938 );
and \U$31435 ( \31778 , \24931 , \24933 );
nor \U$31436 ( \31779 , \31777 , \31778 );
xnor \U$31437 ( \31780 , \24035 , \24345 );
not \U$31438 ( \31781 , \31780 );
not \U$31439 ( \31782 , \24038 );
and \U$31440 ( \31783 , \31781 , \31782 );
and \U$31441 ( \31784 , \31780 , \24038 );
nor \U$31442 ( \31785 , \31783 , \31784 );
xnor \U$31443 ( \31786 , \31779 , \31785 );
or \U$31444 ( \31787 , \31775 , \31786 );
or \U$31445 ( \31788 , \31779 , \31785 );
nand \U$31446 ( \31789 , \31787 , \31788 );
and \U$31447 ( \31790 , \24349 , \31789 );
nor \U$31448 ( \31791 , \24348 , \31790 );
xor \U$31449 ( \31792 , \23694 , \23696 );
and \U$31450 ( \31793 , \31792 , \24024 );
and \U$31451 ( \31794 , \23694 , \23696 );
nor \U$31452 ( \31795 , \31793 , \31794 );
xnor \U$31453 ( \31796 , \23674 , \23664 );
not \U$31454 ( \31797 , \31796 );
not \U$31455 ( \31798 , \23680 );
and \U$31456 ( \31799 , \31797 , \31798 );
and \U$31457 ( \31800 , \31796 , \23680 );
nor \U$31458 ( \31801 , \31799 , \31800 );
xnor \U$31459 ( \31802 , \31795 , \31801 );
or \U$31460 ( \31803 , \31791 , \31802 );
or \U$31461 ( \31804 , \31795 , \31801 );
nand \U$31462 ( \31805 , \31803 , \31804 );
and \U$31463 ( \31806 , \23684 , \31805 );
nor \U$31464 ( \31807 , \23683 , \31806 );
or \U$31465 ( \31808 , \23358 , \31807 );
nand \U$31466 ( \31809 , \23357 , \31808 );
not \U$31467 ( \31810 , \22682 );
not \U$31468 ( \31811 , \23033 );
or \U$31469 ( \31812 , \31810 , \31811 );
or \U$31470 ( \31813 , \23033 , \22682 );
nand \U$31471 ( \31814 , \31813 , \23027 );
nand \U$31472 ( \31815 , \31812 , \31814 );
xor \U$31473 ( \31816 , \22351 , \22353 );
xor \U$31474 ( \31817 , \31816 , \22672 );
xor \U$31475 ( \31818 , \31815 , \31817 );
and \U$31476 ( \31819 , \31809 , \31818 );
and \U$31477 ( \31820 , \31815 , \31817 );
nor \U$31478 ( \31821 , \31819 , \31820 );
or \U$31479 ( \31822 , \22677 , \31821 );
nand \U$31480 ( \31823 , \22676 , \31822 );
and \U$31481 ( \31824 , \22343 , \31823 );
nor \U$31482 ( \31825 , \22342 , \31824 );
or \U$31483 ( \31826 , \21969 , \31825 );
nand \U$31484 ( \31827 , \21968 , \31826 );
not \U$31485 ( \31828 , \21576 );
nor \U$31486 ( \31829 , \31828 , \21941 );
xor \U$31487 ( \31830 , \21197 , \21217 );
and \U$31488 ( \31831 , \31830 , \21575 );
and \U$31489 ( \31832 , \21197 , \21217 );
nor \U$31490 ( \31833 , \31831 , \31832 );
not \U$31491 ( \31834 , \31833 );
xor \U$31492 ( \31835 , \20802 , \21139 );
and \U$31493 ( \31836 , \31835 , \21196 );
and \U$31494 ( \31837 , \20802 , \21139 );
or \U$31495 ( \31838 , \31836 , \31837 );
xor \U$31496 ( \31839 , \19729 , \19749 );
xor \U$31497 ( \31840 , \31839 , \19760 );
and \U$31498 ( \31841 , \21189 , \31840 );
xor \U$31499 ( \31842 , \19729 , \19749 );
xor \U$31500 ( \31843 , \31842 , \19760 );
and \U$31501 ( \31844 , \21193 , \31843 );
and \U$31502 ( \31845 , \21189 , \21193 );
or \U$31503 ( \31846 , \31841 , \31844 , \31845 );
not \U$31504 ( \31847 , \31846 );
not \U$31505 ( \31848 , \31847 );
xor \U$31506 ( \31849 , \21170 , \21174 );
and \U$31507 ( \31850 , \31849 , \21183 );
and \U$31508 ( \31851 , \21170 , \21174 );
nor \U$31509 ( \31852 , \31850 , \31851 );
not \U$31510 ( \31853 , \21150 );
not \U$31511 ( \31854 , \21157 );
and \U$31512 ( \31855 , \31853 , \31854 );
and \U$31513 ( \31856 , \21150 , \21157 );
nor \U$31514 ( \31857 , \31856 , \21161 );
nor \U$31515 ( \31858 , \31855 , \31857 );
xor \U$31516 ( \31859 , \31852 , \31858 );
not \U$31517 ( \31860 , \31859 );
or \U$31518 ( \31861 , \31848 , \31860 );
or \U$31519 ( \31862 , \31859 , \31847 );
nand \U$31520 ( \31863 , \31861 , \31862 );
xor \U$31521 ( \31864 , \31838 , \31863 );
xor \U$31522 ( \31865 , \21166 , \21184 );
and \U$31523 ( \31866 , \31865 , \21195 );
and \U$31524 ( \31867 , \21166 , \21184 );
or \U$31525 ( \31868 , \31866 , \31867 );
xor \U$31526 ( \31869 , \21203 , \21207 );
and \U$31527 ( \31870 , \31869 , \21216 );
and \U$31528 ( \31871 , \21203 , \21207 );
or \U$31529 ( \31872 , \31870 , \31871 );
xor \U$31530 ( \31873 , \31868 , \31872 );
xor \U$31531 ( \31874 , \20038 , \20040 );
xor \U$31532 ( \31875 , \31874 , \20043 );
xor \U$31533 ( \31876 , \19763 , \20014 );
xor \U$31534 ( \31877 , \31876 , \20031 );
xor \U$31535 ( \31878 , \20051 , \20071 );
xor \U$31536 ( \31879 , \31878 , \20076 );
xor \U$31537 ( \31880 , \31877 , \31879 );
xor \U$31538 ( \31881 , \31875 , \31880 );
xor \U$31539 ( \31882 , \31873 , \31881 );
xor \U$31540 ( \31883 , \31864 , \31882 );
not \U$31541 ( \31884 , \31883 );
or \U$31542 ( \31885 , \31834 , \31884 );
or \U$31543 ( \31886 , \31883 , \31833 );
nand \U$31544 ( \31887 , \31885 , \31886 );
xor \U$31545 ( \31888 , \31829 , \31887 );
and \U$31546 ( \31889 , \31827 , \31888 );
and \U$31547 ( \31890 , \31829 , \31887 );
nor \U$31548 ( \31891 , \31889 , \31890 );
not \U$31549 ( \31892 , \31833 );
nand \U$31550 ( \31893 , \31892 , \31883 );
not \U$31551 ( \31894 , \31847 );
not \U$31552 ( \31895 , \31858 );
and \U$31553 ( \31896 , \31894 , \31895 );
and \U$31554 ( \31897 , \31847 , \31858 );
nor \U$31555 ( \31898 , \31897 , \31852 );
nor \U$31556 ( \31899 , \31896 , \31898 );
not \U$31557 ( \31900 , \31899 );
xor \U$31558 ( \31901 , \20038 , \20040 );
xor \U$31559 ( \31902 , \31901 , \20043 );
and \U$31560 ( \31903 , \31877 , \31902 );
xor \U$31561 ( \31904 , \20038 , \20040 );
xor \U$31562 ( \31905 , \31904 , \20043 );
and \U$31563 ( \31906 , \31879 , \31905 );
and \U$31564 ( \31907 , \31877 , \31879 );
or \U$31565 ( \31908 , \31903 , \31906 , \31907 );
not \U$31566 ( \31909 , \31908 );
or \U$31567 ( \31910 , \31900 , \31909 );
or \U$31568 ( \31911 , \31908 , \31899 );
nand \U$31569 ( \31912 , \31910 , \31911 );
not \U$31570 ( \31913 , \31912 );
not \U$31571 ( \31914 , \19655 );
not \U$31572 ( \31915 , \19677 );
or \U$31573 ( \31916 , \31914 , \31915 );
or \U$31574 ( \31917 , \19677 , \19655 );
nand \U$31575 ( \31918 , \31916 , \31917 );
not \U$31576 ( \31919 , \31918 );
not \U$31577 ( \31920 , \19657 );
and \U$31578 ( \31921 , \31919 , \31920 );
and \U$31579 ( \31922 , \31918 , \19657 );
nor \U$31580 ( \31923 , \31921 , \31922 );
not \U$31581 ( \31924 , \31923 );
and \U$31582 ( \31925 , \31913 , \31924 );
and \U$31583 ( \31926 , \31912 , \31923 );
nor \U$31584 ( \31927 , \31925 , \31926 );
not \U$31585 ( \31928 , \31927 );
xor \U$31586 ( \31929 , \31868 , \31872 );
and \U$31587 ( \31930 , \31929 , \31881 );
and \U$31588 ( \31931 , \31868 , \31872 );
or \U$31589 ( \31932 , \31930 , \31931 );
not \U$31590 ( \31933 , \31932 );
and \U$31591 ( \31934 , \31928 , \31933 );
and \U$31592 ( \31935 , \31927 , \31932 );
nor \U$31593 ( \31936 , \31934 , \31935 );
not \U$31594 ( \31937 , \31936 );
xor \U$31595 ( \31938 , \20084 , \20086 );
xor \U$31596 ( \31939 , \31938 , \20091 );
xor \U$31597 ( \31940 , \19544 , \19564 );
xor \U$31598 ( \31941 , \31940 , \19638 );
xor \U$31599 ( \31942 , \20034 , \20046 );
xor \U$31600 ( \31943 , \31942 , \20079 );
xor \U$31601 ( \31944 , \31941 , \31943 );
xor \U$31602 ( \31945 , \31939 , \31944 );
not \U$31603 ( \31946 , \31945 );
and \U$31604 ( \31947 , \31937 , \31946 );
and \U$31605 ( \31948 , \31936 , \31945 );
nor \U$31606 ( \31949 , \31947 , \31948 );
not \U$31607 ( \31950 , \31949 );
xor \U$31608 ( \31951 , \31838 , \31863 );
and \U$31609 ( \31952 , \31951 , \31882 );
and \U$31610 ( \31953 , \31838 , \31863 );
or \U$31611 ( \31954 , \31952 , \31953 );
not \U$31612 ( \31955 , \31954 );
and \U$31613 ( \31956 , \31950 , \31955 );
and \U$31614 ( \31957 , \31949 , \31954 );
nor \U$31615 ( \31958 , \31956 , \31957 );
xnor \U$31616 ( \31959 , \31893 , \31958 );
or \U$31617 ( \31960 , \31891 , \31959 );
or \U$31618 ( \31961 , \31893 , \31958 );
nand \U$31619 ( \31962 , \31960 , \31961 );
not \U$31620 ( \31963 , \31954 );
nor \U$31621 ( \31964 , \31963 , \31949 );
xor \U$31622 ( \31965 , \20082 , \20094 );
xor \U$31623 ( \31966 , \31965 , \20099 );
not \U$31624 ( \31967 , \31945 );
or \U$31625 ( \31968 , \31967 , \31927 );
not \U$31626 ( \31969 , \31927 );
not \U$31627 ( \31970 , \31967 );
or \U$31628 ( \31971 , \31969 , \31970 );
nand \U$31629 ( \31972 , \31971 , \31932 );
nand \U$31630 ( \31973 , \31968 , \31972 );
xor \U$31631 ( \31974 , \31966 , \31973 );
xor \U$31632 ( \31975 , \19296 , \19641 );
xor \U$31633 ( \31976 , \31975 , \19679 );
xor \U$31634 ( \31977 , \20084 , \20086 );
xor \U$31635 ( \31978 , \31977 , \20091 );
and \U$31636 ( \31979 , \31941 , \31978 );
xor \U$31637 ( \31980 , \20084 , \20086 );
xor \U$31638 ( \31981 , \31980 , \20091 );
and \U$31639 ( \31982 , \31943 , \31981 );
and \U$31640 ( \31983 , \31941 , \31943 );
or \U$31641 ( \31984 , \31979 , \31982 , \31983 );
xor \U$31642 ( \31985 , \31976 , \31984 );
or \U$31643 ( \31986 , \31899 , \31923 );
not \U$31644 ( \31987 , \31923 );
not \U$31645 ( \31988 , \31899 );
or \U$31646 ( \31989 , \31987 , \31988 );
nand \U$31647 ( \31990 , \31989 , \31908 );
nand \U$31648 ( \31991 , \31986 , \31990 );
xor \U$31649 ( \31992 , \31985 , \31991 );
xor \U$31650 ( \31993 , \31974 , \31992 );
xor \U$31651 ( \31994 , \31964 , \31993 );
and \U$31652 ( \31995 , \31962 , \31994 );
and \U$31653 ( \31996 , \31964 , \31993 );
nor \U$31654 ( \31997 , \31995 , \31996 );
xor \U$31655 ( \31998 , \19712 , \19714 );
xor \U$31656 ( \31999 , \31998 , \20102 );
not \U$31657 ( \32000 , \31999 );
xor \U$31658 ( \32001 , \31976 , \31984 );
and \U$31659 ( \32002 , \32001 , \31991 );
and \U$31660 ( \32003 , \31976 , \31984 );
nor \U$31661 ( \32004 , \32002 , \32003 );
not \U$31662 ( \32005 , \32004 );
and \U$31663 ( \32006 , \32000 , \32005 );
and \U$31664 ( \32007 , \31999 , \32004 );
nor \U$31665 ( \32008 , \32006 , \32007 );
xor \U$31666 ( \32009 , \31966 , \31973 );
and \U$31667 ( \32010 , \32009 , \31992 );
and \U$31668 ( \32011 , \31966 , \31973 );
nor \U$31669 ( \32012 , \32010 , \32011 );
xnor \U$31670 ( \32013 , \32008 , \32012 );
or \U$31671 ( \32014 , \31997 , \32013 );
or \U$31672 ( \32015 , \32008 , \32012 );
nand \U$31673 ( \32016 , \32014 , \32015 );
not \U$31674 ( \32017 , \31999 );
nor \U$31675 ( \32018 , \32017 , \32004 );
not \U$31676 ( \32019 , \20105 );
not \U$31677 ( \32020 , \20110 );
or \U$31678 ( \32021 , \32019 , \32020 );
or \U$31679 ( \32022 , \20110 , \20105 );
nand \U$31680 ( \32023 , \32021 , \32022 );
xor \U$31681 ( \32024 , \32018 , \32023 );
and \U$31682 ( \32025 , \32016 , \32024 );
and \U$31683 ( \32026 , \32018 , \32023 );
nor \U$31684 ( \32027 , \32025 , \32026 );
or \U$31685 ( \32028 , \20113 , \32027 );
nand \U$31686 ( \32029 , \20112 , \32028 );
and \U$31687 ( \32030 , \19704 , \32029 );
nor \U$31688 ( \32031 , \19703 , \32030 );
xor \U$31689 ( \32032 , \19204 , \19206 );
xor \U$31690 ( \32033 , \32032 , \19209 );
and \U$31691 ( \32034 , \19234 , \32033 );
xor \U$31692 ( \32035 , \19204 , \19206 );
xor \U$31693 ( \32036 , \32035 , \19209 );
and \U$31694 ( \32037 , \19254 , \32036 );
and \U$31695 ( \32038 , \19234 , \19254 );
or \U$31696 ( \32039 , \32034 , \32037 , \32038 );
xor \U$31697 ( \32040 , \17484 , \17527 );
xor \U$31698 ( \32041 , \32040 , \17548 );
not \U$31699 ( \32042 , \32041 );
xor \U$31700 ( \32043 , \17653 , \17659 );
xor \U$31701 ( \32044 , \32043 , \18048 );
not \U$31702 ( \32045 , \32044 );
or \U$31703 ( \32046 , \32042 , \32045 );
or \U$31704 ( \32047 , \32044 , \32041 );
nand \U$31705 ( \32048 , \32046 , \32047 );
xor \U$31706 ( \32049 , \32039 , \32048 );
xor \U$31707 ( \32050 , \19204 , \19206 );
and \U$31708 ( \32051 , \32050 , \19209 );
and \U$31709 ( \32052 , \19204 , \19206 );
or \U$31710 ( \32053 , \32051 , \32052 );
xor \U$31711 ( \32054 , \17567 , \17573 );
xor \U$31712 ( \32055 , \32054 , \17580 );
xor \U$31713 ( \32056 , \32053 , \32055 );
xor \U$31714 ( \32057 , \19238 , \19244 );
and \U$31715 ( \32058 , \32057 , \19253 );
and \U$31716 ( \32059 , \19238 , \19244 );
or \U$31717 ( \32060 , \32058 , \32059 );
xor \U$31718 ( \32061 , \32056 , \32060 );
xor \U$31719 ( \32062 , \32049 , \32061 );
not \U$31720 ( \32063 , \32062 );
not \U$31721 ( \32064 , \19201 );
nand \U$31722 ( \32065 , \32064 , \19256 );
not \U$31723 ( \32066 , \32065 );
and \U$31724 ( \32067 , \32063 , \32066 );
and \U$31725 ( \32068 , \32062 , \32065 );
nor \U$31726 ( \32069 , \32067 , \32068 );
or \U$31727 ( \32070 , \32031 , \32069 );
not \U$31728 ( \32071 , \32062 );
or \U$31729 ( \32072 , \32065 , \32071 );
nand \U$31730 ( \32073 , \32070 , \32072 );
not \U$31731 ( \32074 , \18051 );
not \U$31732 ( \32075 , \17629 );
or \U$31733 ( \32076 , \32074 , \32075 );
or \U$31734 ( \32077 , \17629 , \18051 );
nand \U$31735 ( \32078 , \32076 , \32077 );
not \U$31736 ( \32079 , \32078 );
not \U$31737 ( \32080 , \17635 );
and \U$31738 ( \32081 , \32079 , \32080 );
and \U$31739 ( \32082 , \32078 , \17635 );
nor \U$31740 ( \32083 , \32081 , \32082 );
not \U$31741 ( \32084 , \32083 );
not \U$31742 ( \32085 , \32041 );
nand \U$31743 ( \32086 , \32085 , \32044 );
not \U$31744 ( \32087 , \32086 );
xor \U$31745 ( \32088 , \32053 , \32055 );
and \U$31746 ( \32089 , \32088 , \32060 );
and \U$31747 ( \32090 , \32053 , \32055 );
or \U$31748 ( \32091 , \32089 , \32090 );
not \U$31749 ( \32092 , \32091 );
or \U$31750 ( \32093 , \32087 , \32092 );
or \U$31751 ( \32094 , \32091 , \32086 );
nand \U$31752 ( \32095 , \32093 , \32094 );
not \U$31753 ( \32096 , \32095 );
or \U$31754 ( \32097 , \32084 , \32096 );
or \U$31755 ( \32098 , \32095 , \32083 );
nand \U$31756 ( \32099 , \32097 , \32098 );
xor \U$31757 ( \32100 , \32039 , \32048 );
and \U$31758 ( \32101 , \32100 , \32061 );
and \U$31759 ( \32102 , \32039 , \32048 );
or \U$31760 ( \32103 , \32101 , \32102 );
xor \U$31761 ( \32104 , \32099 , \32103 );
and \U$31762 ( \32105 , \32073 , \32104 );
and \U$31763 ( \32106 , \32103 , \32099 );
nor \U$31764 ( \32107 , \32105 , \32106 );
not \U$31765 ( \32108 , \32083 );
not \U$31766 ( \32109 , \32086 );
and \U$31767 ( \32110 , \32108 , \32109 );
and \U$31768 ( \32111 , \32083 , \32086 );
not \U$31769 ( \32112 , \32091 );
nor \U$31770 ( \32113 , \32111 , \32112 );
nor \U$31771 ( \32114 , \32110 , \32113 );
xnor \U$31772 ( \32115 , \18053 , \17616 );
not \U$31773 ( \32116 , \32115 );
not \U$31774 ( \32117 , \17613 );
and \U$31775 ( \32118 , \32116 , \32117 );
and \U$31776 ( \32119 , \32115 , \17613 );
nor \U$31777 ( \32120 , \32118 , \32119 );
xnor \U$31778 ( \32121 , \32114 , \32120 );
or \U$31779 ( \32122 , \32107 , \32121 );
or \U$31780 ( \32123 , \32114 , \32120 );
nand \U$31781 ( \32124 , \32122 , \32123 );
and \U$31782 ( \32125 , \18057 , \32124 );
nor \U$31783 ( \32126 , \18056 , \32125 );
and \U$31784 ( \32127 , \17607 , \17122 );
not \U$31785 ( \32128 , \17607 );
not \U$31786 ( \32129 , \17122 );
and \U$31787 ( \32130 , \32128 , \32129 );
nor \U$31788 ( \32131 , \32130 , \17116 );
nor \U$31789 ( \32132 , \32127 , \32131 );
xor \U$31790 ( \32133 , \16582 , \16586 );
xor \U$31791 ( \32134 , \32133 , \16594 );
not \U$31792 ( \32135 , \17112 );
not \U$31793 ( \32136 , \17109 );
or \U$31794 ( \32137 , \32135 , \32136 );
or \U$31795 ( \32138 , \17109 , \17112 );
nand \U$31796 ( \32139 , \32138 , \17107 );
nand \U$31797 ( \32140 , \32137 , \32139 );
xnor \U$31798 ( \32141 , \32134 , \32140 );
not \U$31799 ( \32142 , \32141 );
xor \U$31800 ( \32143 , \15622 , \16096 );
not \U$31801 ( \32144 , \32143 );
and \U$31802 ( \32145 , \32142 , \32144 );
and \U$31803 ( \32146 , \32141 , \32143 );
nor \U$31804 ( \32147 , \32145 , \32146 );
xnor \U$31805 ( \32148 , \32132 , \32147 );
or \U$31806 ( \32149 , \32126 , \32148 );
or \U$31807 ( \32150 , \32132 , \32147 );
nand \U$31808 ( \32151 , \32149 , \32150 );
not \U$31809 ( \32152 , \32143 );
not \U$31810 ( \32153 , \32134 );
or \U$31811 ( \32154 , \32152 , \32153 );
or \U$31812 ( \32155 , \32134 , \32143 );
nand \U$31813 ( \32156 , \32155 , \32140 );
nand \U$31814 ( \32157 , \32154 , \32156 );
xor \U$31815 ( \32158 , \16097 , \16597 );
xor \U$31816 ( \32159 , \32158 , \16608 );
xor \U$31817 ( \32160 , \32157 , \32159 );
and \U$31818 ( \32161 , \32151 , \32160 );
and \U$31819 ( \32162 , \32157 , \32159 );
nor \U$31820 ( \32163 , \32161 , \32162 );
xnor \U$31821 ( \32164 , \16611 , \16630 );
or \U$31822 ( \32165 , \32163 , \32164 );
nand \U$31823 ( \32166 , \16632 , \32165 );
xor \U$31824 ( \32167 , \16620 , \16626 );
and \U$31825 ( \32168 , \32167 , \16629 );
and \U$31826 ( \32169 , \16620 , \16626 );
or \U$31827 ( \32170 , \32168 , \32169 );
not \U$31828 ( \32171 , \15613 );
not \U$31829 ( \32172 , \15157 );
or \U$31830 ( \32173 , \32171 , \32172 );
or \U$31831 ( \32174 , \15157 , \15613 );
nand \U$31832 ( \32175 , \32173 , \32174 );
xor \U$31833 ( \32176 , \32170 , \32175 );
and \U$31834 ( \32177 , \32166 , \32176 );
and \U$31835 ( \32178 , \32175 , \32170 );
nor \U$31836 ( \32179 , \32177 , \32178 );
or \U$31837 ( \32180 , \15620 , \32179 );
nand \U$31838 ( \32181 , \15615 , \32180 );
and \U$31839 ( \32182 , \15144 , \32181 );
nor \U$31840 ( \32183 , \15143 , \32182 );
or \U$31841 ( \32184 , \14676 , \32183 );
nand \U$31842 ( \32185 , \14671 , \32184 );
and \U$31843 ( \32186 , \14208 , \14210 );
xor \U$31844 ( \32187 , \13730 , \13732 );
xor \U$31845 ( \32188 , \32187 , \13735 );
xor \U$31846 ( \32189 , \32186 , \32188 );
and \U$31847 ( \32190 , \32185 , \32189 );
and \U$31848 ( \32191 , \32186 , \32188 );
nor \U$31849 ( \32192 , \32190 , \32191 );
xnor \U$31850 ( \32193 , \13291 , \13738 );
or \U$31851 ( \32194 , \32192 , \32193 );
nand \U$31852 ( \32195 , \13740 , \32194 );
and \U$31853 ( \32196 , \13288 , \13290 );
xor \U$31854 ( \32197 , \12865 , \12875 );
xor \U$31855 ( \32198 , \32196 , \32197 );
and \U$31856 ( \32199 , \32195 , \32198 );
and \U$31857 ( \32200 , \32196 , \32197 );
nor \U$31858 ( \32201 , \32199 , \32200 );
xnor \U$31859 ( \32202 , \12876 , \12884 );
or \U$31860 ( \32203 , \32201 , \32202 );
nand \U$31861 ( \32204 , \12886 , \32203 );
and \U$31862 ( \32205 , \12881 , \12883 );
xor \U$31863 ( \32206 , \12054 , \12064 );
xor \U$31864 ( \32207 , \32205 , \32206 );
and \U$31865 ( \32208 , \32204 , \32207 );
and \U$31866 ( \32209 , \32205 , \32206 );
nor \U$31867 ( \32210 , \32208 , \32209 );
xnor \U$31868 ( \32211 , \12065 , \12075 );
or \U$31869 ( \32212 , \32210 , \32211 );
nand \U$31870 ( \32213 , \12077 , \32212 );
and \U$31871 ( \32214 , \12070 , \12074 );
xor \U$31872 ( \32215 , \11169 , \11259 );
xor \U$31873 ( \32216 , \32214 , \32215 );
and \U$31874 ( \32217 , \32213 , \32216 );
and \U$31875 ( \32218 , \32214 , \32215 );
nor \U$31876 ( \32219 , \32217 , \32218 );
xnor \U$31877 ( \32220 , \11260 , \11314 );
or \U$31878 ( \32221 , \32219 , \32220 );
nand \U$31879 ( \32222 , \11316 , \32221 );
and \U$31880 ( \32223 , \11265 , \11313 );
xor \U$31881 ( \32224 , \11269 , \11280 );
and \U$31882 ( \32225 , \32224 , \11312 );
and \U$31883 ( \32226 , \11269 , \11280 );
or \U$31884 ( \32227 , \32225 , \32226 );
not \U$31885 ( \32228 , \32227 );
and \U$31886 ( \32229 , \11307 , \11303 );
not \U$31887 ( \32230 , \11303 );
not \U$31888 ( \32231 , \11307 );
and \U$31889 ( \32232 , \32230 , \32231 );
nor \U$31890 ( \32233 , \32232 , \11294 );
nor \U$31891 ( \32234 , \32229 , \32233 );
xor \U$31892 ( \32235 , \9433 , \9447 );
xor \U$31893 ( \32236 , \32235 , \9472 );
xor \U$31894 ( \32237 , \32234 , \32236 );
xor \U$31895 ( \32238 , \9153 , \9401 );
xor \U$31896 ( \32239 , \32238 , \9430 );
and \U$31897 ( \32240 , \11288 , \32239 );
xor \U$31898 ( \32241 , \9153 , \9401 );
xor \U$31899 ( \32242 , \32241 , \9430 );
and \U$31900 ( \32243 , \11292 , \32242 );
and \U$31901 ( \32244 , \11288 , \11292 );
or \U$31902 ( \32245 , \32240 , \32243 , \32244 );
xor \U$31903 ( \32246 , \11270 , \11274 );
and \U$31904 ( \32247 , \32246 , \11279 );
and \U$31905 ( \32248 , \11270 , \11274 );
nor \U$31906 ( \32249 , \32247 , \32248 );
xor \U$31907 ( \32250 , \32245 , \32249 );
xor \U$31908 ( \32251 , \8635 , \8637 );
xor \U$31909 ( \32252 , \32251 , \8648 );
xor \U$31910 ( \32253 , \9077 , \9084 );
xor \U$31911 ( \32254 , \32252 , \32253 );
xor \U$31912 ( \32255 , \32250 , \32254 );
xor \U$31913 ( \32256 , \32237 , \32255 );
not \U$31914 ( \32257 , \32256 );
or \U$31915 ( \32258 , \32228 , \32257 );
or \U$31916 ( \32259 , \32256 , \32227 );
nand \U$31917 ( \32260 , \32258 , \32259 );
xor \U$31918 ( \32261 , \32223 , \32260 );
and \U$31919 ( \32262 , \32222 , \32261 );
and \U$31920 ( \32263 , \32223 , \32260 );
nor \U$31921 ( \32264 , \32262 , \32263 );
not \U$31922 ( \32265 , \32256 );
nand \U$31923 ( \32266 , \32265 , \32227 );
xor \U$31924 ( \32267 , \9089 , \9475 );
xor \U$31925 ( \32268 , \32267 , \9482 );
not \U$31926 ( \32269 , \32268 );
not \U$31927 ( \32270 , \8651 );
not \U$31928 ( \32271 , \8947 );
or \U$31929 ( \32272 , \32270 , \32271 );
or \U$31930 ( \32273 , \8947 , \8651 );
nand \U$31931 ( \32274 , \32272 , \32273 );
not \U$31932 ( \32275 , \32274 );
not \U$31933 ( \32276 , \8633 );
and \U$31934 ( \32277 , \32275 , \32276 );
and \U$31935 ( \32278 , \32274 , \8633 );
nor \U$31936 ( \32279 , \32277 , \32278 );
xor \U$31937 ( \32280 , \32245 , \32249 );
and \U$31938 ( \32281 , \32280 , \32254 );
and \U$31939 ( \32282 , \32245 , \32249 );
or \U$31940 ( \32283 , \32281 , \32282 );
xor \U$31941 ( \32284 , \32279 , \32283 );
not \U$31942 ( \32285 , \32284 );
or \U$31943 ( \32286 , \32269 , \32285 );
or \U$31944 ( \32287 , \32284 , \32268 );
nand \U$31945 ( \32288 , \32286 , \32287 );
not \U$31946 ( \32289 , \32288 );
xor \U$31947 ( \32290 , \32234 , \32236 );
and \U$31948 ( \32291 , \32290 , \32255 );
and \U$31949 ( \32292 , \32234 , \32236 );
or \U$31950 ( \32293 , \32291 , \32292 );
not \U$31951 ( \32294 , \32293 );
and \U$31952 ( \32295 , \32289 , \32294 );
and \U$31953 ( \32296 , \32288 , \32293 );
nor \U$31954 ( \32297 , \32295 , \32296 );
xnor \U$31955 ( \32298 , \32266 , \32297 );
or \U$31956 ( \32299 , \32264 , \32298 );
or \U$31957 ( \32300 , \32266 , \32297 );
nand \U$31958 ( \32301 , \32299 , \32300 );
not \U$31959 ( \32302 , \32288 );
nor \U$31960 ( \32303 , \32302 , \32293 );
not \U$31961 ( \32304 , \32268 );
not \U$31962 ( \32305 , \32279 );
and \U$31963 ( \32306 , \32304 , \32305 );
and \U$31964 ( \32307 , \32268 , \32279 );
nor \U$31965 ( \32308 , \32307 , \32283 );
nor \U$31966 ( \32309 , \32306 , \32308 );
not \U$31967 ( \32310 , \32309 );
not \U$31968 ( \32311 , \9069 );
not \U$31969 ( \32312 , \9485 );
not \U$31970 ( \32313 , \9071 );
and \U$31971 ( \32314 , \32312 , \32313 );
and \U$31972 ( \32315 , \9485 , \9071 );
nor \U$31973 ( \32316 , \32314 , \32315 );
not \U$31974 ( \32317 , \32316 );
or \U$31975 ( \32318 , \32311 , \32317 );
or \U$31976 ( \32319 , \32316 , \9069 );
nand \U$31977 ( \32320 , \32318 , \32319 );
not \U$31978 ( \32321 , \32320 );
or \U$31979 ( \32322 , \32310 , \32321 );
or \U$31980 ( \32323 , \32320 , \32309 );
nand \U$31981 ( \32324 , \32322 , \32323 );
xor \U$31982 ( \32325 , \32303 , \32324 );
and \U$31983 ( \32326 , \32301 , \32325 );
and \U$31984 ( \32327 , \32303 , \32324 );
nor \U$31985 ( \32328 , \32326 , \32327 );
not \U$31986 ( \32329 , \32309 );
nand \U$31987 ( \32330 , \32329 , \32320 );
not \U$31988 ( \32331 , \9066 );
not \U$31989 ( \32332 , \9487 );
and \U$31990 ( \32333 , \32331 , \32332 );
and \U$31991 ( \32334 , \9066 , \9487 );
nor \U$31992 ( \32335 , \32333 , \32334 );
xnor \U$31993 ( \32336 , \32330 , \32335 );
or \U$31994 ( \32337 , \32328 , \32336 );
or \U$31995 ( \32338 , \32330 , \32335 );
nand \U$31996 ( \32339 , \32337 , \32338 );
and \U$31997 ( \32340 , \9490 , \32339 );
nor \U$31998 ( \32341 , \9489 , \32340 );
xnor \U$31999 ( \32342 , \9061 , \9053 );
or \U$32000 ( \32343 , \32341 , \32342 );
nand \U$32001 ( \32344 , \9063 , \32343 );
and \U$32002 ( \32345 , \9058 , \9060 );
not \U$32003 ( \32346 , \8330 );
not \U$32004 ( \32347 , \7965 );
or \U$32005 ( \32348 , \32346 , \32347 );
or \U$32006 ( \32349 , \7965 , \8330 );
nand \U$32007 ( \32350 , \32348 , \32349 );
xor \U$32008 ( \32351 , \32345 , \32350 );
and \U$32009 ( \32352 , \32344 , \32351 );
and \U$32010 ( \32353 , \32345 , \32350 );
nor \U$32011 ( \32354 , \32352 , \32353 );
or \U$32012 ( \32355 , \8333 , \32354 );
nand \U$32013 ( \32356 , \8332 , \32355 );
xor \U$32014 ( \32357 , \7248 , \7264 );
xor \U$32015 ( \32358 , \32357 , \7280 );
not \U$32016 ( \32359 , \7610 );
or \U$32017 ( \32360 , \7959 , \32359 );
and \U$32018 ( \32361 , \7959 , \32359 );
nor \U$32019 ( \32362 , \32361 , \7948 );
not \U$32020 ( \32363 , \32362 );
nand \U$32021 ( \32364 , \32360 , \32363 );
xor \U$32022 ( \32365 , \32358 , \32364 );
and \U$32023 ( \32366 , \32356 , \32365 );
and \U$32024 ( \32367 , \32358 , \32364 );
nor \U$32025 ( \32368 , \32366 , \32367 );
xnor \U$32026 ( \32369 , \7283 , \7308 );
or \U$32027 ( \32370 , \32368 , \32369 );
nand \U$32028 ( \32371 , \7310 , \32370 );
xor \U$32029 ( \32372 , \7293 , \7297 );
and \U$32030 ( \32373 , \32372 , \7306 );
and \U$32031 ( \32374 , \7293 , \7297 );
nor \U$32032 ( \32375 , \32373 , \32374 );
not \U$32033 ( \32376 , \32375 );
xor \U$32034 ( \32377 , \6349 , \6351 );
xor \U$32035 ( \32378 , \32377 , \6354 );
not \U$32036 ( \32379 , \32378 );
or \U$32037 ( \32380 , \32376 , \32379 );
or \U$32038 ( \32381 , \32378 , \32375 );
nand \U$32039 ( \32382 , \32380 , \32381 );
xor \U$32040 ( \32383 , \7288 , \7290 );
and \U$32041 ( \32384 , \32383 , \7307 );
and \U$32042 ( \32385 , \7288 , \7290 );
or \U$32043 ( \32386 , \32384 , \32385 );
xor \U$32044 ( \32387 , \32382 , \32386 );
and \U$32045 ( \32388 , \32371 , \32387 );
and \U$32046 ( \32389 , \32382 , \32386 );
nor \U$32047 ( \32390 , \32388 , \32389 );
xor \U$32048 ( \32391 , \6357 , \6359 );
not \U$32049 ( \32392 , \32391 );
not \U$32050 ( \32393 , \32375 );
nand \U$32051 ( \32394 , \32393 , \32378 );
not \U$32052 ( \32395 , \32394 );
and \U$32053 ( \32396 , \32392 , \32395 );
and \U$32054 ( \32397 , \32391 , \32394 );
nor \U$32055 ( \32398 , \32396 , \32397 );
or \U$32056 ( \32399 , \32390 , \32398 );
not \U$32057 ( \32400 , \32391 );
or \U$32058 ( \32401 , \32394 , \32400 );
nand \U$32059 ( \32402 , \32399 , \32401 );
and \U$32060 ( \32403 , \6362 , \32402 );
nor \U$32061 ( \32404 , \6361 , \32403 );
or \U$32062 ( \32405 , \6067 , \32404 );
nand \U$32063 ( \32406 , \6066 , \32405 );
not \U$32064 ( \32407 , \5778 );
nor \U$32065 ( \32408 , \32407 , \5527 );
not \U$32066 ( \32409 , \5514 );
not \U$32067 ( \32410 , \5256 );
or \U$32068 ( \32411 , \32409 , \32410 );
or \U$32069 ( \32412 , \5256 , \5514 );
nand \U$32070 ( \32413 , \32411 , \32412 );
xor \U$32071 ( \32414 , \32408 , \32413 );
and \U$32072 ( \32415 , \32406 , \32414 );
and \U$32073 ( \32416 , \32408 , \32413 );
nor \U$32074 ( \32417 , \32415 , \32416 );
or \U$32075 ( \32418 , \5517 , \32417 );
nand \U$32076 ( \32419 , \5516 , \32418 );
and \U$32077 ( \32420 , \5249 , \32419 );
nor \U$32078 ( \32421 , \5248 , \32420 );
xnor \U$32079 ( \32422 , \4147 , \4417 );
not \U$32080 ( \32423 , \32422 );
not \U$32081 ( \32424 , \4154 );
and \U$32082 ( \32425 , \32423 , \32424 );
and \U$32083 ( \32426 , \32422 , \4154 );
nor \U$32084 ( \32427 , \32425 , \32426 );
not \U$32085 ( \32428 , \32427 );
xor \U$32086 ( \32429 , \4176 , \4407 );
xor \U$32087 ( \32430 , \32429 , \4414 );
and \U$32088 ( \32431 , \4957 , \32430 );
xor \U$32089 ( \32432 , \4176 , \4407 );
xor \U$32090 ( \32433 , \32432 , \4414 );
and \U$32091 ( \32434 , \4961 , \32433 );
and \U$32092 ( \32435 , \4957 , \4961 );
or \U$32093 ( \32436 , \32431 , \32434 , \32435 );
not \U$32094 ( \32437 , \32436 );
and \U$32095 ( \32438 , \32428 , \32437 );
and \U$32096 ( \32439 , \32427 , \32436 );
nor \U$32097 ( \32440 , \32438 , \32439 );
nand \U$32098 ( \32441 , \4945 , \4963 );
xnor \U$32099 ( \32442 , \32440 , \32441 );
or \U$32100 ( \32443 , \32421 , \32442 );
or \U$32101 ( \32444 , \32441 , \32440 );
nand \U$32102 ( \32445 , \32443 , \32444 );
not \U$32103 ( \32446 , \32436 );
nor \U$32104 ( \32447 , \32446 , \32427 );
xor \U$32105 ( \32448 , \4419 , \4429 );
xor \U$32106 ( \32449 , \32447 , \32448 );
and \U$32107 ( \32450 , \32445 , \32449 );
and \U$32108 ( \32451 , \32447 , \32448 );
nor \U$32109 ( \32452 , \32450 , \32451 );
not \U$32110 ( \32453 , \32452 );
and \U$32111 ( \32454 , \4437 , \32453 );
nor \U$32112 ( \32455 , \4436 , \32454 );
and \U$32113 ( \32456 , \4145 , \32455 );
and \U$32114 ( \32457 , \4139 , \4144 );
nor \U$32115 ( \32458 , \32456 , \32457 );
and \U$32116 ( \32459 , \3862 , \32458 );
nor \U$32117 ( \32460 , \3861 , \32459 );
not \U$32118 ( \32461 , \3121 );
not \U$32119 ( \32462 , \2919 );
and \U$32120 ( \32463 , \32461 , \32462 );
and \U$32121 ( \32464 , \3121 , \2919 );
nor \U$32122 ( \32465 , \32463 , \32464 );
not \U$32123 ( \32466 , \32465 );
not \U$32124 ( \32467 , \2921 );
and \U$32125 ( \32468 , \32466 , \32467 );
and \U$32126 ( \32469 , \32465 , \2921 );
nor \U$32127 ( \32470 , \32468 , \32469 );
and \U$32128 ( \32471 , \3127 , \3580 );
not \U$32129 ( \32472 , \3127 );
not \U$32130 ( \32473 , \3580 );
and \U$32131 ( \32474 , \32472 , \32473 );
nor \U$32132 ( \32475 , \32474 , \3575 );
nor \U$32133 ( \32476 , \32471 , \32475 );
xnor \U$32134 ( \32477 , \32470 , \32476 );
or \U$32135 ( \32478 , \32460 , \32477 );
or \U$32136 ( \32479 , \32470 , \32476 );
nand \U$32137 ( \32480 , \32478 , \32479 );
and \U$32138 ( \32481 , \3125 , \32480 );
nor \U$32139 ( \32482 , \3124 , \32481 );
and \U$32140 ( \32483 , \2912 , \32482 );
and \U$32141 ( \32484 , \2848 , \2911 );
nor \U$32142 ( \32485 , \32483 , \32484 );
not \U$32143 ( \32486 , \2907 );
nor \U$32144 ( \32487 , \32486 , \2902 );
xor \U$32145 ( \32488 , \2855 , \2871 );
and \U$32146 ( \32489 , \32488 , \2901 );
and \U$32147 ( \32490 , \2855 , \2871 );
or \U$32148 ( \32491 , \32489 , \32490 );
not \U$32149 ( \32492 , \32491 );
xor \U$32150 ( \32493 , \2887 , \2892 );
and \U$32151 ( \32494 , \32493 , \2899 );
and \U$32152 ( \32495 , \2887 , \2892 );
or \U$32153 ( \32496 , \32494 , \32495 );
xor \U$32154 ( \32497 , \2859 , \2861 );
and \U$32155 ( \32498 , \32497 , \2870 );
and \U$32156 ( \32499 , \2859 , \2861 );
or \U$32157 ( \32500 , \32498 , \32499 );
xor \U$32158 ( \32501 , \32496 , \32500 );
xor \U$32159 ( \32502 , \1223 , \1348 );
xor \U$32160 ( \32503 , \32502 , \1442 );
xor \U$32161 ( \32504 , \32501 , \32503 );
not \U$32162 ( \32505 , \32504 );
xnor \U$32163 ( \32506 , \1533 , \1574 );
not \U$32164 ( \32507 , \32506 );
not \U$32165 ( \32508 , \1451 );
and \U$32166 ( \32509 , \32507 , \32508 );
and \U$32167 ( \32510 , \32506 , \1451 );
nor \U$32168 ( \32511 , \32509 , \32510 );
xor \U$32169 ( \32512 , \2880 , \2884 );
and \U$32170 ( \32513 , \32512 , \2900 );
and \U$32171 ( \32514 , \2880 , \2884 );
or \U$32172 ( \32515 , \32513 , \32514 );
xor \U$32173 ( \32516 , \32511 , \32515 );
not \U$32174 ( \32517 , \32516 );
or \U$32175 ( \32518 , \32505 , \32517 );
or \U$32176 ( \32519 , \32516 , \32504 );
nand \U$32177 ( \32520 , \32518 , \32519 );
not \U$32178 ( \32521 , \32520 );
or \U$32179 ( \32522 , \32492 , \32521 );
or \U$32180 ( \32523 , \32520 , \32491 );
nand \U$32181 ( \32524 , \32522 , \32523 );
xor \U$32182 ( \32525 , \32487 , \32524 );
and \U$32183 ( \32526 , \32485 , \32525 );
and \U$32184 ( \32527 , \32487 , \32524 );
nor \U$32185 ( \32528 , \32526 , \32527 );
not \U$32186 ( \32529 , \32491 );
nand \U$32187 ( \32530 , \32529 , \32520 );
xor \U$32188 ( \32531 , \1445 , \1576 );
xor \U$32189 ( \32532 , \32531 , \1684 );
not \U$32190 ( \32533 , \32532 );
xor \U$32191 ( \32534 , \32496 , \32500 );
and \U$32192 ( \32535 , \32534 , \32503 );
and \U$32193 ( \32536 , \32496 , \32500 );
or \U$32194 ( \32537 , \32535 , \32536 );
not \U$32195 ( \32538 , \32537 );
xor \U$32196 ( \32539 , \1705 , \1711 );
xor \U$32197 ( \32540 , \32539 , \1716 );
not \U$32198 ( \32541 , \32540 );
and \U$32199 ( \32542 , \32538 , \32541 );
and \U$32200 ( \32543 , \32537 , \32540 );
nor \U$32201 ( \32544 , \32542 , \32543 );
not \U$32202 ( \32545 , \32544 );
or \U$32203 ( \32546 , \32533 , \32545 );
or \U$32204 ( \32547 , \32544 , \32532 );
nand \U$32205 ( \32548 , \32546 , \32547 );
not \U$32206 ( \32549 , \32548 );
not \U$32207 ( \32550 , \32504 );
not \U$32208 ( \32551 , \32511 );
and \U$32209 ( \32552 , \32550 , \32551 );
and \U$32210 ( \32553 , \32504 , \32511 );
nor \U$32211 ( \32554 , \32553 , \32515 );
nor \U$32212 ( \32555 , \32552 , \32554 );
not \U$32213 ( \32556 , \32555 );
and \U$32214 ( \32557 , \32549 , \32556 );
and \U$32215 ( \32558 , \32548 , \32555 );
nor \U$32216 ( \32559 , \32557 , \32558 );
xnor \U$32217 ( \32560 , \32530 , \32559 );
or \U$32218 ( \32561 , \32528 , \32560 );
or \U$32219 ( \32562 , \32530 , \32559 );
nand \U$32220 ( \32563 , \32561 , \32562 );
not \U$32221 ( \32564 , \32548 );
nor \U$32222 ( \32565 , \32564 , \32555 );
and \U$32223 ( \32566 , \32532 , \32540 );
not \U$32224 ( \32567 , \32532 );
not \U$32225 ( \32568 , \32540 );
and \U$32226 ( \32569 , \32567 , \32568 );
nor \U$32227 ( \32570 , \32569 , \32537 );
nor \U$32228 ( \32571 , \32566 , \32570 );
not \U$32229 ( \32572 , \32571 );
xor \U$32230 ( \32573 , \1687 , \1694 );
xor \U$32231 ( \32574 , \32573 , \1820 );
not \U$32232 ( \32575 , \32574 );
or \U$32233 ( \32576 , \32572 , \32575 );
or \U$32234 ( \32577 , \32574 , \32571 );
nand \U$32235 ( \32578 , \32576 , \32577 );
xor \U$32236 ( \32579 , \32565 , \32578 );
and \U$32237 ( \32580 , \32563 , \32579 );
and \U$32238 ( \32581 , \32565 , \32578 );
nor \U$32239 ( \32582 , \32580 , \32581 );
not \U$32240 ( \32583 , \32571 );
nand \U$32241 ( \32584 , \32583 , \32574 );
not \U$32242 ( \32585 , \1957 );
not \U$32243 ( \32586 , \1823 );
and \U$32244 ( \32587 , \32585 , \32586 );
and \U$32245 ( \32588 , \1957 , \1823 );
nor \U$32246 ( \32589 , \32587 , \32588 );
xnor \U$32247 ( \32590 , \32584 , \32589 );
or \U$32248 ( \32591 , \32582 , \32590 );
or \U$32249 ( \32592 , \32584 , \32589 );
nand \U$32250 ( \32593 , \32591 , \32592 );
and \U$32251 ( \32594 , \2026 , \32593 );
nor \U$32252 ( \32595 , \2025 , \32594 );
not \U$32253 ( \32596 , \2013 );
nand \U$32254 ( \32597 , \32596 , \2020 );
xor \U$32255 ( \32598 , \1976 , \1992 );
and \U$32256 ( \32599 , \32598 , \2008 );
and \U$32257 ( \32600 , \1976 , \1992 );
or \U$32258 ( \32601 , \32599 , \32600 );
not \U$32259 ( \32602 , \32601 );
or \U$32260 ( \32603 , \2009 , \1960 );
not \U$32261 ( \32604 , \1960 );
not \U$32262 ( \32605 , \2009 );
or \U$32263 ( \32606 , \32604 , \32605 );
nand \U$32264 ( \32607 , \32606 , \1965 );
nand \U$32265 ( \32608 , \32603 , \32607 );
not \U$32266 ( \32609 , \32608 );
or \U$32267 ( \32610 , \32602 , \32609 );
or \U$32268 ( \32611 , \32608 , \32601 );
nand \U$32269 ( \32612 , \32610 , \32611 );
not \U$32270 ( \32613 , \32612 );
xor \U$32271 ( \32614 , \1997 , \1998 );
and \U$32272 ( \32615 , \32614 , \2007 );
and \U$32273 ( \32616 , \1997 , \1998 );
or \U$32274 ( \32617 , \32615 , \32616 );
xor \U$32275 ( \32618 , \1119 , \1139 );
xor \U$32276 ( \32619 , \32618 , \1168 );
xor \U$32277 ( \32620 , \32617 , \32619 );
xor \U$32278 ( \32621 , \1126 , \1128 );
xor \U$32279 ( \32622 , \32621 , \1136 );
and \U$32280 ( \32623 , \2003 , \32622 );
xor \U$32281 ( \32624 , \1126 , \1128 );
xor \U$32282 ( \32625 , \32624 , \1136 );
and \U$32283 ( \32626 , \2005 , \32625 );
and \U$32284 ( \32627 , \2003 , \2005 );
or \U$32285 ( \32628 , \32623 , \32626 , \32627 );
xor \U$32286 ( \32629 , \1980 , \1984 );
and \U$32287 ( \32630 , \32629 , \1991 );
and \U$32288 ( \32631 , \1980 , \1984 );
or \U$32289 ( \32632 , \32630 , \32631 );
xor \U$32290 ( \32633 , \32628 , \32632 );
xnor \U$32291 ( \32634 , \1091 , \1089 );
not \U$32292 ( \32635 , \32634 );
not \U$32293 ( \32636 , \1097 );
and \U$32294 ( \32637 , \32635 , \32636 );
and \U$32295 ( \32638 , \32634 , \1097 );
nor \U$32296 ( \32639 , \32637 , \32638 );
xor \U$32297 ( \32640 , \32633 , \32639 );
xor \U$32298 ( \32641 , \32620 , \32640 );
not \U$32299 ( \32642 , \32641 );
and \U$32300 ( \32643 , \32613 , \32642 );
and \U$32301 ( \32644 , \32612 , \32641 );
nor \U$32302 ( \32645 , \32643 , \32644 );
xnor \U$32303 ( \32646 , \32597 , \32645 );
or \U$32304 ( \32647 , \32595 , \32646 );
or \U$32305 ( \32648 , \32597 , \32645 );
nand \U$32306 ( \32649 , \32647 , \32648 );
xor \U$32307 ( \32650 , \32617 , \32619 );
and \U$32308 ( \32651 , \32650 , \32640 );
and \U$32309 ( \32652 , \32617 , \32619 );
or \U$32310 ( \32653 , \32651 , \32652 );
not \U$32311 ( \32654 , \32653 );
xor \U$32312 ( \32655 , \1099 , \1171 );
xor \U$32313 ( \32656 , \32655 , \1174 );
not \U$32314 ( \32657 , \32656 );
xor \U$32315 ( \32658 , \32628 , \32632 );
and \U$32316 ( \32659 , \32658 , \32639 );
and \U$32317 ( \32660 , \32628 , \32632 );
or \U$32318 ( \32661 , \32659 , \32660 );
not \U$32319 ( \32662 , \32661 );
xor \U$32320 ( \32663 , \740 , \749 );
xor \U$32321 ( \32664 , \32663 , \783 );
not \U$32322 ( \32665 , \32664 );
and \U$32323 ( \32666 , \32662 , \32665 );
and \U$32324 ( \32667 , \32661 , \32664 );
nor \U$32325 ( \32668 , \32666 , \32667 );
not \U$32326 ( \32669 , \32668 );
or \U$32327 ( \32670 , \32657 , \32669 );
or \U$32328 ( \32671 , \32668 , \32656 );
nand \U$32329 ( \32672 , \32670 , \32671 );
not \U$32330 ( \32673 , \32672 );
or \U$32331 ( \32674 , \32654 , \32673 );
or \U$32332 ( \32675 , \32653 , \32672 );
nand \U$32333 ( \32676 , \32674 , \32675 );
or \U$32334 ( \32677 , \32641 , \32601 );
not \U$32335 ( \32678 , \32601 );
not \U$32336 ( \32679 , \32641 );
or \U$32337 ( \32680 , \32678 , \32679 );
nand \U$32338 ( \32681 , \32680 , \32608 );
nand \U$32339 ( \32682 , \32677 , \32681 );
xor \U$32340 ( \32683 , \32676 , \32682 );
and \U$32341 ( \32684 , \32649 , \32683 );
and \U$32342 ( \32685 , \32676 , \32682 );
nor \U$32343 ( \32686 , \32684 , \32685 );
not \U$32344 ( \32687 , \32653 );
nand \U$32345 ( \32688 , \32687 , \32672 );
xor \U$32346 ( \32689 , \1177 , \1187 );
xor \U$32347 ( \32690 , \32689 , \1190 );
not \U$32348 ( \32691 , \32690 );
and \U$32349 ( \32692 , \32656 , \32664 );
not \U$32350 ( \32693 , \32656 );
not \U$32351 ( \32694 , \32664 );
and \U$32352 ( \32695 , \32693 , \32694 );
nor \U$32353 ( \32696 , \32695 , \32661 );
nor \U$32354 ( \32697 , \32692 , \32696 );
not \U$32355 ( \32698 , \32697 );
and \U$32356 ( \32699 , \32691 , \32698 );
and \U$32357 ( \32700 , \32690 , \32697 );
nor \U$32358 ( \32701 , \32699 , \32700 );
xnor \U$32359 ( \32702 , \32688 , \32701 );
or \U$32360 ( \32703 , \32686 , \32702 );
or \U$32361 ( \32704 , \32688 , \32701 );
nand \U$32362 ( \32705 , \32703 , \32704 );
not \U$32363 ( \32706 , \32690 );
nor \U$32364 ( \32707 , \32706 , \32697 );
not \U$32365 ( \32708 , \1193 );
not \U$32366 ( \32709 , \1078 );
or \U$32367 ( \32710 , \32708 , \32709 );
or \U$32368 ( \32711 , \1078 , \1193 );
nand \U$32369 ( \32712 , \32710 , \32711 );
xor \U$32370 ( \32713 , \32707 , \32712 );
and \U$32371 ( \32714 , \32705 , \32713 );
and \U$32372 ( \32715 , \32707 , \32712 );
nor \U$32373 ( \32716 , \32714 , \32715 );
or \U$32374 ( \32717 , \1196 , \32716 );
nand \U$32375 ( \32718 , \1195 , \32717 );
not \U$32376 ( \32719 , \32718 );
or \U$32377 ( \32720 , \1063 , \32719 );
or \U$32378 ( \32721 , \32718 , \1062 );
nand \U$32379 ( \32722 , \32720 , \32721 );
not \U$32380 ( \32723 , \32722 );
or \U$32381 ( \32724 , \803 , \32723 );
or \U$32382 ( \32725 , \32722 , \802 );
nand \U$32383 ( \32726 , \32724 , \32725 );
not \U$32384 ( \32727 , \32726 );
xor \U$32385 ( \32728 , \1023 , \1049 );
and \U$32386 ( \32729 , \32728 , \1058 );
and \U$32387 ( \32730 , \1023 , \1049 );
or \U$32388 ( \32731 , \32729 , \32730 );
not \U$32389 ( \32732 , \32731 );
not \U$32390 ( \32733 , \981 );
nor \U$32391 ( \32734 , \32733 , \1006 );
not \U$32392 ( \32735 , \32734 );
and \U$32393 ( \32736 , \32732 , \32735 );
and \U$32394 ( \32737 , \32731 , \32734 );
nor \U$32395 ( \32738 , \32736 , \32737 );
not \U$32396 ( \32739 , \32738 );
xor \U$32397 ( \32740 , \990 , \996 );
and \U$32398 ( \32741 , \32740 , \1005 );
and \U$32399 ( \32742 , \990 , \996 );
or \U$32400 ( \32743 , \32741 , \32742 );
not \U$32401 ( \32744 , \32743 );
not \U$32402 ( \32745 , \980 );
or \U$32403 ( \32746 , \32744 , \32745 );
or \U$32404 ( \32747 , \980 , \32743 );
nand \U$32405 ( \32748 , \32746 , \32747 );
not \U$32406 ( \32749 , \32748 );
and \U$32407 ( \32750 , \32739 , \32749 );
and \U$32408 ( \32751 , \32738 , \32748 );
nor \U$32409 ( \32752 , \32750 , \32751 );
not \U$32410 ( \32753 , \32752 );
and \U$32411 ( \32754 , \32727 , \32753 );
and \U$32412 ( \32755 , \32726 , \32752 );
nor \U$32413 ( \32756 , \32754 , \32755 );
not \U$32414 ( \32757 , \32756 );
not \U$32415 ( \32758 , \679 );
nand \U$32416 ( \32759 , \32758 , \646 );
not \U$32417 ( \32760 , \32759 );
not \U$32418 ( \32761 , \645 );
and \U$32419 ( \32762 , \32760 , \32761 );
and \U$32420 ( \32763 , \32759 , \645 );
nor \U$32421 ( \32764 , \32762 , \32763 );
not \U$32422 ( \32765 , \32764 );
or \U$32423 ( \32766 , \662 , \675 );
not \U$32424 ( \32767 , \675 );
not \U$32425 ( \32768 , \662 );
or \U$32426 ( \32769 , \32767 , \32768 );
nand \U$32427 ( \32770 , \32769 , \653 );
nand \U$32428 ( \32771 , \32766 , \32770 );
not \U$32429 ( \32772 , \32771 );
xor \U$32430 ( \32773 , \609 , \610 );
and \U$32431 ( \32774 , \32773 , \619 );
and \U$32432 ( \32775 , \609 , \610 );
or \U$32433 ( \32776 , \32774 , \32775 );
not \U$32434 ( \32777 , \32776 );
or \U$32435 ( \32778 , \32772 , \32777 );
or \U$32436 ( \32779 , \32776 , \32771 );
nand \U$32437 ( \32780 , \32778 , \32779 );
not \U$32438 ( \32781 , \32780 );
and \U$32439 ( \32782 , \32765 , \32781 );
and \U$32440 ( \32783 , \32764 , \32780 );
nor \U$32441 ( \32784 , \32782 , \32783 );
not \U$32442 ( \32785 , \32784 );
and \U$32443 ( \32786 , \354 , RI986de28_4);
and \U$32444 ( \32787 , RI986dd38_2, \352 );
nor \U$32445 ( \32788 , \32786 , \32787 );
and \U$32446 ( \32789 , \416 , RI986e008_8);
and \U$32447 ( \32790 , RI986df18_6, \414 );
nor \U$32448 ( \32791 , \32789 , \32790 );
xor \U$32449 ( \32792 , \32788 , \32791 );
not \U$32450 ( \32793 , \32792 );
or \U$32451 ( \32794 , \630 , \683 );
not \U$32452 ( \32795 , \683 );
not \U$32453 ( \32796 , \630 );
or \U$32454 ( \32797 , \32795 , \32796 );
nand \U$32455 ( \32798 , \32797 , \587 );
nand \U$32456 ( \32799 , \32794 , \32798 );
not \U$32457 ( \32800 , \32799 );
xor \U$32458 ( \32801 , \602 , \620 );
and \U$32459 ( \32802 , \32801 , \629 );
and \U$32460 ( \32803 , \602 , \620 );
or \U$32461 ( \32804 , \32802 , \32803 );
not \U$32462 ( \32805 , \32804 );
and \U$32463 ( \32806 , \32800 , \32805 );
and \U$32464 ( \32807 , \32799 , \32804 );
nor \U$32465 ( \32808 , \32806 , \32807 );
not \U$32466 ( \32809 , \32808 );
or \U$32467 ( \32810 , \32793 , \32809 );
or \U$32468 ( \32811 , \32808 , \32792 );
nand \U$32469 ( \32812 , \32810 , \32811 );
not \U$32470 ( \32813 , \32812 );
or \U$32471 ( \32814 , \32785 , \32813 );
or \U$32472 ( \32815 , \32812 , \32784 );
nand \U$32473 ( \32816 , \32814 , \32815 );
not \U$32474 ( \32817 , \32816 );
and \U$32475 ( \32818 , \32757 , \32817 );
and \U$32476 ( \32819 , \32756 , \32816 );
nor \U$32477 ( \32820 , \32818 , \32819 );
not \U$32478 ( \32821 , \32820 );
or \U$32479 ( \32822 , \1030 , \1045 );
not \U$32480 ( \32823 , \1045 );
not \U$32481 ( \32824 , \1030 );
or \U$32482 ( \32825 , \32823 , \32824 );
nand \U$32483 ( \32826 , \32825 , \1039 );
nand \U$32484 ( \32827 , \32822 , \32826 );
not \U$32485 ( \32828 , \32827 );
nand \U$32486 ( \32829 , RI986f688_56, RI9871fc8_144);
not \U$32487 ( \32830 , \32829 );
and \U$32488 ( \32831 , \32828 , \32830 );
and \U$32489 ( \32832 , \32827 , \32829 );
nor \U$32490 ( \32833 , \32831 , \32832 );
not \U$32491 ( \32834 , \32833 );
nand \U$32492 ( \32835 , RI986e3c8_16, \776 );
and \U$32493 ( \32836 , \32835 , \474 );
not \U$32494 ( \32837 , \32835 );
and \U$32495 ( \32838 , \32837 , \451 );
nor \U$32496 ( \32839 , \32836 , \32838 );
not \U$32497 ( \32840 , \32839 );
and \U$32498 ( \32841 , \438 , RI986e0f8_10);
and \U$32499 ( \32842 , RI986e2d8_14, \436 );
nor \U$32500 ( \32843 , \32841 , \32842 );
and \U$32501 ( \32844 , \32843 , \443 );
not \U$32502 ( \32845 , \32843 );
and \U$32503 ( \32846 , \32845 , \444 );
nor \U$32504 ( \32847 , \32844 , \32846 );
not \U$32505 ( \32848 , \32847 );
or \U$32506 ( \32849 , \32840 , \32848 );
or \U$32507 ( \32850 , \32847 , \32839 );
nand \U$32508 ( \32851 , \32849 , \32850 );
not \U$32509 ( \32852 , \32851 );
and \U$32510 ( \32853 , \465 , RI986dd38_2);
and \U$32511 ( \32854 , RI986e1e8_12, \463 );
nor \U$32512 ( \32855 , \32853 , \32854 );
not \U$32513 ( \32856 , \32855 );
not \U$32514 ( \32857 , \454 );
and \U$32515 ( \32858 , \32856 , \32857 );
and \U$32516 ( \32859 , \32855 , \454 );
nor \U$32517 ( \32860 , \32858 , \32859 );
not \U$32518 ( \32861 , \32860 );
and \U$32519 ( \32862 , \32852 , \32861 );
and \U$32520 ( \32863 , \32851 , \32860 );
nor \U$32521 ( \32864 , \32862 , \32863 );
and \U$32522 ( \32865 , \376 , RI986df18_6);
and \U$32523 ( \32866 , RI986de28_4, \374 );
nor \U$32524 ( \32867 , \32865 , \32866 );
not \U$32525 ( \32868 , \32867 );
not \U$32526 ( \32869 , \367 );
and \U$32527 ( \32870 , \32868 , \32869 );
and \U$32528 ( \32871 , \32867 , \367 );
nor \U$32529 ( \32872 , \32870 , \32871 );
not \U$32530 ( \32873 , \32872 );
not \U$32531 ( \32874 , \487 );
and \U$32532 ( \32875 , \395 , RI986f688_56);
and \U$32533 ( \32876 , RI986e008_8, \393 );
nor \U$32534 ( \32877 , \32875 , \32876 );
not \U$32535 ( \32878 , \32877 );
or \U$32536 ( \32879 , \32874 , \32878 );
or \U$32537 ( \32880 , \32877 , \386 );
nand \U$32538 ( \32881 , \32879 , \32880 );
not \U$32539 ( \32882 , \32881 );
or \U$32540 ( \32883 , \32873 , \32882 );
or \U$32541 ( \32884 , \32872 , \32881 );
nand \U$32542 ( \32885 , \32883 , \32884 );
not \U$32543 ( \32886 , \32885 );
and \U$32544 ( \32887 , \354 , RI986f3b8_50);
and \U$32545 ( \32888 , RI986f598_54, \352 );
nor \U$32546 ( \32889 , \32887 , \32888 );
not \U$32547 ( \32890 , \32889 );
not \U$32548 ( \32891 , \345 );
and \U$32549 ( \32892 , \32890 , \32891 );
and \U$32550 ( \32893 , \32889 , \361 );
nor \U$32551 ( \32894 , \32892 , \32893 );
not \U$32552 ( \32895 , \32894 );
and \U$32553 ( \32896 , \32886 , \32895 );
and \U$32554 ( \32897 , \32885 , \32894 );
nor \U$32555 ( \32898 , \32896 , \32897 );
or \U$32556 ( \32899 , \32864 , \32898 );
not \U$32557 ( \32900 , \32898 );
not \U$32558 ( \32901 , \32864 );
or \U$32559 ( \32902 , \32900 , \32901 );
and \U$32560 ( \32903 , \416 , RI986f958_62);
and \U$32561 ( \32904 , RI986f4a8_52, \414 );
nor \U$32562 ( \32905 , \32903 , \32904 );
and \U$32563 ( \32906 , \32905 , \421 );
not \U$32564 ( \32907 , \32905 );
and \U$32565 ( \32908 , \32907 , \422 );
nor \U$32566 ( \32909 , \32906 , \32908 );
nand \U$32567 ( \32910 , RI986fa48_64, RI9871fc8_144);
or \U$32568 ( \32911 , \32909 , \32910 );
nand \U$32569 ( \32912 , \32910 , \32909 );
nand \U$32570 ( \32913 , \32911 , \32912 );
nand \U$32571 ( \32914 , \32902 , \32913 );
nand \U$32572 ( \32915 , \32899 , \32914 );
and \U$32573 ( \32916 , \354 , RI986f4a8_52);
and \U$32574 ( \32917 , RI986f3b8_50, \352 );
nor \U$32575 ( \32918 , \32916 , \32917 );
not \U$32576 ( \32919 , \32918 );
not \U$32577 ( \32920 , \361 );
and \U$32578 ( \32921 , \32919 , \32920 );
and \U$32579 ( \32922 , \32918 , \345 );
nor \U$32580 ( \32923 , \32921 , \32922 );
nand \U$32581 ( \32924 , RI986f778_58, RI9871fc8_144);
xor \U$32582 ( \32925 , \32923 , \32924 );
and \U$32583 ( \32926 , \416 , RI986fa48_64);
and \U$32584 ( \32927 , RI986f958_62, \414 );
nor \U$32585 ( \32928 , \32926 , \32927 );
and \U$32586 ( \32929 , \32928 , \421 );
not \U$32587 ( \32930 , \32928 );
and \U$32588 ( \32931 , \32930 , \422 );
nor \U$32589 ( \32932 , \32929 , \32931 );
and \U$32590 ( \32933 , \32925 , \32932 );
and \U$32591 ( \32934 , \32923 , \32924 );
or \U$32592 ( \32935 , \32933 , \32934 );
and \U$32593 ( \32936 , \776 , RI986e2d8_14);
and \U$32594 ( \32937 , RI986e3c8_16, \774 );
nor \U$32595 ( \32938 , \32936 , \32937 );
and \U$32596 ( \32939 , \32938 , \451 );
not \U$32597 ( \32940 , \32938 );
and \U$32598 ( \32941 , \32940 , \474 );
nor \U$32599 ( \32942 , \32939 , \32941 );
xor \U$32600 ( \32943 , \32942 , \1301 );
and \U$32601 ( \32944 , \438 , RI986e1e8_12);
and \U$32602 ( \32945 , RI986e0f8_10, \436 );
nor \U$32603 ( \32946 , \32944 , \32945 );
and \U$32604 ( \32947 , \32946 , \443 );
not \U$32605 ( \32948 , \32946 );
and \U$32606 ( \32949 , \32948 , \444 );
nor \U$32607 ( \32950 , \32947 , \32949 );
and \U$32608 ( \32951 , \32943 , \32950 );
and \U$32609 ( \32952 , \32942 , \1301 );
or \U$32610 ( \32953 , \32951 , \32952 );
xor \U$32611 ( \32954 , \32935 , \32953 );
and \U$32612 ( \32955 , \395 , RI986f598_54);
and \U$32613 ( \32956 , RI986f688_56, \393 );
nor \U$32614 ( \32957 , \32955 , \32956 );
not \U$32615 ( \32958 , \32957 );
not \U$32616 ( \32959 , \487 );
and \U$32617 ( \32960 , \32958 , \32959 );
and \U$32618 ( \32961 , \32957 , \386 );
nor \U$32619 ( \32962 , \32960 , \32961 );
and \U$32620 ( \32963 , \465 , RI986de28_4);
and \U$32621 ( \32964 , RI986dd38_2, \463 );
nor \U$32622 ( \32965 , \32963 , \32964 );
not \U$32623 ( \32966 , \32965 );
not \U$32624 ( \32967 , \456 );
and \U$32625 ( \32968 , \32966 , \32967 );
and \U$32626 ( \32969 , \32965 , \454 );
nor \U$32627 ( \32970 , \32968 , \32969 );
xor \U$32628 ( \32971 , \32962 , \32970 );
and \U$32629 ( \32972 , \376 , RI986e008_8);
and \U$32630 ( \32973 , RI986df18_6, \374 );
nor \U$32631 ( \32974 , \32972 , \32973 );
not \U$32632 ( \32975 , \32974 );
not \U$32633 ( \32976 , \365 );
and \U$32634 ( \32977 , \32975 , \32976 );
and \U$32635 ( \32978 , \32974 , \367 );
nor \U$32636 ( \32979 , \32977 , \32978 );
and \U$32637 ( \32980 , \32971 , \32979 );
and \U$32638 ( \32981 , \32962 , \32970 );
or \U$32639 ( \32982 , \32980 , \32981 );
and \U$32640 ( \32983 , \32954 , \32982 );
and \U$32641 ( \32984 , \32935 , \32953 );
nor \U$32642 ( \32985 , \32983 , \32984 );
xor \U$32643 ( \32986 , \32915 , \32985 );
xor \U$32644 ( \32987 , \894 , \474 );
xor \U$32645 ( \32988 , \32987 , \903 );
xor \U$32646 ( \32989 , \909 , \916 );
xor \U$32647 ( \32990 , \867 , \875 );
xor \U$32648 ( \32991 , \32990 , \884 );
xor \U$32649 ( \32992 , \32989 , \32991 );
xor \U$32650 ( \32993 , \32988 , \32992 );
and \U$32651 ( \32994 , \32986 , \32993 );
and \U$32652 ( \32995 , \32915 , \32985 );
or \U$32653 ( \32996 , \32994 , \32995 );
xor \U$32654 ( \32997 , \887 , \906 );
xor \U$32655 ( \32998 , \32997 , \917 );
xor \U$32656 ( \32999 , \32996 , \32998 );
xor \U$32657 ( \33000 , \894 , \474 );
xor \U$32658 ( \33001 , \33000 , \903 );
and \U$32659 ( \33002 , \32989 , \33001 );
xor \U$32660 ( \33003 , \894 , \474 );
xor \U$32661 ( \33004 , \33003 , \903 );
and \U$32662 ( \33005 , \32991 , \33004 );
and \U$32663 ( \33006 , \32989 , \32991 );
or \U$32664 ( \33007 , \33002 , \33005 , \33006 );
or \U$32665 ( \33008 , \32872 , \32894 );
not \U$32666 ( \33009 , \32894 );
not \U$32667 ( \33010 , \32872 );
or \U$32668 ( \33011 , \33009 , \33010 );
nand \U$32669 ( \33012 , \33011 , \32881 );
nand \U$32670 ( \33013 , \33008 , \33012 );
xor \U$32671 ( \33014 , \33013 , \32912 );
or \U$32672 ( \33015 , \32847 , \32860 );
not \U$32673 ( \33016 , \32860 );
not \U$32674 ( \33017 , \32847 );
or \U$32675 ( \33018 , \33016 , \33017 );
nand \U$32676 ( \33019 , \33018 , \32839 );
nand \U$32677 ( \33020 , \33015 , \33019 );
and \U$32678 ( \33021 , \33014 , \33020 );
and \U$32679 ( \33022 , \33013 , \32912 );
or \U$32680 ( \33023 , \33021 , \33022 );
xor \U$32681 ( \33024 , \33007 , \33023 );
not \U$32682 ( \33025 , \828 );
xnor \U$32683 ( \33026 , \826 , \857 );
not \U$32684 ( \33027 , \33026 );
or \U$32685 ( \33028 , \33025 , \33027 );
or \U$32686 ( \33029 , \33026 , \828 );
nand \U$32687 ( \33030 , \33028 , \33029 );
xor \U$32688 ( \33031 , \33024 , \33030 );
and \U$32689 ( \33032 , \32999 , \33031 );
and \U$32690 ( \33033 , \32996 , \32998 );
or \U$32691 ( \33034 , \33032 , \33033 );
not \U$32692 ( \33035 , \33034 );
xor \U$32693 ( \33036 , \33007 , \33023 );
and \U$32694 ( \33037 , \33036 , \33030 );
and \U$32695 ( \33038 , \33007 , \33023 );
nor \U$32696 ( \33039 , \33037 , \33038 );
xor \U$32697 ( \33040 , \1015 , \828 );
xor \U$32698 ( \33041 , \33040 , \1020 );
xor \U$32699 ( \33042 , \33039 , \33041 );
xor \U$32700 ( \33043 , \859 , \920 );
xor \U$32701 ( \33044 , \33043 , \967 );
xor \U$32702 ( \33045 , \33042 , \33044 );
not \U$32703 ( \33046 , \33045 );
or \U$32704 ( \33047 , \33035 , \33046 );
or \U$32705 ( \33048 , \33045 , \33034 );
nand \U$32706 ( \33049 , \33047 , \33048 );
xor \U$32707 ( \33050 , \32996 , \32998 );
xor \U$32708 ( \33051 , \33050 , \33031 );
not \U$32709 ( \33052 , \33051 );
xor \U$32710 ( \33053 , \32915 , \32985 );
xor \U$32711 ( \33054 , \33053 , \32993 );
xor \U$32712 ( \33055 , \33013 , \32912 );
xor \U$32713 ( \33056 , \33055 , \33020 );
and \U$32714 ( \33057 , \33054 , \33056 );
not \U$32715 ( \33058 , \33054 );
not \U$32716 ( \33059 , \33056 );
and \U$32717 ( \33060 , \33058 , \33059 );
xor \U$32718 ( \33061 , \32923 , \32924 );
xor \U$32719 ( \33062 , \33061 , \32932 );
xor \U$32720 ( \33063 , \32942 , \1301 );
xor \U$32721 ( \33064 , \33063 , \32950 );
and \U$32722 ( \33065 , \33062 , \33064 );
xor \U$32723 ( \33066 , \32962 , \32970 );
xor \U$32724 ( \33067 , \33066 , \32979 );
xor \U$32725 ( \33068 , \32942 , \1301 );
xor \U$32726 ( \33069 , \33068 , \32950 );
and \U$32727 ( \33070 , \33067 , \33069 );
and \U$32728 ( \33071 , \33062 , \33067 );
or \U$32729 ( \33072 , \33065 , \33070 , \33071 );
and \U$32730 ( \33073 , \376 , RI986f688_56);
and \U$32731 ( \33074 , RI986e008_8, \374 );
nor \U$32732 ( \33075 , \33073 , \33074 );
not \U$32733 ( \33076 , \33075 );
not \U$32734 ( \33077 , \367 );
and \U$32735 ( \33078 , \33076 , \33077 );
and \U$32736 ( \33079 , \33075 , \367 );
nor \U$32737 ( \33080 , \33078 , \33079 );
and \U$32738 ( \33081 , \465 , RI986df18_6);
and \U$32739 ( \33082 , RI986de28_4, \463 );
nor \U$32740 ( \33083 , \33081 , \33082 );
not \U$32741 ( \33084 , \33083 );
not \U$32742 ( \33085 , \454 );
and \U$32743 ( \33086 , \33084 , \33085 );
and \U$32744 ( \33087 , \33083 , \456 );
nor \U$32745 ( \33088 , \33086 , \33087 );
xor \U$32746 ( \33089 , \33080 , \33088 );
and \U$32747 ( \33090 , \395 , RI986f3b8_50);
and \U$32748 ( \33091 , RI986f598_54, \393 );
nor \U$32749 ( \33092 , \33090 , \33091 );
not \U$32750 ( \33093 , \33092 );
not \U$32751 ( \33094 , \386 );
and \U$32752 ( \33095 , \33093 , \33094 );
and \U$32753 ( \33096 , \33092 , \487 );
nor \U$32754 ( \33097 , \33095 , \33096 );
and \U$32755 ( \33098 , \33089 , \33097 );
and \U$32756 ( \33099 , \33080 , \33088 );
or \U$32757 ( \33100 , \33098 , \33099 );
and \U$32758 ( \33101 , \416 , RI986f778_58);
and \U$32759 ( \33102 , RI986fa48_64, \414 );
nor \U$32760 ( \33103 , \33101 , \33102 );
and \U$32761 ( \33104 , \33103 , \421 );
not \U$32762 ( \33105 , \33103 );
and \U$32763 ( \33106 , \33105 , \422 );
nor \U$32764 ( \33107 , \33104 , \33106 );
nand \U$32765 ( \33108 , RI986f868_60, RI9871fc8_144);
xor \U$32766 ( \33109 , \33107 , \33108 );
and \U$32767 ( \33110 , \354 , RI986f958_62);
and \U$32768 ( \33111 , RI986f4a8_52, \352 );
nor \U$32769 ( \33112 , \33110 , \33111 );
not \U$32770 ( \33113 , \33112 );
not \U$32771 ( \33114 , \361 );
and \U$32772 ( \33115 , \33113 , \33114 );
and \U$32773 ( \33116 , \33112 , \345 );
nor \U$32774 ( \33117 , \33115 , \33116 );
and \U$32775 ( \33118 , \33109 , \33117 );
and \U$32776 ( \33119 , \33107 , \33108 );
or \U$32777 ( \33120 , \33118 , \33119 );
xor \U$32778 ( \33121 , \33100 , \33120 );
and \U$32779 ( \33122 , \776 , RI986e0f8_10);
and \U$32780 ( \33123 , RI986e2d8_14, \774 );
nor \U$32781 ( \33124 , \33122 , \33123 );
and \U$32782 ( \33125 , \33124 , \451 );
not \U$32783 ( \33126 , \33124 );
and \U$32784 ( \33127 , \33126 , \474 );
nor \U$32785 ( \33128 , \33125 , \33127 );
nand \U$32786 ( \33129 , RI986e3c8_16, \1293 );
not \U$32787 ( \33130 , \33129 );
not \U$32788 ( \33131 , \1301 );
and \U$32789 ( \33132 , \33130 , \33131 );
and \U$32790 ( \33133 , \33129 , \1301 );
nor \U$32791 ( \33134 , \33132 , \33133 );
xor \U$32792 ( \33135 , \33128 , \33134 );
and \U$32793 ( \33136 , \438 , RI986dd38_2);
and \U$32794 ( \33137 , RI986e1e8_12, \436 );
nor \U$32795 ( \33138 , \33136 , \33137 );
and \U$32796 ( \33139 , \33138 , \443 );
not \U$32797 ( \33140 , \33138 );
and \U$32798 ( \33141 , \33140 , \444 );
nor \U$32799 ( \33142 , \33139 , \33141 );
and \U$32800 ( \33143 , \33135 , \33142 );
and \U$32801 ( \33144 , \33128 , \33134 );
or \U$32802 ( \33145 , \33143 , \33144 );
and \U$32803 ( \33146 , \33121 , \33145 );
and \U$32804 ( \33147 , \33100 , \33120 );
or \U$32805 ( \33148 , \33146 , \33147 );
xor \U$32806 ( \33149 , \33072 , \33148 );
xnor \U$32807 ( \33150 , \32898 , \32864 );
not \U$32808 ( \33151 , \33150 );
not \U$32809 ( \33152 , \32913 );
and \U$32810 ( \33153 , \33151 , \33152 );
and \U$32811 ( \33154 , \33150 , \32913 );
nor \U$32812 ( \33155 , \33153 , \33154 );
and \U$32813 ( \33156 , \33149 , \33155 );
and \U$32814 ( \33157 , \33072 , \33148 );
or \U$32815 ( \33158 , \33156 , \33157 );
nor \U$32816 ( \33159 , \33060 , \33158 );
nor \U$32817 ( \33160 , \33057 , \33159 );
nor \U$32818 ( \33161 , \33052 , \33160 );
and \U$32819 ( \33162 , \33049 , \33161 );
xor \U$32820 ( \33163 , \33161 , \33049 );
and \U$32821 ( \33164 , \416 , RI986f868_60);
and \U$32822 ( \33165 , RI986f778_58, \414 );
nor \U$32823 ( \33166 , \33164 , \33165 );
and \U$32824 ( \33167 , \33166 , \421 );
not \U$32825 ( \33168 , \33166 );
and \U$32826 ( \33169 , \33168 , \422 );
nor \U$32827 ( \33170 , \33167 , \33169 );
and \U$32828 ( \33171 , \395 , RI986f4a8_52);
and \U$32829 ( \33172 , RI986f3b8_50, \393 );
nor \U$32830 ( \33173 , \33171 , \33172 );
not \U$32831 ( \33174 , \33173 );
not \U$32832 ( \33175 , \487 );
and \U$32833 ( \33176 , \33174 , \33175 );
and \U$32834 ( \33177 , \33173 , \487 );
nor \U$32835 ( \33178 , \33176 , \33177 );
xor \U$32836 ( \33179 , \33170 , \33178 );
and \U$32837 ( \33180 , \354 , RI986fa48_64);
and \U$32838 ( \33181 , RI986f958_62, \352 );
nor \U$32839 ( \33182 , \33180 , \33181 );
not \U$32840 ( \33183 , \33182 );
not \U$32841 ( \33184 , \361 );
and \U$32842 ( \33185 , \33183 , \33184 );
and \U$32843 ( \33186 , \33182 , \361 );
nor \U$32844 ( \33187 , \33185 , \33186 );
and \U$32845 ( \33188 , \33179 , \33187 );
and \U$32846 ( \33189 , \33170 , \33178 );
or \U$32847 ( \33190 , \33188 , \33189 );
not \U$32848 ( \33191 , \1301 );
and \U$32849 ( \33192 , \1293 , RI986e2d8_14);
and \U$32850 ( \33193 , RI986e3c8_16, \1291 );
nor \U$32851 ( \33194 , \33192 , \33193 );
not \U$32852 ( \33195 , \33194 );
or \U$32853 ( \33196 , \33191 , \33195 );
or \U$32854 ( \33197 , \33194 , \1128 );
nand \U$32855 ( \33198 , \33196 , \33197 );
not \U$32856 ( \33199 , \33198 );
nand \U$32857 ( \33200 , \33199 , \1337 );
and \U$32858 ( \33201 , \776 , RI986e1e8_12);
and \U$32859 ( \33202 , RI986e0f8_10, \774 );
nor \U$32860 ( \33203 , \33201 , \33202 );
and \U$32861 ( \33204 , \33203 , \474 );
not \U$32862 ( \33205 , \33203 );
and \U$32863 ( \33206 , \33205 , \451 );
nor \U$32864 ( \33207 , \33204 , \33206 );
and \U$32865 ( \33208 , \33200 , \33207 );
and \U$32866 ( \33209 , \1336 , \33198 );
nor \U$32867 ( \33210 , \33208 , \33209 );
xor \U$32868 ( \33211 , \33190 , \33210 );
and \U$32869 ( \33212 , \376 , RI986f598_54);
and \U$32870 ( \33213 , RI986f688_56, \374 );
nor \U$32871 ( \33214 , \33212 , \33213 );
not \U$32872 ( \33215 , \33214 );
not \U$32873 ( \33216 , \367 );
and \U$32874 ( \33217 , \33215 , \33216 );
and \U$32875 ( \33218 , \33214 , \365 );
nor \U$32876 ( \33219 , \33217 , \33218 );
and \U$32877 ( \33220 , \438 , RI986de28_4);
and \U$32878 ( \33221 , RI986dd38_2, \436 );
nor \U$32879 ( \33222 , \33220 , \33221 );
and \U$32880 ( \33223 , \33222 , \443 );
not \U$32881 ( \33224 , \33222 );
and \U$32882 ( \33225 , \33224 , \444 );
nor \U$32883 ( \33226 , \33223 , \33225 );
xor \U$32884 ( \33227 , \33219 , \33226 );
and \U$32885 ( \33228 , \465 , RI986e008_8);
and \U$32886 ( \33229 , RI986df18_6, \463 );
nor \U$32887 ( \33230 , \33228 , \33229 );
not \U$32888 ( \33231 , \33230 );
not \U$32889 ( \33232 , \456 );
and \U$32890 ( \33233 , \33231 , \33232 );
and \U$32891 ( \33234 , \33230 , \456 );
nor \U$32892 ( \33235 , \33233 , \33234 );
and \U$32893 ( \33236 , \33227 , \33235 );
and \U$32894 ( \33237 , \33219 , \33226 );
or \U$32895 ( \33238 , \33236 , \33237 );
xor \U$32896 ( \33239 , \33211 , \33238 );
not \U$32897 ( \33240 , \33239 );
xor \U$32898 ( \33241 , \33128 , \33134 );
xor \U$32899 ( \33242 , \33241 , \33142 );
not \U$32900 ( \33243 , \33242 );
and \U$32901 ( \33244 , \776 , RI986dd38_2);
and \U$32902 ( \33245 , RI986e1e8_12, \774 );
nor \U$32903 ( \33246 , \33244 , \33245 );
and \U$32904 ( \33247 , \33246 , \474 );
not \U$32905 ( \33248 , \33246 );
and \U$32906 ( \33249 , \33248 , \451 );
nor \U$32907 ( \33250 , \33247 , \33249 );
nand \U$32908 ( \33251 , RI986e3c8_16, \1329 );
and \U$32909 ( \33252 , \33251 , \1336 );
not \U$32910 ( \33253 , \33251 );
and \U$32911 ( \33254 , \33253 , \1337 );
nor \U$32912 ( \33255 , \33252 , \33254 );
xor \U$32913 ( \33256 , \33250 , \33255 );
not \U$32914 ( \33257 , \1301 );
and \U$32915 ( \33258 , \1293 , RI986e0f8_10);
and \U$32916 ( \33259 , RI986e2d8_14, \1291 );
nor \U$32917 ( \33260 , \33258 , \33259 );
not \U$32918 ( \33261 , \33260 );
or \U$32919 ( \33262 , \33257 , \33261 );
or \U$32920 ( \33263 , \33260 , \1301 );
nand \U$32921 ( \33264 , \33262 , \33263 );
and \U$32922 ( \33265 , \33256 , \33264 );
and \U$32923 ( \33266 , \33250 , \33255 );
or \U$32924 ( \33267 , \33265 , \33266 );
not \U$32925 ( \33268 , \456 );
and \U$32926 ( \33269 , \465 , RI986f688_56);
and \U$32927 ( \33270 , RI986e008_8, \463 );
nor \U$32928 ( \33271 , \33269 , \33270 );
not \U$32929 ( \33272 , \33271 );
or \U$32930 ( \33273 , \33268 , \33272 );
or \U$32931 ( \33274 , \33271 , \456 );
nand \U$32932 ( \33275 , \33273 , \33274 );
and \U$32933 ( \33276 , \438 , RI986df18_6);
and \U$32934 ( \33277 , RI986de28_4, \436 );
nor \U$32935 ( \33278 , \33276 , \33277 );
and \U$32936 ( \33279 , \33278 , \444 );
not \U$32937 ( \33280 , \33278 );
and \U$32938 ( \33281 , \33280 , \443 );
nor \U$32939 ( \33282 , \33279 , \33281 );
xor \U$32940 ( \33283 , \33275 , \33282 );
not \U$32941 ( \33284 , \365 );
and \U$32942 ( \33285 , \376 , RI986f3b8_50);
and \U$32943 ( \33286 , RI986f598_54, \374 );
nor \U$32944 ( \33287 , \33285 , \33286 );
not \U$32945 ( \33288 , \33287 );
or \U$32946 ( \33289 , \33284 , \33288 );
or \U$32947 ( \33290 , \33287 , \365 );
nand \U$32948 ( \33291 , \33289 , \33290 );
and \U$32949 ( \33292 , \33283 , \33291 );
and \U$32950 ( \33293 , \33275 , \33282 );
or \U$32951 ( \33294 , \33292 , \33293 );
xor \U$32952 ( \33295 , \33267 , \33294 );
and \U$32953 ( \33296 , \395 , RI986f958_62);
and \U$32954 ( \33297 , RI986f4a8_52, \393 );
nor \U$32955 ( \33298 , \33296 , \33297 );
not \U$32956 ( \33299 , \33298 );
not \U$32957 ( \33300 , \386 );
and \U$32958 ( \33301 , \33299 , \33300 );
and \U$32959 ( \33302 , \33298 , \487 );
nor \U$32960 ( \33303 , \33301 , \33302 );
and \U$32961 ( \33304 , \354 , RI986f778_58);
and \U$32962 ( \33305 , RI986fa48_64, \352 );
nor \U$32963 ( \33306 , \33304 , \33305 );
not \U$32964 ( \33307 , \33306 );
not \U$32965 ( \33308 , \361 );
and \U$32966 ( \33309 , \33307 , \33308 );
and \U$32967 ( \33310 , \33306 , \361 );
nor \U$32968 ( \33311 , \33309 , \33310 );
xor \U$32969 ( \33312 , \33303 , \33311 );
and \U$32970 ( \33313 , \416 , RI986e698_22);
and \U$32971 ( \33314 , RI986f868_60, \414 );
nor \U$32972 ( \33315 , \33313 , \33314 );
and \U$32973 ( \33316 , \33315 , \421 );
not \U$32974 ( \33317 , \33315 );
and \U$32975 ( \33318 , \33317 , \422 );
nor \U$32976 ( \33319 , \33316 , \33318 );
and \U$32977 ( \33320 , \33312 , \33319 );
and \U$32978 ( \33321 , \33303 , \33311 );
nor \U$32979 ( \33322 , \33320 , \33321 );
and \U$32980 ( \33323 , \33295 , \33322 );
and \U$32981 ( \33324 , \33267 , \33294 );
nor \U$32982 ( \33325 , \33323 , \33324 );
xor \U$32983 ( \33326 , \33170 , \33178 );
xor \U$32984 ( \33327 , \33326 , \33187 );
not \U$32985 ( \33328 , \33327 );
nand \U$32986 ( \33329 , RI986e698_22, RI9871fc8_144);
not \U$32987 ( \33330 , \33329 );
and \U$32988 ( \33331 , \33328 , \33330 );
and \U$32989 ( \33332 , \33327 , \33329 );
xor \U$32990 ( \33333 , \33219 , \33226 );
xor \U$32991 ( \33334 , \33333 , \33235 );
nor \U$32992 ( \33335 , \33332 , \33334 );
nor \U$32993 ( \33336 , \33331 , \33335 );
xor \U$32994 ( \33337 , \33325 , \33336 );
not \U$32995 ( \33338 , \33337 );
or \U$32996 ( \33339 , \33243 , \33338 );
or \U$32997 ( \33340 , \33337 , \33242 );
nand \U$32998 ( \33341 , \33339 , \33340 );
nand \U$32999 ( \33342 , \33240 , \33341 );
not \U$33000 ( \33343 , \33342 );
xor \U$33001 ( \33344 , \33275 , \33282 );
xor \U$33002 ( \33345 , \33344 , \33291 );
xor \U$33003 ( \33346 , \33250 , \33255 );
xor \U$33004 ( \33347 , \33346 , \33264 );
and \U$33005 ( \33348 , \33345 , \33347 );
nand \U$33006 ( \33349 , RI986e788_24, RI9871fc8_144);
xor \U$33007 ( \33350 , \33303 , \33311 );
xor \U$33008 ( \33351 , \33350 , \33319 );
nand \U$33009 ( \33352 , \33349 , \33351 );
xor \U$33010 ( \33353 , \33348 , \33352 );
and \U$33011 ( \33354 , \376 , RI986f4a8_52);
and \U$33012 ( \33355 , RI986f3b8_50, \374 );
nor \U$33013 ( \33356 , \33354 , \33355 );
not \U$33014 ( \33357 , \33356 );
not \U$33015 ( \33358 , \367 );
and \U$33016 ( \33359 , \33357 , \33358 );
and \U$33017 ( \33360 , \33356 , \365 );
nor \U$33018 ( \33361 , \33359 , \33360 );
and \U$33019 ( \33362 , \395 , RI986fa48_64);
and \U$33020 ( \33363 , RI986f958_62, \393 );
nor \U$33021 ( \33364 , \33362 , \33363 );
not \U$33022 ( \33365 , \33364 );
not \U$33023 ( \33366 , \487 );
and \U$33024 ( \33367 , \33365 , \33366 );
and \U$33025 ( \33368 , \33364 , \487 );
nor \U$33026 ( \33369 , \33367 , \33368 );
xor \U$33027 ( \33370 , \33361 , \33369 );
and \U$33028 ( \33371 , \354 , RI986f868_60);
and \U$33029 ( \33372 , RI986f778_58, \352 );
nor \U$33030 ( \33373 , \33371 , \33372 );
not \U$33031 ( \33374 , \33373 );
not \U$33032 ( \33375 , \345 );
and \U$33033 ( \33376 , \33374 , \33375 );
and \U$33034 ( \33377 , \33373 , \361 );
nor \U$33035 ( \33378 , \33376 , \33377 );
and \U$33036 ( \33379 , \33370 , \33378 );
and \U$33037 ( \33380 , \33361 , \33369 );
nor \U$33038 ( \33381 , \33379 , \33380 );
and \U$33039 ( \33382 , \1293 , RI986e1e8_12);
and \U$33040 ( \33383 , RI986e0f8_10, \1291 );
nor \U$33041 ( \33384 , \33382 , \33383 );
not \U$33042 ( \33385 , \33384 );
not \U$33043 ( \33386 , \1128 );
and \U$33044 ( \33387 , \33385 , \33386 );
and \U$33045 ( \33388 , \33384 , \1301 );
nor \U$33046 ( \33389 , \33387 , \33388 );
or \U$33047 ( \33390 , \33389 , \1318 );
not \U$33048 ( \33391 , \1318 );
not \U$33049 ( \33392 , \33389 );
or \U$33050 ( \33393 , \33391 , \33392 );
and \U$33051 ( \33394 , \1329 , RI986e2d8_14);
and \U$33052 ( \33395 , RI986e3c8_16, \1327 );
nor \U$33053 ( \33396 , \33394 , \33395 );
and \U$33054 ( \33397 , \33396 , \1336 );
not \U$33055 ( \33398 , \33396 );
and \U$33056 ( \33399 , \33398 , \1337 );
nor \U$33057 ( \33400 , \33397 , \33399 );
nand \U$33058 ( \33401 , \33393 , \33400 );
nand \U$33059 ( \33402 , \33390 , \33401 );
xor \U$33060 ( \33403 , \33381 , \33402 );
not \U$33061 ( \33404 , \454 );
and \U$33062 ( \33405 , \465 , RI986f598_54);
and \U$33063 ( \33406 , RI986f688_56, \463 );
nor \U$33064 ( \33407 , \33405 , \33406 );
not \U$33065 ( \33408 , \33407 );
or \U$33066 ( \33409 , \33404 , \33408 );
or \U$33067 ( \33410 , \33407 , \456 );
nand \U$33068 ( \33411 , \33409 , \33410 );
and \U$33069 ( \33412 , \776 , RI986de28_4);
and \U$33070 ( \33413 , RI986dd38_2, \774 );
nor \U$33071 ( \33414 , \33412 , \33413 );
and \U$33072 ( \33415 , \33414 , \474 );
not \U$33073 ( \33416 , \33414 );
and \U$33074 ( \33417 , \33416 , \451 );
nor \U$33075 ( \33418 , \33415 , \33417 );
xor \U$33076 ( \33419 , \33411 , \33418 );
and \U$33077 ( \33420 , \438 , RI986e008_8);
and \U$33078 ( \33421 , RI986df18_6, \436 );
nor \U$33079 ( \33422 , \33420 , \33421 );
and \U$33080 ( \33423 , \33422 , \444 );
not \U$33081 ( \33424 , \33422 );
and \U$33082 ( \33425 , \33424 , \443 );
nor \U$33083 ( \33426 , \33423 , \33425 );
and \U$33084 ( \33427 , \33419 , \33426 );
and \U$33085 ( \33428 , \33411 , \33418 );
or \U$33086 ( \33429 , \33427 , \33428 );
and \U$33087 ( \33430 , \33403 , \33429 );
and \U$33088 ( \33431 , \33381 , \33402 );
or \U$33089 ( \33432 , \33430 , \33431 );
and \U$33090 ( \33433 , \33353 , \33432 );
and \U$33091 ( \33434 , \33348 , \33352 );
or \U$33092 ( \33435 , \33433 , \33434 );
xor \U$33093 ( \33436 , \33107 , \33108 );
xor \U$33094 ( \33437 , \33436 , \33117 );
xor \U$33095 ( \33438 , \33080 , \33088 );
xor \U$33096 ( \33439 , \33438 , \33097 );
or \U$33097 ( \33440 , \33437 , \33439 );
nand \U$33098 ( \33441 , \33437 , \33439 );
nand \U$33099 ( \33442 , \33440 , \33441 );
xor \U$33100 ( \33443 , \33435 , \33442 );
xor \U$33101 ( \33444 , \33267 , \33294 );
xor \U$33102 ( \33445 , \33444 , \33322 );
not \U$33103 ( \33446 , \33207 );
and \U$33104 ( \33447 , \33198 , \1337 );
not \U$33105 ( \33448 , \33198 );
and \U$33106 ( \33449 , \33448 , \1336 );
nor \U$33107 ( \33450 , \33447 , \33449 );
not \U$33108 ( \33451 , \33450 );
or \U$33109 ( \33452 , \33446 , \33451 );
or \U$33110 ( \33453 , \33450 , \33207 );
nand \U$33111 ( \33454 , \33452 , \33453 );
xor \U$33112 ( \33455 , \33445 , \33454 );
not \U$33113 ( \33456 , \33327 );
xor \U$33114 ( \33457 , \33329 , \33334 );
not \U$33115 ( \33458 , \33457 );
or \U$33116 ( \33459 , \33456 , \33458 );
or \U$33117 ( \33460 , \33457 , \33327 );
nand \U$33118 ( \33461 , \33459 , \33460 );
and \U$33119 ( \33462 , \33455 , \33461 );
and \U$33120 ( \33463 , \33445 , \33454 );
or \U$33121 ( \33464 , \33462 , \33463 );
and \U$33122 ( \33465 , \33443 , \33464 );
and \U$33123 ( \33466 , \33435 , \33442 );
or \U$33124 ( \33467 , \33465 , \33466 );
not \U$33125 ( \33468 , \33467 );
or \U$33126 ( \33469 , \33343 , \33468 );
or \U$33127 ( \33470 , \33467 , \33342 );
nand \U$33128 ( \33471 , \33469 , \33470 );
not \U$33129 ( \33472 , \33471 );
not \U$33130 ( \33473 , \33325 );
not \U$33131 ( \33474 , \33242 );
and \U$33132 ( \33475 , \33473 , \33474 );
and \U$33133 ( \33476 , \33325 , \33242 );
nor \U$33134 ( \33477 , \33476 , \33336 );
nor \U$33135 ( \33478 , \33475 , \33477 );
xor \U$33136 ( \33479 , \33100 , \33120 );
xor \U$33137 ( \33480 , \33479 , \33145 );
xor \U$33138 ( \33481 , \33478 , \33480 );
xor \U$33139 ( \33482 , \33190 , \33210 );
and \U$33140 ( \33483 , \33482 , \33238 );
and \U$33141 ( \33484 , \33190 , \33210 );
or \U$33142 ( \33485 , \33483 , \33484 );
not \U$33143 ( \33486 , \33441 );
xor \U$33144 ( \33487 , \33485 , \33486 );
xor \U$33145 ( \33488 , \32942 , \1301 );
xor \U$33146 ( \33489 , \33488 , \32950 );
xor \U$33147 ( \33490 , \33062 , \33067 );
xor \U$33148 ( \33491 , \33489 , \33490 );
xor \U$33149 ( \33492 , \33487 , \33491 );
xor \U$33150 ( \33493 , \33481 , \33492 );
not \U$33151 ( \33494 , \33493 );
and \U$33152 ( \33495 , \33472 , \33494 );
and \U$33153 ( \33496 , \33471 , \33493 );
nor \U$33154 ( \33497 , \33495 , \33496 );
not \U$33155 ( \33498 , \33497 );
not \U$33156 ( \33499 , \33239 );
not \U$33157 ( \33500 , \33341 );
or \U$33158 ( \33501 , \33499 , \33500 );
or \U$33159 ( \33502 , \33341 , \33239 );
nand \U$33160 ( \33503 , \33501 , \33502 );
not \U$33161 ( \33504 , \33503 );
xor \U$33162 ( \33505 , \33435 , \33442 );
xor \U$33163 ( \33506 , \33505 , \33464 );
not \U$33164 ( \33507 , \33506 );
or \U$33165 ( \33508 , \33504 , \33507 );
or \U$33166 ( \33509 , \33506 , \33503 );
or \U$33167 ( \33510 , \33351 , \33349 );
nand \U$33168 ( \33511 , \33510 , \33352 );
xor \U$33169 ( \33512 , \33345 , \33347 );
xor \U$33170 ( \33513 , \33511 , \33512 );
xor \U$33171 ( \33514 , \33381 , \33402 );
xor \U$33172 ( \33515 , \33514 , \33429 );
and \U$33173 ( \33516 , \33513 , \33515 );
and \U$33174 ( \33517 , \33511 , \33512 );
or \U$33175 ( \33518 , \33516 , \33517 );
and \U$33176 ( \33519 , \1293 , RI986dd38_2);
and \U$33177 ( \33520 , RI986e1e8_12, \1291 );
nor \U$33178 ( \33521 , \33519 , \33520 );
not \U$33179 ( \33522 , \33521 );
not \U$33180 ( \33523 , \1301 );
and \U$33181 ( \33524 , \33522 , \33523 );
and \U$33182 ( \33525 , \33521 , \1128 );
nor \U$33183 ( \33526 , \33524 , \33525 );
nand \U$33184 ( \33527 , RI986e3c8_16, \1311 );
and \U$33185 ( \33528 , \33527 , \1315 );
not \U$33186 ( \33529 , \33527 );
and \U$33187 ( \33530 , \33529 , \1458 );
nor \U$33188 ( \33531 , \33528 , \33530 );
xor \U$33189 ( \33532 , \33526 , \33531 );
and \U$33190 ( \33533 , \1329 , RI986e0f8_10);
and \U$33191 ( \33534 , RI986e2d8_14, \1327 );
nor \U$33192 ( \33535 , \33533 , \33534 );
and \U$33193 ( \33536 , \33535 , \1337 );
not \U$33194 ( \33537 , \33535 );
and \U$33195 ( \33538 , \33537 , \1336 );
nor \U$33196 ( \33539 , \33536 , \33538 );
and \U$33197 ( \33540 , \33532 , \33539 );
and \U$33198 ( \33541 , \33526 , \33531 );
or \U$33199 ( \33542 , \33540 , \33541 );
and \U$33200 ( \33543 , \395 , RI986f778_58);
and \U$33201 ( \33544 , RI986fa48_64, \393 );
nor \U$33202 ( \33545 , \33543 , \33544 );
not \U$33203 ( \33546 , \33545 );
not \U$33204 ( \33547 , \487 );
and \U$33205 ( \33548 , \33546 , \33547 );
and \U$33206 ( \33549 , \33545 , \386 );
nor \U$33207 ( \33550 , \33548 , \33549 );
and \U$33208 ( \33551 , \376 , RI986f958_62);
and \U$33209 ( \33552 , RI986f4a8_52, \374 );
nor \U$33210 ( \33553 , \33551 , \33552 );
not \U$33211 ( \33554 , \33553 );
not \U$33212 ( \33555 , \365 );
and \U$33213 ( \33556 , \33554 , \33555 );
and \U$33214 ( \33557 , \33553 , \367 );
nor \U$33215 ( \33558 , \33556 , \33557 );
xor \U$33216 ( \33559 , \33550 , \33558 );
and \U$33217 ( \33560 , \354 , RI986e698_22);
and \U$33218 ( \33561 , RI986f868_60, \352 );
nor \U$33219 ( \33562 , \33560 , \33561 );
not \U$33220 ( \33563 , \33562 );
not \U$33221 ( \33564 , \345 );
and \U$33222 ( \33565 , \33563 , \33564 );
and \U$33223 ( \33566 , \33562 , \345 );
nor \U$33224 ( \33567 , \33565 , \33566 );
and \U$33225 ( \33568 , \33559 , \33567 );
and \U$33226 ( \33569 , \33550 , \33558 );
or \U$33227 ( \33570 , \33568 , \33569 );
or \U$33228 ( \33571 , \33542 , \33570 );
not \U$33229 ( \33572 , \33542 );
not \U$33230 ( \33573 , \33570 );
or \U$33231 ( \33574 , \33572 , \33573 );
and \U$33232 ( \33575 , \438 , RI986f688_56);
and \U$33233 ( \33576 , RI986e008_8, \436 );
nor \U$33234 ( \33577 , \33575 , \33576 );
and \U$33235 ( \33578 , \33577 , \444 );
not \U$33236 ( \33579 , \33577 );
and \U$33237 ( \33580 , \33579 , \443 );
nor \U$33238 ( \33581 , \33578 , \33580 );
and \U$33239 ( \33582 , \776 , RI986df18_6);
and \U$33240 ( \33583 , RI986de28_4, \774 );
nor \U$33241 ( \33584 , \33582 , \33583 );
and \U$33242 ( \33585 , \33584 , \474 );
not \U$33243 ( \33586 , \33584 );
and \U$33244 ( \33587 , \33586 , \451 );
nor \U$33245 ( \33588 , \33585 , \33587 );
xor \U$33246 ( \33589 , \33581 , \33588 );
not \U$33247 ( \33590 , \456 );
and \U$33248 ( \33591 , \465 , RI986f3b8_50);
and \U$33249 ( \33592 , RI986f598_54, \463 );
nor \U$33250 ( \33593 , \33591 , \33592 );
not \U$33251 ( \33594 , \33593 );
or \U$33252 ( \33595 , \33590 , \33594 );
or \U$33253 ( \33596 , \33593 , \456 );
nand \U$33254 ( \33597 , \33595 , \33596 );
and \U$33255 ( \33598 , \33589 , \33597 );
and \U$33256 ( \33599 , \33581 , \33588 );
or \U$33257 ( \33600 , \33598 , \33599 );
nand \U$33258 ( \33601 , \33574 , \33600 );
nand \U$33259 ( \33602 , \33571 , \33601 );
and \U$33260 ( \33603 , \416 , RI986e788_24);
and \U$33261 ( \33604 , RI986e698_22, \414 );
nor \U$33262 ( \33605 , \33603 , \33604 );
and \U$33263 ( \33606 , \33605 , \421 );
not \U$33264 ( \33607 , \33605 );
and \U$33265 ( \33608 , \33607 , \422 );
nor \U$33266 ( \33609 , \33606 , \33608 );
nand \U$33267 ( \33610 , RI986e4b8_18, RI9871fc8_144);
or \U$33268 ( \33611 , \33609 , \33610 );
not \U$33269 ( \33612 , \33610 );
not \U$33270 ( \33613 , \33609 );
or \U$33271 ( \33614 , \33612 , \33613 );
nand \U$33272 ( \33615 , RI986e5a8_20, RI9871fc8_144);
and \U$33273 ( \33616 , \416 , RI986e4b8_18);
and \U$33274 ( \33617 , RI986e788_24, \414 );
nor \U$33275 ( \33618 , \33616 , \33617 );
and \U$33276 ( \33619 , \33618 , \421 );
not \U$33277 ( \33620 , \33618 );
and \U$33278 ( \33621 , \33620 , \422 );
nor \U$33279 ( \33622 , \33619 , \33621 );
nand \U$33280 ( \33623 , \33615 , \33622 );
nand \U$33281 ( \33624 , \33614 , \33623 );
nand \U$33282 ( \33625 , \33611 , \33624 );
xor \U$33283 ( \33626 , \33602 , \33625 );
not \U$33284 ( \33627 , \1315 );
not \U$33285 ( \33628 , \33400 );
or \U$33286 ( \33629 , \33627 , \33628 );
or \U$33287 ( \33630 , \33400 , \1318 );
nand \U$33288 ( \33631 , \33629 , \33630 );
not \U$33289 ( \33632 , \33631 );
not \U$33290 ( \33633 , \33389 );
and \U$33291 ( \33634 , \33632 , \33633 );
and \U$33292 ( \33635 , \33631 , \33389 );
nor \U$33293 ( \33636 , \33634 , \33635 );
xor \U$33294 ( \33637 , \33361 , \33369 );
xor \U$33295 ( \33638 , \33637 , \33378 );
or \U$33296 ( \33639 , \33636 , \33638 );
not \U$33297 ( \33640 , \33638 );
not \U$33298 ( \33641 , \33636 );
or \U$33299 ( \33642 , \33640 , \33641 );
xor \U$33300 ( \33643 , \33411 , \33418 );
xor \U$33301 ( \33644 , \33643 , \33426 );
nand \U$33302 ( \33645 , \33642 , \33644 );
nand \U$33303 ( \33646 , \33639 , \33645 );
and \U$33304 ( \33647 , \33626 , \33646 );
and \U$33305 ( \33648 , \33602 , \33625 );
or \U$33306 ( \33649 , \33647 , \33648 );
xor \U$33307 ( \33650 , \33518 , \33649 );
xor \U$33308 ( \33651 , \33445 , \33454 );
xor \U$33309 ( \33652 , \33651 , \33461 );
and \U$33310 ( \33653 , \33650 , \33652 );
and \U$33311 ( \33654 , \33518 , \33649 );
or \U$33312 ( \33655 , \33653 , \33654 );
nand \U$33313 ( \33656 , \33509 , \33655 );
nand \U$33314 ( \33657 , \33508 , \33656 );
nand \U$33315 ( \33658 , \33498 , \33657 );
xor \U$33316 ( \33659 , \33478 , \33480 );
and \U$33317 ( \33660 , \33659 , \33492 );
and \U$33318 ( \33661 , \33478 , \33480 );
or \U$33319 ( \33662 , \33660 , \33661 );
not \U$33320 ( \33663 , \33662 );
or \U$33321 ( \33664 , \33493 , \33342 );
not \U$33322 ( \33665 , \33342 );
not \U$33323 ( \33666 , \33493 );
or \U$33324 ( \33667 , \33665 , \33666 );
nand \U$33325 ( \33668 , \33667 , \33467 );
nand \U$33326 ( \33669 , \33664 , \33668 );
not \U$33327 ( \33670 , \33669 );
or \U$33328 ( \33671 , \33663 , \33670 );
or \U$33329 ( \33672 , \33669 , \33662 );
nand \U$33330 ( \33673 , \33671 , \33672 );
not \U$33331 ( \33674 , \33673 );
xor \U$33332 ( \33675 , \33485 , \33486 );
and \U$33333 ( \33676 , \33675 , \33491 );
and \U$33334 ( \33677 , \33485 , \33486 );
or \U$33335 ( \33678 , \33676 , \33677 );
xor \U$33336 ( \33679 , \32935 , \32953 );
xor \U$33337 ( \33680 , \33679 , \32982 );
xor \U$33338 ( \33681 , \33678 , \33680 );
xor \U$33339 ( \33682 , \33072 , \33148 );
xor \U$33340 ( \33683 , \33682 , \33155 );
xor \U$33341 ( \33684 , \33681 , \33683 );
not \U$33342 ( \33685 , \33684 );
and \U$33343 ( \33686 , \33674 , \33685 );
and \U$33344 ( \33687 , \33673 , \33684 );
nor \U$33345 ( \33688 , \33686 , \33687 );
xor \U$33346 ( \33689 , \33658 , \33688 );
not \U$33347 ( \33690 , \33609 );
not \U$33348 ( \33691 , \33623 );
or \U$33349 ( \33692 , \33690 , \33691 );
or \U$33350 ( \33693 , \33623 , \33609 );
nand \U$33351 ( \33694 , \33692 , \33693 );
not \U$33352 ( \33695 , \33694 );
not \U$33353 ( \33696 , \33610 );
and \U$33354 ( \33697 , \33695 , \33696 );
and \U$33355 ( \33698 , \33694 , \33610 );
nor \U$33356 ( \33699 , \33697 , \33698 );
not \U$33357 ( \33700 , \33600 );
not \U$33358 ( \33701 , \33570 );
or \U$33359 ( \33702 , \33700 , \33701 );
or \U$33360 ( \33703 , \33570 , \33600 );
nand \U$33361 ( \33704 , \33702 , \33703 );
not \U$33362 ( \33705 , \33704 );
not \U$33363 ( \33706 , \33542 );
and \U$33364 ( \33707 , \33705 , \33706 );
and \U$33365 ( \33708 , \33704 , \33542 );
nor \U$33366 ( \33709 , \33707 , \33708 );
xor \U$33367 ( \33710 , \33699 , \33709 );
not \U$33368 ( \33711 , \33644 );
not \U$33369 ( \33712 , \33636 );
or \U$33370 ( \33713 , \33711 , \33712 );
or \U$33371 ( \33714 , \33636 , \33644 );
nand \U$33372 ( \33715 , \33713 , \33714 );
not \U$33373 ( \33716 , \33715 );
not \U$33374 ( \33717 , \33638 );
and \U$33375 ( \33718 , \33716 , \33717 );
and \U$33376 ( \33719 , \33715 , \33638 );
nor \U$33377 ( \33720 , \33718 , \33719 );
and \U$33378 ( \33721 , \33710 , \33720 );
and \U$33379 ( \33722 , \33699 , \33709 );
nor \U$33380 ( \33723 , \33721 , \33722 );
and \U$33381 ( \33724 , \465 , RI986f4a8_52);
and \U$33382 ( \33725 , RI986f3b8_50, \463 );
nor \U$33383 ( \33726 , \33724 , \33725 );
not \U$33384 ( \33727 , \33726 );
not \U$33385 ( \33728 , \456 );
and \U$33386 ( \33729 , \33727 , \33728 );
and \U$33387 ( \33730 , \33726 , \454 );
nor \U$33388 ( \33731 , \33729 , \33730 );
and \U$33389 ( \33732 , \376 , RI986fa48_64);
and \U$33390 ( \33733 , RI986f958_62, \374 );
nor \U$33391 ( \33734 , \33732 , \33733 );
not \U$33392 ( \33735 , \33734 );
not \U$33393 ( \33736 , \367 );
and \U$33394 ( \33737 , \33735 , \33736 );
and \U$33395 ( \33738 , \33734 , \367 );
nor \U$33396 ( \33739 , \33737 , \33738 );
xor \U$33397 ( \33740 , \33731 , \33739 );
and \U$33398 ( \33741 , \395 , RI986f868_60);
and \U$33399 ( \33742 , RI986f778_58, \393 );
nor \U$33400 ( \33743 , \33741 , \33742 );
not \U$33401 ( \33744 , \33743 );
not \U$33402 ( \33745 , \386 );
and \U$33403 ( \33746 , \33744 , \33745 );
and \U$33404 ( \33747 , \33743 , \487 );
nor \U$33405 ( \33748 , \33746 , \33747 );
and \U$33406 ( \33749 , \33740 , \33748 );
and \U$33407 ( \33750 , \33731 , \33739 );
or \U$33408 ( \33751 , \33749 , \33750 );
and \U$33409 ( \33752 , \1311 , RI986e2d8_14);
and \U$33410 ( \33753 , RI986e3c8_16, \1309 );
nor \U$33411 ( \33754 , \33752 , \33753 );
and \U$33412 ( \33755 , \33754 , \1315 );
not \U$33413 ( \33756 , \33754 );
and \U$33414 ( \33757 , \33756 , \1319 );
nor \U$33415 ( \33758 , \33755 , \33757 );
xor \U$33416 ( \33759 , \33758 , \2034 );
and \U$33417 ( \33760 , \1329 , RI986e1e8_12);
and \U$33418 ( \33761 , RI986e0f8_10, \1327 );
nor \U$33419 ( \33762 , \33760 , \33761 );
and \U$33420 ( \33763 , \33762 , \1337 );
not \U$33421 ( \33764 , \33762 );
and \U$33422 ( \33765 , \33764 , \1336 );
nor \U$33423 ( \33766 , \33763 , \33765 );
and \U$33424 ( \33767 , \33759 , \33766 );
and \U$33425 ( \33768 , \33758 , \2034 );
or \U$33426 ( \33769 , \33767 , \33768 );
xor \U$33427 ( \33770 , \33751 , \33769 );
and \U$33428 ( \33771 , \438 , RI986f598_54);
and \U$33429 ( \33772 , RI986f688_56, \436 );
nor \U$33430 ( \33773 , \33771 , \33772 );
and \U$33431 ( \33774 , \33773 , \443 );
not \U$33432 ( \33775 , \33773 );
and \U$33433 ( \33776 , \33775 , \444 );
nor \U$33434 ( \33777 , \33774 , \33776 );
not \U$33435 ( \33778 , \33777 );
and \U$33436 ( \33779 , \1293 , RI986de28_4);
and \U$33437 ( \33780 , RI986dd38_2, \1291 );
nor \U$33438 ( \33781 , \33779 , \33780 );
not \U$33439 ( \33782 , \33781 );
not \U$33440 ( \33783 , \1128 );
and \U$33441 ( \33784 , \33782 , \33783 );
and \U$33442 ( \33785 , \33781 , \1128 );
nor \U$33443 ( \33786 , \33784 , \33785 );
not \U$33444 ( \33787 , \33786 );
and \U$33445 ( \33788 , \33778 , \33787 );
and \U$33446 ( \33789 , \33786 , \33777 );
and \U$33447 ( \33790 , \776 , RI986e008_8);
and \U$33448 ( \33791 , RI986df18_6, \774 );
nor \U$33449 ( \33792 , \33790 , \33791 );
and \U$33450 ( \33793 , \33792 , \451 );
not \U$33451 ( \33794 , \33792 );
and \U$33452 ( \33795 , \33794 , \474 );
nor \U$33453 ( \33796 , \33793 , \33795 );
nor \U$33454 ( \33797 , \33789 , \33796 );
nor \U$33455 ( \33798 , \33788 , \33797 );
and \U$33456 ( \33799 , \33770 , \33798 );
and \U$33457 ( \33800 , \33751 , \33769 );
or \U$33458 ( \33801 , \33799 , \33800 );
xor \U$33459 ( \33802 , \33526 , \33531 );
xor \U$33460 ( \33803 , \33802 , \33539 );
not \U$33461 ( \33804 , \33803 );
xor \U$33462 ( \33805 , \33581 , \33588 );
xor \U$33463 ( \33806 , \33805 , \33597 );
nand \U$33464 ( \33807 , \33804 , \33806 );
or \U$33465 ( \33808 , \33801 , \33807 );
not \U$33466 ( \33809 , \33807 );
not \U$33467 ( \33810 , \33801 );
or \U$33468 ( \33811 , \33809 , \33810 );
xor \U$33469 ( \33812 , \33550 , \33558 );
xor \U$33470 ( \33813 , \33812 , \33567 );
and \U$33471 ( \33814 , \354 , RI986e788_24);
and \U$33472 ( \33815 , RI986e698_22, \352 );
nor \U$33473 ( \33816 , \33814 , \33815 );
not \U$33474 ( \33817 , \33816 );
not \U$33475 ( \33818 , \361 );
and \U$33476 ( \33819 , \33817 , \33818 );
and \U$33477 ( \33820 , \33816 , \361 );
nor \U$33478 ( \33821 , \33819 , \33820 );
nand \U$33479 ( \33822 , RI986f1d8_46, RI9871fc8_144);
xor \U$33480 ( \33823 , \33821 , \33822 );
and \U$33481 ( \33824 , \416 , RI986e5a8_20);
and \U$33482 ( \33825 , RI986e4b8_18, \414 );
nor \U$33483 ( \33826 , \33824 , \33825 );
and \U$33484 ( \33827 , \33826 , \421 );
not \U$33485 ( \33828 , \33826 );
and \U$33486 ( \33829 , \33828 , \422 );
nor \U$33487 ( \33830 , \33827 , \33829 );
and \U$33488 ( \33831 , \33823 , \33830 );
and \U$33489 ( \33832 , \33821 , \33822 );
or \U$33490 ( \33833 , \33831 , \33832 );
or \U$33491 ( \33834 , \33813 , \33833 );
not \U$33492 ( \33835 , \33833 );
not \U$33493 ( \33836 , \33813 );
or \U$33494 ( \33837 , \33835 , \33836 );
or \U$33495 ( \33838 , \33622 , \33615 );
nand \U$33496 ( \33839 , \33838 , \33623 );
nand \U$33497 ( \33840 , \33837 , \33839 );
nand \U$33498 ( \33841 , \33834 , \33840 );
nand \U$33499 ( \33842 , \33811 , \33841 );
nand \U$33500 ( \33843 , \33808 , \33842 );
xor \U$33501 ( \33844 , \33723 , \33843 );
xor \U$33502 ( \33845 , \33511 , \33512 );
xor \U$33503 ( \33846 , \33845 , \33515 );
xor \U$33504 ( \33847 , \33844 , \33846 );
xor \U$33505 ( \33848 , \33602 , \33625 );
xor \U$33506 ( \33849 , \33848 , \33646 );
and \U$33507 ( \33850 , \33847 , \33849 );
not \U$33508 ( \33851 , \33847 );
not \U$33509 ( \33852 , \33849 );
and \U$33510 ( \33853 , \33851 , \33852 );
not \U$33511 ( \33854 , \33803 );
not \U$33512 ( \33855 , \33806 );
and \U$33513 ( \33856 , \33854 , \33855 );
and \U$33514 ( \33857 , \33803 , \33806 );
nor \U$33515 ( \33858 , \33856 , \33857 );
xor \U$33516 ( \33859 , \33751 , \33769 );
xor \U$33517 ( \33860 , \33859 , \33798 );
and \U$33518 ( \33861 , \33858 , \33860 );
xnor \U$33519 ( \33862 , \33833 , \33813 );
not \U$33520 ( \33863 , \33862 );
not \U$33521 ( \33864 , \33839 );
and \U$33522 ( \33865 , \33863 , \33864 );
and \U$33523 ( \33866 , \33862 , \33839 );
nor \U$33524 ( \33867 , \33865 , \33866 );
xor \U$33525 ( \33868 , \33751 , \33769 );
xor \U$33526 ( \33869 , \33868 , \33798 );
and \U$33527 ( \33870 , \33867 , \33869 );
and \U$33528 ( \33871 , \33858 , \33867 );
or \U$33529 ( \33872 , \33861 , \33870 , \33871 );
not \U$33530 ( \33873 , \454 );
and \U$33531 ( \33874 , \465 , RI986f958_62);
and \U$33532 ( \33875 , RI986f4a8_52, \463 );
nor \U$33533 ( \33876 , \33874 , \33875 );
not \U$33534 ( \33877 , \33876 );
or \U$33535 ( \33878 , \33873 , \33877 );
or \U$33536 ( \33879 , \33876 , \454 );
nand \U$33537 ( \33880 , \33878 , \33879 );
not \U$33538 ( \33881 , \365 );
and \U$33539 ( \33882 , \376 , RI986f778_58);
and \U$33540 ( \33883 , RI986fa48_64, \374 );
nor \U$33541 ( \33884 , \33882 , \33883 );
not \U$33542 ( \33885 , \33884 );
or \U$33543 ( \33886 , \33881 , \33885 );
or \U$33544 ( \33887 , \33884 , \367 );
nand \U$33545 ( \33888 , \33886 , \33887 );
xor \U$33546 ( \33889 , \33880 , \33888 );
not \U$33547 ( \33890 , \386 );
and \U$33548 ( \33891 , \395 , RI986e698_22);
and \U$33549 ( \33892 , RI986f868_60, \393 );
nor \U$33550 ( \33893 , \33891 , \33892 );
not \U$33551 ( \33894 , \33893 );
or \U$33552 ( \33895 , \33890 , \33894 );
or \U$33553 ( \33896 , \33893 , \487 );
nand \U$33554 ( \33897 , \33895 , \33896 );
and \U$33555 ( \33898 , \33889 , \33897 );
and \U$33556 ( \33899 , \33880 , \33888 );
nor \U$33557 ( \33900 , \33898 , \33899 );
and \U$33558 ( \33901 , \1329 , RI986dd38_2);
and \U$33559 ( \33902 , RI986e1e8_12, \1327 );
nor \U$33560 ( \33903 , \33901 , \33902 );
and \U$33561 ( \33904 , \33903 , \1337 );
not \U$33562 ( \33905 , \33903 );
and \U$33563 ( \33906 , \33905 , \1336 );
nor \U$33564 ( \33907 , \33904 , \33906 );
not \U$33565 ( \33908 , \33907 );
and \U$33566 ( \33909 , \1311 , RI986e0f8_10);
and \U$33567 ( \33910 , RI986e2d8_14, \1309 );
nor \U$33568 ( \33911 , \33909 , \33910 );
and \U$33569 ( \33912 , \33911 , \1315 );
not \U$33570 ( \33913 , \33911 );
and \U$33571 ( \33914 , \33913 , \1458 );
nor \U$33572 ( \33915 , \33912 , \33914 );
not \U$33573 ( \33916 , \33915 );
and \U$33574 ( \33917 , \33908 , \33916 );
and \U$33575 ( \33918 , \33915 , \33907 );
nand \U$33576 ( \33919 , RI986e3c8_16, \2042 );
not \U$33577 ( \33920 , \33919 );
not \U$33578 ( \33921 , \2034 );
and \U$33579 ( \33922 , \33920 , \33921 );
and \U$33580 ( \33923 , \33919 , \1462 );
nor \U$33581 ( \33924 , \33922 , \33923 );
nor \U$33582 ( \33925 , \33918 , \33924 );
nor \U$33583 ( \33926 , \33917 , \33925 );
xor \U$33584 ( \33927 , \33900 , \33926 );
and \U$33585 ( \33928 , \776 , RI986f688_56);
and \U$33586 ( \33929 , RI986e008_8, \774 );
nor \U$33587 ( \33930 , \33928 , \33929 );
and \U$33588 ( \33931 , \33930 , \474 );
not \U$33589 ( \33932 , \33930 );
and \U$33590 ( \33933 , \33932 , \451 );
nor \U$33591 ( \33934 , \33931 , \33933 );
not \U$33592 ( \33935 , \1128 );
and \U$33593 ( \33936 , \1293 , RI986df18_6);
and \U$33594 ( \33937 , RI986de28_4, \1291 );
nor \U$33595 ( \33938 , \33936 , \33937 );
not \U$33596 ( \33939 , \33938 );
or \U$33597 ( \33940 , \33935 , \33939 );
or \U$33598 ( \33941 , \33938 , \1128 );
nand \U$33599 ( \33942 , \33940 , \33941 );
xor \U$33600 ( \33943 , \33934 , \33942 );
and \U$33601 ( \33944 , \438 , RI986f3b8_50);
and \U$33602 ( \33945 , RI986f598_54, \436 );
nor \U$33603 ( \33946 , \33944 , \33945 );
and \U$33604 ( \33947 , \33946 , \444 );
not \U$33605 ( \33948 , \33946 );
and \U$33606 ( \33949 , \33948 , \443 );
nor \U$33607 ( \33950 , \33947 , \33949 );
and \U$33608 ( \33951 , \33943 , \33950 );
and \U$33609 ( \33952 , \33934 , \33942 );
nor \U$33610 ( \33953 , \33951 , \33952 );
and \U$33611 ( \33954 , \33927 , \33953 );
and \U$33612 ( \33955 , \33900 , \33926 );
or \U$33613 ( \33956 , \33954 , \33955 );
xor \U$33614 ( \33957 , \33758 , \2034 );
xor \U$33615 ( \33958 , \33957 , \33766 );
not \U$33616 ( \33959 , \33958 );
not \U$33617 ( \33960 , \33777 );
xor \U$33618 ( \33961 , \33796 , \33786 );
not \U$33619 ( \33962 , \33961 );
or \U$33620 ( \33963 , \33960 , \33962 );
or \U$33621 ( \33964 , \33961 , \33777 );
nand \U$33622 ( \33965 , \33963 , \33964 );
nand \U$33623 ( \33966 , \33959 , \33965 );
xor \U$33624 ( \33967 , \33956 , \33966 );
and \U$33625 ( \33968 , \416 , RI986f1d8_46);
and \U$33626 ( \33969 , RI986e5a8_20, \414 );
nor \U$33627 ( \33970 , \33968 , \33969 );
and \U$33628 ( \33971 , \33970 , \421 );
not \U$33629 ( \33972 , \33970 );
and \U$33630 ( \33973 , \33972 , \422 );
nor \U$33631 ( \33974 , \33971 , \33973 );
nand \U$33632 ( \33975 , RI986f2c8_48, RI9871fc8_144);
xor \U$33633 ( \33976 , \33974 , \33975 );
and \U$33634 ( \33977 , \354 , RI986e4b8_18);
and \U$33635 ( \33978 , RI986e788_24, \352 );
nor \U$33636 ( \33979 , \33977 , \33978 );
not \U$33637 ( \33980 , \33979 );
not \U$33638 ( \33981 , \345 );
and \U$33639 ( \33982 , \33980 , \33981 );
and \U$33640 ( \33983 , \33979 , \345 );
nor \U$33641 ( \33984 , \33982 , \33983 );
and \U$33642 ( \33985 , \33976 , \33984 );
and \U$33643 ( \33986 , \33974 , \33975 );
or \U$33644 ( \33987 , \33985 , \33986 );
xor \U$33645 ( \33988 , \33821 , \33822 );
xor \U$33646 ( \33989 , \33988 , \33830 );
and \U$33647 ( \33990 , \33987 , \33989 );
xor \U$33648 ( \33991 , \33731 , \33739 );
xor \U$33649 ( \33992 , \33991 , \33748 );
xor \U$33650 ( \33993 , \33821 , \33822 );
xor \U$33651 ( \33994 , \33993 , \33830 );
and \U$33652 ( \33995 , \33992 , \33994 );
and \U$33653 ( \33996 , \33987 , \33992 );
or \U$33654 ( \33997 , \33990 , \33995 , \33996 );
and \U$33655 ( \33998 , \33967 , \33997 );
and \U$33656 ( \33999 , \33956 , \33966 );
or \U$33657 ( \34000 , \33998 , \33999 );
xor \U$33658 ( \34001 , \33872 , \34000 );
xor \U$33659 ( \34002 , \33699 , \33709 );
xor \U$33660 ( \34003 , \34002 , \33720 );
and \U$33661 ( \34004 , \34001 , \34003 );
and \U$33662 ( \34005 , \33872 , \34000 );
or \U$33663 ( \34006 , \34004 , \34005 );
nor \U$33664 ( \34007 , \33853 , \34006 );
nor \U$33665 ( \34008 , \33850 , \34007 );
not \U$33666 ( \34009 , \34008 );
xor \U$33667 ( \34010 , \33723 , \33843 );
and \U$33668 ( \34011 , \34010 , \33846 );
and \U$33669 ( \34012 , \33723 , \33843 );
or \U$33670 ( \34013 , \34011 , \34012 );
xor \U$33671 ( \34014 , \33348 , \33352 );
xor \U$33672 ( \34015 , \34014 , \33432 );
xor \U$33673 ( \34016 , \34013 , \34015 );
xor \U$33674 ( \34017 , \33518 , \33649 );
xor \U$33675 ( \34018 , \34017 , \33652 );
xor \U$33676 ( \34019 , \34016 , \34018 );
nand \U$33677 ( \34020 , \34009 , \34019 );
xnor \U$33678 ( \34021 , \33655 , \33506 );
not \U$33679 ( \34022 , \34021 );
not \U$33680 ( \34023 , \33503 );
and \U$33681 ( \34024 , \34022 , \34023 );
and \U$33682 ( \34025 , \34021 , \33503 );
nor \U$33683 ( \34026 , \34024 , \34025 );
not \U$33684 ( \34027 , \34026 );
xor \U$33685 ( \34028 , \34013 , \34015 );
and \U$33686 ( \34029 , \34028 , \34018 );
and \U$33687 ( \34030 , \34013 , \34015 );
or \U$33688 ( \34031 , \34029 , \34030 );
not \U$33689 ( \34032 , \34031 );
and \U$33690 ( \34033 , \34027 , \34032 );
and \U$33691 ( \34034 , \34026 , \34031 );
nor \U$33692 ( \34035 , \34033 , \34034 );
xor \U$33693 ( \34036 , \34020 , \34035 );
not \U$33694 ( \34037 , \33847 );
not \U$33695 ( \34038 , \34006 );
not \U$33696 ( \34039 , \33849 );
and \U$33697 ( \34040 , \34038 , \34039 );
and \U$33698 ( \34041 , \34006 , \33849 );
nor \U$33699 ( \34042 , \34040 , \34041 );
not \U$33700 ( \34043 , \34042 );
or \U$33701 ( \34044 , \34037 , \34043 );
or \U$33702 ( \34045 , \34042 , \33847 );
nand \U$33703 ( \34046 , \34044 , \34045 );
not \U$33704 ( \34047 , \34046 );
xor \U$33705 ( \34048 , \33872 , \34000 );
xor \U$33706 ( \34049 , \34048 , \34003 );
not \U$33707 ( \34050 , \34049 );
not \U$33708 ( \34051 , \33841 );
not \U$33709 ( \34052 , \33801 );
and \U$33710 ( \34053 , \34051 , \34052 );
and \U$33711 ( \34054 , \33841 , \33801 );
nor \U$33712 ( \34055 , \34053 , \34054 );
xnor \U$33713 ( \34056 , \34055 , \33807 );
not \U$33714 ( \34057 , \34056 );
and \U$33715 ( \34058 , \34050 , \34057 );
and \U$33716 ( \34059 , \34049 , \34056 );
xor \U$33717 ( \34060 , \33900 , \33926 );
xor \U$33718 ( \34061 , \34060 , \33953 );
not \U$33719 ( \34062 , \34061 );
not \U$33720 ( \34063 , \33958 );
not \U$33721 ( \34064 , \33965 );
and \U$33722 ( \34065 , \34063 , \34064 );
and \U$33723 ( \34066 , \33958 , \33965 );
nor \U$33724 ( \34067 , \34065 , \34066 );
not \U$33725 ( \34068 , \34067 );
and \U$33726 ( \34069 , \34062 , \34068 );
and \U$33727 ( \34070 , \34061 , \34067 );
xor \U$33728 ( \34071 , \33821 , \33822 );
xor \U$33729 ( \34072 , \34071 , \33830 );
xor \U$33730 ( \34073 , \33987 , \33992 );
xor \U$33731 ( \34074 , \34072 , \34073 );
nor \U$33732 ( \34075 , \34070 , \34074 );
nor \U$33733 ( \34076 , \34069 , \34075 );
and \U$33734 ( \34077 , \354 , RI986e5a8_20);
and \U$33735 ( \34078 , RI986e4b8_18, \352 );
nor \U$33736 ( \34079 , \34077 , \34078 );
not \U$33737 ( \34080 , \34079 );
not \U$33738 ( \34081 , \345 );
and \U$33739 ( \34082 , \34080 , \34081 );
and \U$33740 ( \34083 , \34079 , \361 );
nor \U$33741 ( \34084 , \34082 , \34083 );
and \U$33742 ( \34085 , \395 , RI986e788_24);
and \U$33743 ( \34086 , RI986e698_22, \393 );
nor \U$33744 ( \34087 , \34085 , \34086 );
not \U$33745 ( \34088 , \34087 );
not \U$33746 ( \34089 , \386 );
and \U$33747 ( \34090 , \34088 , \34089 );
and \U$33748 ( \34091 , \34087 , \386 );
nor \U$33749 ( \34092 , \34090 , \34091 );
xor \U$33750 ( \34093 , \34084 , \34092 );
and \U$33751 ( \34094 , \416 , RI986f2c8_48);
and \U$33752 ( \34095 , RI986f1d8_46, \414 );
nor \U$33753 ( \34096 , \34094 , \34095 );
and \U$33754 ( \34097 , \34096 , \421 );
not \U$33755 ( \34098 , \34096 );
and \U$33756 ( \34099 , \34098 , \422 );
nor \U$33757 ( \34100 , \34097 , \34099 );
and \U$33758 ( \34101 , \34093 , \34100 );
and \U$33759 ( \34102 , \34084 , \34092 );
or \U$33760 ( \34103 , \34101 , \34102 );
xor \U$33761 ( \34104 , \33974 , \33975 );
xor \U$33762 ( \34105 , \34104 , \33984 );
nand \U$33763 ( \34106 , \34103 , \34105 );
and \U$33764 ( \34107 , \465 , RI986fa48_64);
and \U$33765 ( \34108 , RI986f958_62, \463 );
nor \U$33766 ( \34109 , \34107 , \34108 );
not \U$33767 ( \34110 , \34109 );
not \U$33768 ( \34111 , \456 );
and \U$33769 ( \34112 , \34110 , \34111 );
and \U$33770 ( \34113 , \34109 , \454 );
nor \U$33771 ( \34114 , \34112 , \34113 );
and \U$33772 ( \34115 , \376 , RI986f868_60);
and \U$33773 ( \34116 , RI986f778_58, \374 );
nor \U$33774 ( \34117 , \34115 , \34116 );
not \U$33775 ( \34118 , \34117 );
not \U$33776 ( \34119 , \367 );
and \U$33777 ( \34120 , \34118 , \34119 );
and \U$33778 ( \34121 , \34117 , \365 );
nor \U$33779 ( \34122 , \34120 , \34121 );
or \U$33780 ( \34123 , \34114 , \34122 );
not \U$33781 ( \34124 , \34122 );
not \U$33782 ( \34125 , \34114 );
or \U$33783 ( \34126 , \34124 , \34125 );
and \U$33784 ( \34127 , \438 , RI986f4a8_52);
and \U$33785 ( \34128 , RI986f3b8_50, \436 );
nor \U$33786 ( \34129 , \34127 , \34128 );
and \U$33787 ( \34130 , \34129 , \444 );
not \U$33788 ( \34131 , \34129 );
and \U$33789 ( \34132 , \34131 , \443 );
nor \U$33790 ( \34133 , \34130 , \34132 );
nand \U$33791 ( \34134 , \34126 , \34133 );
nand \U$33792 ( \34135 , \34123 , \34134 );
and \U$33793 ( \34136 , \2042 , RI986e2d8_14);
and \U$33794 ( \34137 , RI986e3c8_16, \2040 );
nor \U$33795 ( \34138 , \34136 , \34137 );
not \U$33796 ( \34139 , \34138 );
not \U$33797 ( \34140 , \2034 );
and \U$33798 ( \34141 , \34139 , \34140 );
and \U$33799 ( \34142 , \34138 , \2034 );
nor \U$33800 ( \34143 , \34141 , \34142 );
or \U$33801 ( \34144 , \34143 , \2031 );
and \U$33802 ( \34145 , \34143 , \2031 );
and \U$33803 ( \34146 , \1311 , RI986e1e8_12);
and \U$33804 ( \34147 , RI986e0f8_10, \1309 );
nor \U$33805 ( \34148 , \34146 , \34147 );
and \U$33806 ( \34149 , \34148 , \1315 );
not \U$33807 ( \34150 , \34148 );
and \U$33808 ( \34151 , \34150 , \1458 );
nor \U$33809 ( \34152 , \34149 , \34151 );
nor \U$33810 ( \34153 , \34145 , \34152 );
not \U$33811 ( \34154 , \34153 );
nand \U$33812 ( \34155 , \34144 , \34154 );
xor \U$33813 ( \34156 , \34135 , \34155 );
and \U$33814 ( \34157 , \776 , RI986f598_54);
and \U$33815 ( \34158 , RI986f688_56, \774 );
nor \U$33816 ( \34159 , \34157 , \34158 );
and \U$33817 ( \34160 , \34159 , \451 );
not \U$33818 ( \34161 , \34159 );
and \U$33819 ( \34162 , \34161 , \474 );
nor \U$33820 ( \34163 , \34160 , \34162 );
and \U$33821 ( \34164 , \1293 , RI986e008_8);
and \U$33822 ( \34165 , RI986df18_6, \1291 );
nor \U$33823 ( \34166 , \34164 , \34165 );
not \U$33824 ( \34167 , \34166 );
not \U$33825 ( \34168 , \1128 );
and \U$33826 ( \34169 , \34167 , \34168 );
and \U$33827 ( \34170 , \34166 , \1301 );
nor \U$33828 ( \34171 , \34169 , \34170 );
or \U$33829 ( \34172 , \34163 , \34171 );
not \U$33830 ( \34173 , \34171 );
not \U$33831 ( \34174 , \34163 );
or \U$33832 ( \34175 , \34173 , \34174 );
and \U$33833 ( \34176 , \1329 , RI986de28_4);
and \U$33834 ( \34177 , RI986dd38_2, \1327 );
nor \U$33835 ( \34178 , \34176 , \34177 );
and \U$33836 ( \34179 , \34178 , \1336 );
not \U$33837 ( \34180 , \34178 );
and \U$33838 ( \34181 , \34180 , \1337 );
nor \U$33839 ( \34182 , \34179 , \34181 );
nand \U$33840 ( \34183 , \34175 , \34182 );
nand \U$33841 ( \34184 , \34172 , \34183 );
and \U$33842 ( \34185 , \34156 , \34184 );
and \U$33843 ( \34186 , \34135 , \34155 );
or \U$33844 ( \34187 , \34185 , \34186 );
xor \U$33845 ( \34188 , \34106 , \34187 );
not \U$33846 ( \34189 , \33907 );
xor \U$33847 ( \34190 , \33924 , \33915 );
not \U$33848 ( \34191 , \34190 );
or \U$33849 ( \34192 , \34189 , \34191 );
or \U$33850 ( \34193 , \34190 , \33907 );
nand \U$33851 ( \34194 , \34192 , \34193 );
xor \U$33852 ( \34195 , \33880 , \33888 );
xor \U$33853 ( \34196 , \34195 , \33897 );
xor \U$33854 ( \34197 , \34194 , \34196 );
xor \U$33855 ( \34198 , \33934 , \33942 );
xor \U$33856 ( \34199 , \34198 , \33950 );
and \U$33857 ( \34200 , \34197 , \34199 );
and \U$33858 ( \34201 , \34194 , \34196 );
or \U$33859 ( \34202 , \34200 , \34201 );
and \U$33860 ( \34203 , \34188 , \34202 );
and \U$33861 ( \34204 , \34106 , \34187 );
nor \U$33862 ( \34205 , \34203 , \34204 );
xor \U$33863 ( \34206 , \34076 , \34205 );
xor \U$33864 ( \34207 , \33751 , \33769 );
xor \U$33865 ( \34208 , \34207 , \33798 );
xor \U$33866 ( \34209 , \33858 , \33867 );
xor \U$33867 ( \34210 , \34208 , \34209 );
and \U$33868 ( \34211 , \34206 , \34210 );
and \U$33869 ( \34212 , \34076 , \34205 );
or \U$33870 ( \34213 , \34211 , \34212 );
nor \U$33871 ( \34214 , \34059 , \34213 );
nor \U$33872 ( \34215 , \34058 , \34214 );
not \U$33873 ( \34216 , \34215 );
and \U$33874 ( \34217 , \34047 , \34216 );
and \U$33875 ( \34218 , \34046 , \34215 );
nor \U$33876 ( \34219 , \34217 , \34218 );
or \U$33877 ( \34220 , \34105 , \34103 );
nand \U$33878 ( \34221 , \34220 , \34106 );
xor \U$33879 ( \34222 , \34135 , \34155 );
xor \U$33880 ( \34223 , \34222 , \34184 );
and \U$33881 ( \34224 , \34221 , \34223 );
xor \U$33882 ( \34225 , \34194 , \34196 );
xor \U$33883 ( \34226 , \34225 , \34199 );
xor \U$33884 ( \34227 , \34135 , \34155 );
xor \U$33885 ( \34228 , \34227 , \34184 );
and \U$33886 ( \34229 , \34226 , \34228 );
and \U$33887 ( \34230 , \34221 , \34226 );
or \U$33888 ( \34231 , \34224 , \34229 , \34230 );
nand \U$33889 ( \34232 , RI986f0e8_44, RI9871fc8_144);
nand \U$33890 ( \34233 , RI986eff8_42, RI9871fc8_144);
xor \U$33891 ( \34234 , \34232 , \34233 );
and \U$33892 ( \34235 , \395 , RI986e4b8_18);
and \U$33893 ( \34236 , RI986e788_24, \393 );
nor \U$33894 ( \34237 , \34235 , \34236 );
not \U$33895 ( \34238 , \34237 );
not \U$33896 ( \34239 , \386 );
and \U$33897 ( \34240 , \34238 , \34239 );
and \U$33898 ( \34241 , \34237 , \487 );
nor \U$33899 ( \34242 , \34240 , \34241 );
not \U$33900 ( \34243 , \34242 );
and \U$33901 ( \34244 , \416 , RI986eff8_42);
and \U$33902 ( \34245 , RI986f2c8_48, \414 );
nor \U$33903 ( \34246 , \34244 , \34245 );
and \U$33904 ( \34247 , \34246 , \421 );
not \U$33905 ( \34248 , \34246 );
and \U$33906 ( \34249 , \34248 , \422 );
nor \U$33907 ( \34250 , \34247 , \34249 );
not \U$33908 ( \34251 , \34250 );
and \U$33909 ( \34252 , \34243 , \34251 );
and \U$33910 ( \34253 , \34242 , \34250 );
and \U$33911 ( \34254 , \354 , RI986f1d8_46);
and \U$33912 ( \34255 , RI986e5a8_20, \352 );
nor \U$33913 ( \34256 , \34254 , \34255 );
not \U$33914 ( \34257 , \34256 );
not \U$33915 ( \34258 , \345 );
and \U$33916 ( \34259 , \34257 , \34258 );
and \U$33917 ( \34260 , \34256 , \345 );
nor \U$33918 ( \34261 , \34259 , \34260 );
nor \U$33919 ( \34262 , \34253 , \34261 );
nor \U$33920 ( \34263 , \34252 , \34262 );
and \U$33921 ( \34264 , \34234 , \34263 );
and \U$33922 ( \34265 , \34232 , \34233 );
or \U$33923 ( \34266 , \34264 , \34265 );
and \U$33924 ( \34267 , \1311 , RI986dd38_2);
and \U$33925 ( \34268 , RI986e1e8_12, \1309 );
nor \U$33926 ( \34269 , \34267 , \34268 );
and \U$33927 ( \34270 , \34269 , \1315 );
not \U$33928 ( \34271 , \34269 );
and \U$33929 ( \34272 , \34271 , \1458 );
nor \U$33930 ( \34273 , \34270 , \34272 );
not \U$33931 ( \34274 , \34273 );
and \U$33932 ( \34275 , \2042 , RI986e0f8_10);
and \U$33933 ( \34276 , RI986e2d8_14, \2040 );
nor \U$33934 ( \34277 , \34275 , \34276 );
not \U$33935 ( \34278 , \34277 );
not \U$33936 ( \34279 , \1462 );
and \U$33937 ( \34280 , \34278 , \34279 );
and \U$33938 ( \34281 , \34277 , \2034 );
nor \U$33939 ( \34282 , \34280 , \34281 );
not \U$33940 ( \34283 , \34282 );
and \U$33941 ( \34284 , \34274 , \34283 );
and \U$33942 ( \34285 , \34282 , \34273 );
nand \U$33943 ( \34286 , RI986e3c8_16, \2274 );
and \U$33944 ( \34287 , \34286 , \2031 );
not \U$33945 ( \34288 , \34286 );
and \U$33946 ( \34289 , \34288 , \2030 );
nor \U$33947 ( \34290 , \34287 , \34289 );
nor \U$33948 ( \34291 , \34285 , \34290 );
nor \U$33949 ( \34292 , \34284 , \34291 );
and \U$33950 ( \34293 , \438 , RI986f958_62);
and \U$33951 ( \34294 , RI986f4a8_52, \436 );
nor \U$33952 ( \34295 , \34293 , \34294 );
and \U$33953 ( \34296 , \34295 , \443 );
not \U$33954 ( \34297 , \34295 );
and \U$33955 ( \34298 , \34297 , \444 );
nor \U$33956 ( \34299 , \34296 , \34298 );
not \U$33957 ( \34300 , \34299 );
and \U$33958 ( \34301 , \376 , RI986e698_22);
and \U$33959 ( \34302 , RI986f868_60, \374 );
nor \U$33960 ( \34303 , \34301 , \34302 );
not \U$33961 ( \34304 , \34303 );
not \U$33962 ( \34305 , \365 );
and \U$33963 ( \34306 , \34304 , \34305 );
and \U$33964 ( \34307 , \34303 , \367 );
nor \U$33965 ( \34308 , \34306 , \34307 );
not \U$33966 ( \34309 , \34308 );
and \U$33967 ( \34310 , \34300 , \34309 );
and \U$33968 ( \34311 , \34299 , \34308 );
and \U$33969 ( \34312 , \465 , RI986f778_58);
and \U$33970 ( \34313 , RI986fa48_64, \463 );
nor \U$33971 ( \34314 , \34312 , \34313 );
not \U$33972 ( \34315 , \34314 );
not \U$33973 ( \34316 , \454 );
and \U$33974 ( \34317 , \34315 , \34316 );
and \U$33975 ( \34318 , \34314 , \456 );
nor \U$33976 ( \34319 , \34317 , \34318 );
nor \U$33977 ( \34320 , \34311 , \34319 );
nor \U$33978 ( \34321 , \34310 , \34320 );
xor \U$33979 ( \34322 , \34292 , \34321 );
not \U$33980 ( \34323 , \1128 );
and \U$33981 ( \34324 , \1293 , RI986f688_56);
and \U$33982 ( \34325 , RI986e008_8, \1291 );
nor \U$33983 ( \34326 , \34324 , \34325 );
not \U$33984 ( \34327 , \34326 );
or \U$33985 ( \34328 , \34323 , \34327 );
or \U$33986 ( \34329 , \34326 , \1128 );
nand \U$33987 ( \34330 , \34328 , \34329 );
and \U$33988 ( \34331 , \1329 , RI986df18_6);
and \U$33989 ( \34332 , RI986de28_4, \1327 );
nor \U$33990 ( \34333 , \34331 , \34332 );
and \U$33991 ( \34334 , \34333 , \1336 );
not \U$33992 ( \34335 , \34333 );
and \U$33993 ( \34336 , \34335 , \1337 );
nor \U$33994 ( \34337 , \34334 , \34336 );
xor \U$33995 ( \34338 , \34330 , \34337 );
and \U$33996 ( \34339 , \776 , RI986f3b8_50);
and \U$33997 ( \34340 , RI986f598_54, \774 );
nor \U$33998 ( \34341 , \34339 , \34340 );
and \U$33999 ( \34342 , \34341 , \474 );
not \U$34000 ( \34343 , \34341 );
and \U$34001 ( \34344 , \34343 , \451 );
nor \U$34002 ( \34345 , \34342 , \34344 );
and \U$34003 ( \34346 , \34338 , \34345 );
and \U$34004 ( \34347 , \34330 , \34337 );
nor \U$34005 ( \34348 , \34346 , \34347 );
and \U$34006 ( \34349 , \34322 , \34348 );
and \U$34007 ( \34350 , \34292 , \34321 );
or \U$34008 ( \34351 , \34349 , \34350 );
xor \U$34009 ( \34352 , \34266 , \34351 );
not \U$34010 ( \34353 , \34114 );
not \U$34011 ( \34354 , \34133 );
or \U$34012 ( \34355 , \34353 , \34354 );
or \U$34013 ( \34356 , \34114 , \34133 );
nand \U$34014 ( \34357 , \34355 , \34356 );
not \U$34015 ( \34358 , \34357 );
not \U$34016 ( \34359 , \34122 );
and \U$34017 ( \34360 , \34358 , \34359 );
and \U$34018 ( \34361 , \34357 , \34122 );
nor \U$34019 ( \34362 , \34360 , \34361 );
xor \U$34020 ( \34363 , \34084 , \34092 );
xor \U$34021 ( \34364 , \34363 , \34100 );
xor \U$34022 ( \34365 , \34362 , \34364 );
not \U$34023 ( \34366 , \34171 );
not \U$34024 ( \34367 , \34182 );
or \U$34025 ( \34368 , \34366 , \34367 );
or \U$34026 ( \34369 , \34171 , \34182 );
nand \U$34027 ( \34370 , \34368 , \34369 );
not \U$34028 ( \34371 , \34370 );
not \U$34029 ( \34372 , \34163 );
and \U$34030 ( \34373 , \34371 , \34372 );
and \U$34031 ( \34374 , \34370 , \34163 );
nor \U$34032 ( \34375 , \34373 , \34374 );
and \U$34033 ( \34376 , \34365 , \34375 );
and \U$34034 ( \34377 , \34362 , \34364 );
or \U$34035 ( \34378 , \34376 , \34377 );
and \U$34036 ( \34379 , \34352 , \34378 );
and \U$34037 ( \34380 , \34266 , \34351 );
nor \U$34038 ( \34381 , \34379 , \34380 );
xor \U$34039 ( \34382 , \34231 , \34381 );
not \U$34040 ( \34383 , \34067 );
xor \U$34041 ( \34384 , \34061 , \34074 );
not \U$34042 ( \34385 , \34384 );
or \U$34043 ( \34386 , \34383 , \34385 );
or \U$34044 ( \34387 , \34384 , \34067 );
nand \U$34045 ( \34388 , \34386 , \34387 );
and \U$34046 ( \34389 , \34382 , \34388 );
and \U$34047 ( \34390 , \34231 , \34381 );
nor \U$34048 ( \34391 , \34389 , \34390 );
xor \U$34049 ( \34392 , \33956 , \33966 );
xor \U$34050 ( \34393 , \34392 , \33997 );
xor \U$34051 ( \34394 , \34391 , \34393 );
xor \U$34052 ( \34395 , \34076 , \34205 );
xor \U$34053 ( \34396 , \34395 , \34210 );
and \U$34054 ( \34397 , \34394 , \34396 );
and \U$34055 ( \34398 , \34391 , \34393 );
or \U$34056 ( \34399 , \34397 , \34398 );
not \U$34057 ( \34400 , \34399 );
not \U$34058 ( \34401 , \34049 );
xor \U$34059 ( \34402 , \34056 , \34213 );
not \U$34060 ( \34403 , \34402 );
or \U$34061 ( \34404 , \34401 , \34403 );
or \U$34062 ( \34405 , \34402 , \34049 );
nand \U$34063 ( \34406 , \34404 , \34405 );
nand \U$34064 ( \34407 , \34400 , \34406 );
or \U$34065 ( \34408 , \34219 , \34407 );
xnor \U$34066 ( \34409 , \34407 , \34219 );
not \U$34067 ( \34410 , \34399 );
not \U$34068 ( \34411 , \34406 );
or \U$34069 ( \34412 , \34410 , \34411 );
or \U$34070 ( \34413 , \34406 , \34399 );
nand \U$34071 ( \34414 , \34412 , \34413 );
and \U$34072 ( \34415 , \376 , RI986e788_24);
and \U$34073 ( \34416 , RI986e698_22, \374 );
nor \U$34074 ( \34417 , \34415 , \34416 );
not \U$34075 ( \34418 , \34417 );
not \U$34076 ( \34419 , \367 );
and \U$34077 ( \34420 , \34418 , \34419 );
and \U$34078 ( \34421 , \34417 , \365 );
nor \U$34079 ( \34422 , \34420 , \34421 );
and \U$34080 ( \34423 , \395 , RI986e5a8_20);
and \U$34081 ( \34424 , RI986e4b8_18, \393 );
nor \U$34082 ( \34425 , \34423 , \34424 );
not \U$34083 ( \34426 , \34425 );
not \U$34084 ( \34427 , \487 );
and \U$34085 ( \34428 , \34426 , \34427 );
and \U$34086 ( \34429 , \34425 , \386 );
nor \U$34087 ( \34430 , \34428 , \34429 );
xor \U$34088 ( \34431 , \34422 , \34430 );
and \U$34089 ( \34432 , \354 , RI986f2c8_48);
and \U$34090 ( \34433 , RI986f1d8_46, \352 );
nor \U$34091 ( \34434 , \34432 , \34433 );
not \U$34092 ( \34435 , \34434 );
not \U$34093 ( \34436 , \345 );
and \U$34094 ( \34437 , \34435 , \34436 );
and \U$34095 ( \34438 , \34434 , \361 );
nor \U$34096 ( \34439 , \34437 , \34438 );
and \U$34097 ( \34440 , \34431 , \34439 );
and \U$34098 ( \34441 , \34422 , \34430 );
nor \U$34099 ( \34442 , \34440 , \34441 );
xor \U$34100 ( \34443 , \34442 , \34232 );
not \U$34101 ( \34444 , \34250 );
xor \U$34102 ( \34445 , \34242 , \34261 );
not \U$34103 ( \34446 , \34445 );
or \U$34104 ( \34447 , \34444 , \34446 );
or \U$34105 ( \34448 , \34445 , \34250 );
nand \U$34106 ( \34449 , \34447 , \34448 );
and \U$34107 ( \34450 , \34443 , \34449 );
and \U$34108 ( \34451 , \34442 , \34232 );
or \U$34109 ( \34452 , \34450 , \34451 );
and \U$34110 ( \34453 , \776 , RI986f4a8_52);
and \U$34111 ( \34454 , RI986f3b8_50, \774 );
nor \U$34112 ( \34455 , \34453 , \34454 );
and \U$34113 ( \34456 , \34455 , \451 );
not \U$34114 ( \34457 , \34455 );
and \U$34115 ( \34458 , \34457 , \474 );
nor \U$34116 ( \34459 , \34456 , \34458 );
and \U$34117 ( \34460 , \465 , RI986f868_60);
and \U$34118 ( \34461 , RI986f778_58, \463 );
nor \U$34119 ( \34462 , \34460 , \34461 );
not \U$34120 ( \34463 , \34462 );
not \U$34121 ( \34464 , \456 );
and \U$34122 ( \34465 , \34463 , \34464 );
and \U$34123 ( \34466 , \34462 , \456 );
nor \U$34124 ( \34467 , \34465 , \34466 );
or \U$34125 ( \34468 , \34459 , \34467 );
not \U$34126 ( \34469 , \34467 );
not \U$34127 ( \34470 , \34459 );
or \U$34128 ( \34471 , \34469 , \34470 );
and \U$34129 ( \34472 , \438 , RI986fa48_64);
and \U$34130 ( \34473 , RI986f958_62, \436 );
nor \U$34131 ( \34474 , \34472 , \34473 );
and \U$34132 ( \34475 , \34474 , \444 );
not \U$34133 ( \34476 , \34474 );
and \U$34134 ( \34477 , \34476 , \443 );
nor \U$34135 ( \34478 , \34475 , \34477 );
nand \U$34136 ( \34479 , \34471 , \34478 );
nand \U$34137 ( \34480 , \34468 , \34479 );
and \U$34138 ( \34481 , \2274 , RI986e2d8_14);
and \U$34139 ( \34482 , RI986e3c8_16, \2272 );
nor \U$34140 ( \34483 , \34481 , \34482 );
and \U$34141 ( \34484 , \34483 , \2031 );
not \U$34142 ( \34485 , \34483 );
and \U$34143 ( \34486 , \34485 , \2030 );
nor \U$34144 ( \34487 , \34484 , \34486 );
or \U$34145 ( \34488 , \34487 , \2263 );
and \U$34146 ( \34489 , \34487 , \2263 );
and \U$34147 ( \34490 , \2042 , RI986e1e8_12);
and \U$34148 ( \34491 , RI986e0f8_10, \2040 );
nor \U$34149 ( \34492 , \34490 , \34491 );
not \U$34150 ( \34493 , \34492 );
not \U$34151 ( \34494 , \1462 );
and \U$34152 ( \34495 , \34493 , \34494 );
and \U$34153 ( \34496 , \34492 , \2034 );
nor \U$34154 ( \34497 , \34495 , \34496 );
nor \U$34155 ( \34498 , \34489 , \34497 );
not \U$34156 ( \34499 , \34498 );
nand \U$34157 ( \34500 , \34488 , \34499 );
xor \U$34158 ( \34501 , \34480 , \34500 );
and \U$34159 ( \34502 , \1293 , RI986f598_54);
and \U$34160 ( \34503 , RI986f688_56, \1291 );
nor \U$34161 ( \34504 , \34502 , \34503 );
not \U$34162 ( \34505 , \34504 );
not \U$34163 ( \34506 , \1128 );
and \U$34164 ( \34507 , \34505 , \34506 );
and \U$34165 ( \34508 , \34504 , \1128 );
nor \U$34166 ( \34509 , \34507 , \34508 );
and \U$34167 ( \34510 , \1329 , RI986e008_8);
and \U$34168 ( \34511 , RI986df18_6, \1327 );
nor \U$34169 ( \34512 , \34510 , \34511 );
and \U$34170 ( \34513 , \34512 , \1337 );
not \U$34171 ( \34514 , \34512 );
and \U$34172 ( \34515 , \34514 , \1336 );
nor \U$34173 ( \34516 , \34513 , \34515 );
or \U$34174 ( \34517 , \34509 , \34516 );
not \U$34175 ( \34518 , \34516 );
not \U$34176 ( \34519 , \34509 );
or \U$34177 ( \34520 , \34518 , \34519 );
and \U$34178 ( \34521 , \1311 , RI986de28_4);
and \U$34179 ( \34522 , RI986dd38_2, \1309 );
nor \U$34180 ( \34523 , \34521 , \34522 );
and \U$34181 ( \34524 , \34523 , \1458 );
not \U$34182 ( \34525 , \34523 );
and \U$34183 ( \34526 , \34525 , \1318 );
nor \U$34184 ( \34527 , \34524 , \34526 );
nand \U$34185 ( \34528 , \34520 , \34527 );
nand \U$34186 ( \34529 , \34517 , \34528 );
and \U$34187 ( \34530 , \34501 , \34529 );
and \U$34188 ( \34531 , \34480 , \34500 );
or \U$34189 ( \34532 , \34530 , \34531 );
xor \U$34190 ( \34533 , \34452 , \34532 );
xor \U$34191 ( \34534 , \34330 , \34337 );
xor \U$34192 ( \34535 , \34534 , \34345 );
not \U$34193 ( \34536 , \34273 );
xor \U$34194 ( \34537 , \34290 , \34282 );
not \U$34195 ( \34538 , \34537 );
or \U$34196 ( \34539 , \34536 , \34538 );
or \U$34197 ( \34540 , \34537 , \34273 );
nand \U$34198 ( \34541 , \34539 , \34540 );
xor \U$34199 ( \34542 , \34535 , \34541 );
not \U$34200 ( \34543 , \34308 );
xor \U$34201 ( \34544 , \34319 , \34299 );
not \U$34202 ( \34545 , \34544 );
or \U$34203 ( \34546 , \34543 , \34545 );
or \U$34204 ( \34547 , \34544 , \34308 );
nand \U$34205 ( \34548 , \34546 , \34547 );
and \U$34206 ( \34549 , \34542 , \34548 );
and \U$34207 ( \34550 , \34535 , \34541 );
or \U$34208 ( \34551 , \34549 , \34550 );
and \U$34209 ( \34552 , \34533 , \34551 );
and \U$34210 ( \34553 , \34452 , \34532 );
or \U$34211 ( \34554 , \34552 , \34553 );
and \U$34212 ( \34555 , \34143 , \2031 );
not \U$34213 ( \34556 , \34143 );
and \U$34214 ( \34557 , \34556 , \2030 );
nor \U$34215 ( \34558 , \34555 , \34557 );
not \U$34216 ( \34559 , \34558 );
not \U$34217 ( \34560 , \34152 );
and \U$34218 ( \34561 , \34559 , \34560 );
and \U$34219 ( \34562 , \34558 , \34152 );
nor \U$34220 ( \34563 , \34561 , \34562 );
xor \U$34221 ( \34564 , \34232 , \34233 );
xor \U$34222 ( \34565 , \34564 , \34263 );
xor \U$34223 ( \34566 , \34563 , \34565 );
xor \U$34224 ( \34567 , \34362 , \34364 );
xor \U$34225 ( \34568 , \34567 , \34375 );
and \U$34226 ( \34569 , \34566 , \34568 );
and \U$34227 ( \34570 , \34563 , \34565 );
nor \U$34228 ( \34571 , \34569 , \34570 );
xor \U$34229 ( \34572 , \34554 , \34571 );
xor \U$34230 ( \34573 , \34135 , \34155 );
xor \U$34231 ( \34574 , \34573 , \34184 );
xor \U$34232 ( \34575 , \34221 , \34226 );
xor \U$34233 ( \34576 , \34574 , \34575 );
and \U$34234 ( \34577 , \34572 , \34576 );
and \U$34235 ( \34578 , \34554 , \34571 );
or \U$34236 ( \34579 , \34577 , \34578 );
xor \U$34237 ( \34580 , \34106 , \34187 );
xor \U$34238 ( \34581 , \34580 , \34202 );
xor \U$34239 ( \34582 , \34579 , \34581 );
xor \U$34240 ( \34583 , \34231 , \34381 );
xor \U$34241 ( \34584 , \34583 , \34388 );
and \U$34242 ( \34585 , \34582 , \34584 );
and \U$34243 ( \34586 , \34579 , \34581 );
or \U$34244 ( \34587 , \34585 , \34586 );
not \U$34245 ( \34588 , \34587 );
xor \U$34246 ( \34589 , \34391 , \34393 );
xor \U$34247 ( \34590 , \34589 , \34396 );
nor \U$34248 ( \34591 , \34588 , \34590 );
and \U$34249 ( \34592 , \34414 , \34591 );
xor \U$34250 ( \34593 , \34591 , \34414 );
xor \U$34251 ( \34594 , \34563 , \34565 );
xor \U$34252 ( \34595 , \34594 , \34568 );
not \U$34253 ( \34596 , \34595 );
xor \U$34254 ( \34597 , \34452 , \34532 );
xor \U$34255 ( \34598 , \34597 , \34551 );
nand \U$34256 ( \34599 , \34596 , \34598 );
xor \U$34257 ( \34600 , \34266 , \34351 );
xor \U$34258 ( \34601 , \34600 , \34378 );
xor \U$34259 ( \34602 , \34599 , \34601 );
xor \U$34260 ( \34603 , \34535 , \34541 );
xor \U$34261 ( \34604 , \34603 , \34548 );
xor \U$34262 ( \34605 , \34480 , \34500 );
xor \U$34263 ( \34606 , \34605 , \34529 );
xor \U$34264 ( \34607 , \34604 , \34606 );
xor \U$34265 ( \34608 , \34442 , \34232 );
xor \U$34266 ( \34609 , \34608 , \34449 );
and \U$34267 ( \34610 , \34607 , \34609 );
and \U$34268 ( \34611 , \34604 , \34606 );
nor \U$34269 ( \34612 , \34610 , \34611 );
not \U$34270 ( \34613 , \34612 );
xor \U$34271 ( \34614 , \34292 , \34321 );
xor \U$34272 ( \34615 , \34614 , \34348 );
not \U$34273 ( \34616 , \34615 );
and \U$34274 ( \34617 , \34613 , \34616 );
and \U$34275 ( \34618 , \34612 , \34615 );
and \U$34276 ( \34619 , \2042 , RI986dd38_2);
and \U$34277 ( \34620 , RI986e1e8_12, \2040 );
nor \U$34278 ( \34621 , \34619 , \34620 );
not \U$34279 ( \34622 , \34621 );
not \U$34280 ( \34623 , \1462 );
and \U$34281 ( \34624 , \34622 , \34623 );
and \U$34282 ( \34625 , \34621 , \2034 );
nor \U$34283 ( \34626 , \34624 , \34625 );
not \U$34284 ( \34627 , \34626 );
and \U$34285 ( \34628 , \2274 , RI986e0f8_10);
and \U$34286 ( \34629 , RI986e2d8_14, \2272 );
nor \U$34287 ( \34630 , \34628 , \34629 );
and \U$34288 ( \34631 , \34630 , \2031 );
not \U$34289 ( \34632 , \34630 );
and \U$34290 ( \34633 , \34632 , \2030 );
nor \U$34291 ( \34634 , \34631 , \34633 );
not \U$34292 ( \34635 , \34634 );
and \U$34293 ( \34636 , \34627 , \34635 );
and \U$34294 ( \34637 , \34634 , \34626 );
nand \U$34295 ( \34638 , RI986e3c8_16, \2464 );
and \U$34296 ( \34639 , \34638 , \2263 );
not \U$34297 ( \34640 , \34638 );
and \U$34298 ( \34641 , \34640 , \2468 );
nor \U$34299 ( \34642 , \34639 , \34641 );
nor \U$34300 ( \34643 , \34637 , \34642 );
nor \U$34301 ( \34644 , \34636 , \34643 );
and \U$34302 ( \34645 , \776 , RI986f958_62);
and \U$34303 ( \34646 , RI986f4a8_52, \774 );
nor \U$34304 ( \34647 , \34645 , \34646 );
and \U$34305 ( \34648 , \34647 , \474 );
not \U$34306 ( \34649 , \34647 );
and \U$34307 ( \34650 , \34649 , \451 );
nor \U$34308 ( \34651 , \34648 , \34650 );
and \U$34309 ( \34652 , \438 , RI986f778_58);
and \U$34310 ( \34653 , RI986fa48_64, \436 );
nor \U$34311 ( \34654 , \34652 , \34653 );
and \U$34312 ( \34655 , \34654 , \444 );
not \U$34313 ( \34656 , \34654 );
and \U$34314 ( \34657 , \34656 , \443 );
nor \U$34315 ( \34658 , \34655 , \34657 );
xor \U$34316 ( \34659 , \34651 , \34658 );
not \U$34317 ( \34660 , \456 );
and \U$34318 ( \34661 , \465 , RI986e698_22);
and \U$34319 ( \34662 , RI986f868_60, \463 );
nor \U$34320 ( \34663 , \34661 , \34662 );
not \U$34321 ( \34664 , \34663 );
or \U$34322 ( \34665 , \34660 , \34664 );
or \U$34323 ( \34666 , \34663 , \454 );
nand \U$34324 ( \34667 , \34665 , \34666 );
and \U$34325 ( \34668 , \34659 , \34667 );
and \U$34326 ( \34669 , \34651 , \34658 );
nor \U$34327 ( \34670 , \34668 , \34669 );
or \U$34328 ( \34671 , \34644 , \34670 );
not \U$34329 ( \34672 , \34644 );
not \U$34330 ( \34673 , \34670 );
or \U$34331 ( \34674 , \34672 , \34673 );
and \U$34332 ( \34675 , \1311 , RI986df18_6);
and \U$34333 ( \34676 , RI986de28_4, \1309 );
nor \U$34334 ( \34677 , \34675 , \34676 );
and \U$34335 ( \34678 , \34677 , \1458 );
not \U$34336 ( \34679 , \34677 );
and \U$34337 ( \34680 , \34679 , \1315 );
nor \U$34338 ( \34681 , \34678 , \34680 );
not \U$34339 ( \34682 , \1301 );
and \U$34340 ( \34683 , \1293 , RI986f3b8_50);
and \U$34341 ( \34684 , RI986f598_54, \1291 );
nor \U$34342 ( \34685 , \34683 , \34684 );
not \U$34343 ( \34686 , \34685 );
or \U$34344 ( \34687 , \34682 , \34686 );
or \U$34345 ( \34688 , \34685 , \1301 );
nand \U$34346 ( \34689 , \34687 , \34688 );
xor \U$34347 ( \34690 , \34681 , \34689 );
and \U$34348 ( \34691 , \1329 , RI986f688_56);
and \U$34349 ( \34692 , RI986e008_8, \1327 );
nor \U$34350 ( \34693 , \34691 , \34692 );
and \U$34351 ( \34694 , \34693 , \1336 );
not \U$34352 ( \34695 , \34693 );
and \U$34353 ( \34696 , \34695 , \1337 );
nor \U$34354 ( \34697 , \34694 , \34696 );
and \U$34355 ( \34698 , \34690 , \34697 );
and \U$34356 ( \34699 , \34681 , \34689 );
or \U$34357 ( \34700 , \34698 , \34699 );
nand \U$34358 ( \34701 , \34674 , \34700 );
nand \U$34359 ( \34702 , \34671 , \34701 );
nand \U$34360 ( \34703 , RI986ec38_34, RI9871fc8_144);
and \U$34361 ( \34704 , \416 , RI986ed28_36);
and \U$34362 ( \34705 , RI986f0e8_44, \414 );
nor \U$34363 ( \34706 , \34704 , \34705 );
and \U$34364 ( \34707 , \34706 , \421 );
not \U$34365 ( \34708 , \34706 );
and \U$34366 ( \34709 , \34708 , \422 );
nor \U$34367 ( \34710 , \34707 , \34709 );
nand \U$34368 ( \34711 , \34703 , \34710 );
and \U$34369 ( \34712 , \416 , RI986f0e8_44);
and \U$34370 ( \34713 , RI986eff8_42, \414 );
nor \U$34371 ( \34714 , \34712 , \34713 );
and \U$34372 ( \34715 , \34714 , \422 );
not \U$34373 ( \34716 , \34714 );
and \U$34374 ( \34717 , \34716 , \421 );
nor \U$34375 ( \34718 , \34715 , \34717 );
xor \U$34376 ( \34719 , \34711 , \34718 );
not \U$34377 ( \34720 , \365 );
and \U$34378 ( \34721 , \376 , RI986e4b8_18);
and \U$34379 ( \34722 , RI986e788_24, \374 );
nor \U$34380 ( \34723 , \34721 , \34722 );
not \U$34381 ( \34724 , \34723 );
or \U$34382 ( \34725 , \34720 , \34724 );
or \U$34383 ( \34726 , \34723 , \365 );
nand \U$34384 ( \34727 , \34725 , \34726 );
not \U$34385 ( \34728 , \386 );
and \U$34386 ( \34729 , \395 , RI986f1d8_46);
and \U$34387 ( \34730 , RI986e5a8_20, \393 );
nor \U$34388 ( \34731 , \34729 , \34730 );
not \U$34389 ( \34732 , \34731 );
or \U$34390 ( \34733 , \34728 , \34732 );
or \U$34391 ( \34734 , \34731 , \487 );
nand \U$34392 ( \34735 , \34733 , \34734 );
xor \U$34393 ( \34736 , \34727 , \34735 );
not \U$34394 ( \34737 , \361 );
and \U$34395 ( \34738 , \354 , RI986eff8_42);
and \U$34396 ( \34739 , RI986f2c8_48, \352 );
nor \U$34397 ( \34740 , \34738 , \34739 );
not \U$34398 ( \34741 , \34740 );
or \U$34399 ( \34742 , \34737 , \34741 );
or \U$34400 ( \34743 , \34740 , \361 );
nand \U$34401 ( \34744 , \34742 , \34743 );
and \U$34402 ( \34745 , \34736 , \34744 );
and \U$34403 ( \34746 , \34727 , \34735 );
or \U$34404 ( \34747 , \34745 , \34746 );
and \U$34405 ( \34748 , \34719 , \34747 );
and \U$34406 ( \34749 , \34711 , \34718 );
or \U$34407 ( \34750 , \34748 , \34749 );
and \U$34408 ( \34751 , \34702 , \34750 );
not \U$34409 ( \34752 , \34702 );
not \U$34410 ( \34753 , \34750 );
and \U$34411 ( \34754 , \34752 , \34753 );
not \U$34412 ( \34755 , \34459 );
not \U$34413 ( \34756 , \34478 );
or \U$34414 ( \34757 , \34755 , \34756 );
or \U$34415 ( \34758 , \34459 , \34478 );
nand \U$34416 ( \34759 , \34757 , \34758 );
not \U$34417 ( \34760 , \34759 );
not \U$34418 ( \34761 , \34467 );
and \U$34419 ( \34762 , \34760 , \34761 );
and \U$34420 ( \34763 , \34759 , \34467 );
nor \U$34421 ( \34764 , \34762 , \34763 );
nand \U$34422 ( \34765 , RI986ed28_36, RI9871fc8_144);
xor \U$34423 ( \34766 , \34764 , \34765 );
xor \U$34424 ( \34767 , \34422 , \34430 );
xor \U$34425 ( \34768 , \34767 , \34439 );
and \U$34426 ( \34769 , \34766 , \34768 );
and \U$34427 ( \34770 , \34764 , \34765 );
or \U$34428 ( \34771 , \34769 , \34770 );
nor \U$34429 ( \34772 , \34754 , \34771 );
nor \U$34430 ( \34773 , \34751 , \34772 );
nor \U$34431 ( \34774 , \34618 , \34773 );
nor \U$34432 ( \34775 , \34617 , \34774 );
and \U$34433 ( \34776 , \34602 , \34775 );
and \U$34434 ( \34777 , \34599 , \34601 );
or \U$34435 ( \34778 , \34776 , \34777 );
not \U$34436 ( \34779 , \34778 );
xor \U$34437 ( \34780 , \34579 , \34581 );
xor \U$34438 ( \34781 , \34780 , \34584 );
nand \U$34439 ( \34782 , \34779 , \34781 );
not \U$34440 ( \34783 , \34590 );
not \U$34441 ( \34784 , \34587 );
and \U$34442 ( \34785 , \34783 , \34784 );
and \U$34443 ( \34786 , \34590 , \34587 );
nor \U$34444 ( \34787 , \34785 , \34786 );
xor \U$34445 ( \34788 , \34782 , \34787 );
and \U$34446 ( \34789 , \2464 , RI986e2d8_14);
and \U$34447 ( \34790 , RI986e3c8_16, \2462 );
nor \U$34448 ( \34791 , \34789 , \34790 );
and \U$34449 ( \34792 , \34791 , \2263 );
not \U$34450 ( \34793 , \34791 );
and \U$34451 ( \34794 , \34793 , \2468 );
nor \U$34452 ( \34795 , \34792 , \34794 );
xor \U$34453 ( \34796 , \34795 , \3406 );
and \U$34454 ( \34797 , \2274 , RI986e1e8_12);
and \U$34455 ( \34798 , RI986e0f8_10, \2272 );
nor \U$34456 ( \34799 , \34797 , \34798 );
and \U$34457 ( \34800 , \34799 , \2031 );
not \U$34458 ( \34801 , \34799 );
and \U$34459 ( \34802 , \34801 , \2030 );
nor \U$34460 ( \34803 , \34800 , \34802 );
and \U$34461 ( \34804 , \34796 , \34803 );
and \U$34462 ( \34805 , \34795 , \3406 );
or \U$34463 ( \34806 , \34804 , \34805 );
and \U$34464 ( \34807 , \1329 , RI986f598_54);
and \U$34465 ( \34808 , RI986f688_56, \1327 );
nor \U$34466 ( \34809 , \34807 , \34808 );
and \U$34467 ( \34810 , \34809 , \1337 );
not \U$34468 ( \34811 , \34809 );
and \U$34469 ( \34812 , \34811 , \1336 );
nor \U$34470 ( \34813 , \34810 , \34812 );
not \U$34471 ( \34814 , \34813 );
and \U$34472 ( \34815 , \1311 , RI986e008_8);
and \U$34473 ( \34816 , RI986df18_6, \1309 );
nor \U$34474 ( \34817 , \34815 , \34816 );
and \U$34475 ( \34818 , \34817 , \1315 );
not \U$34476 ( \34819 , \34817 );
and \U$34477 ( \34820 , \34819 , \1458 );
nor \U$34478 ( \34821 , \34818 , \34820 );
not \U$34479 ( \34822 , \34821 );
and \U$34480 ( \34823 , \34814 , \34822 );
and \U$34481 ( \34824 , \34821 , \34813 );
and \U$34482 ( \34825 , \2042 , RI986de28_4);
and \U$34483 ( \34826 , RI986dd38_2, \2040 );
nor \U$34484 ( \34827 , \34825 , \34826 );
not \U$34485 ( \34828 , \34827 );
not \U$34486 ( \34829 , \2034 );
and \U$34487 ( \34830 , \34828 , \34829 );
and \U$34488 ( \34831 , \34827 , \1462 );
nor \U$34489 ( \34832 , \34830 , \34831 );
nor \U$34490 ( \34833 , \34824 , \34832 );
nor \U$34491 ( \34834 , \34823 , \34833 );
xor \U$34492 ( \34835 , \34806 , \34834 );
and \U$34493 ( \34836 , \1293 , RI986f4a8_52);
and \U$34494 ( \34837 , RI986f3b8_50, \1291 );
nor \U$34495 ( \34838 , \34836 , \34837 );
not \U$34496 ( \34839 , \34838 );
not \U$34497 ( \34840 , \1301 );
and \U$34498 ( \34841 , \34839 , \34840 );
and \U$34499 ( \34842 , \34838 , \1301 );
nor \U$34500 ( \34843 , \34841 , \34842 );
and \U$34501 ( \34844 , \776 , RI986fa48_64);
and \U$34502 ( \34845 , RI986f958_62, \774 );
nor \U$34503 ( \34846 , \34844 , \34845 );
and \U$34504 ( \34847 , \34846 , \451 );
not \U$34505 ( \34848 , \34846 );
and \U$34506 ( \34849 , \34848 , \474 );
nor \U$34507 ( \34850 , \34847 , \34849 );
xor \U$34508 ( \34851 , \34843 , \34850 );
and \U$34509 ( \34852 , \438 , RI986f868_60);
and \U$34510 ( \34853 , RI986f778_58, \436 );
nor \U$34511 ( \34854 , \34852 , \34853 );
and \U$34512 ( \34855 , \34854 , \443 );
not \U$34513 ( \34856 , \34854 );
and \U$34514 ( \34857 , \34856 , \444 );
nor \U$34515 ( \34858 , \34855 , \34857 );
and \U$34516 ( \34859 , \34851 , \34858 );
and \U$34517 ( \34860 , \34843 , \34850 );
or \U$34518 ( \34861 , \34859 , \34860 );
and \U$34519 ( \34862 , \34835 , \34861 );
and \U$34520 ( \34863 , \34806 , \34834 );
nor \U$34521 ( \34864 , \34862 , \34863 );
and \U$34522 ( \34865 , \416 , RI986ec38_34);
and \U$34523 ( \34866 , RI986ed28_36, \414 );
nor \U$34524 ( \34867 , \34865 , \34866 );
and \U$34525 ( \34868 , \34867 , \421 );
not \U$34526 ( \34869 , \34867 );
and \U$34527 ( \34870 , \34869 , \422 );
nor \U$34528 ( \34871 , \34868 , \34870 );
nand \U$34529 ( \34872 , RI986ee18_38, RI9871fc8_144);
or \U$34530 ( \34873 , \34871 , \34872 );
not \U$34531 ( \34874 , \34872 );
not \U$34532 ( \34875 , \34871 );
or \U$34533 ( \34876 , \34874 , \34875 );
not \U$34534 ( \34877 , \361 );
and \U$34535 ( \34878 , \354 , RI986f0e8_44);
and \U$34536 ( \34879 , RI986eff8_42, \352 );
nor \U$34537 ( \34880 , \34878 , \34879 );
not \U$34538 ( \34881 , \34880 );
or \U$34539 ( \34882 , \34877 , \34881 );
or \U$34540 ( \34883 , \34880 , \345 );
nand \U$34541 ( \34884 , \34882 , \34883 );
nand \U$34542 ( \34885 , \34876 , \34884 );
nand \U$34543 ( \34886 , \34873 , \34885 );
or \U$34544 ( \34887 , \34710 , \34703 );
nand \U$34545 ( \34888 , \34887 , \34711 );
xor \U$34546 ( \34889 , \34886 , \34888 );
and \U$34547 ( \34890 , \465 , RI986e788_24);
and \U$34548 ( \34891 , RI986e698_22, \463 );
nor \U$34549 ( \34892 , \34890 , \34891 );
not \U$34550 ( \34893 , \34892 );
not \U$34551 ( \34894 , \456 );
and \U$34552 ( \34895 , \34893 , \34894 );
and \U$34553 ( \34896 , \34892 , \454 );
nor \U$34554 ( \34897 , \34895 , \34896 );
and \U$34555 ( \34898 , \395 , RI986f2c8_48);
and \U$34556 ( \34899 , RI986f1d8_46, \393 );
nor \U$34557 ( \34900 , \34898 , \34899 );
not \U$34558 ( \34901 , \34900 );
not \U$34559 ( \34902 , \487 );
and \U$34560 ( \34903 , \34901 , \34902 );
and \U$34561 ( \34904 , \34900 , \487 );
nor \U$34562 ( \34905 , \34903 , \34904 );
or \U$34563 ( \34906 , \34897 , \34905 );
not \U$34564 ( \34907 , \34905 );
not \U$34565 ( \34908 , \34897 );
or \U$34566 ( \34909 , \34907 , \34908 );
not \U$34567 ( \34910 , \365 );
and \U$34568 ( \34911 , \376 , RI986e5a8_20);
and \U$34569 ( \34912 , RI986e4b8_18, \374 );
nor \U$34570 ( \34913 , \34911 , \34912 );
not \U$34571 ( \34914 , \34913 );
or \U$34572 ( \34915 , \34910 , \34914 );
or \U$34573 ( \34916 , \34913 , \365 );
nand \U$34574 ( \34917 , \34915 , \34916 );
nand \U$34575 ( \34918 , \34909 , \34917 );
nand \U$34576 ( \34919 , \34906 , \34918 );
and \U$34577 ( \34920 , \34889 , \34919 );
and \U$34578 ( \34921 , \34886 , \34888 );
or \U$34579 ( \34922 , \34920 , \34921 );
xor \U$34580 ( \34923 , \34864 , \34922 );
xor \U$34581 ( \34924 , \34651 , \34658 );
xor \U$34582 ( \34925 , \34924 , \34667 );
xor \U$34583 ( \34926 , \34727 , \34735 );
xor \U$34584 ( \34927 , \34926 , \34744 );
and \U$34585 ( \34928 , \34925 , \34927 );
xor \U$34586 ( \34929 , \34681 , \34689 );
xor \U$34587 ( \34930 , \34929 , \34697 );
xor \U$34588 ( \34931 , \34727 , \34735 );
xor \U$34589 ( \34932 , \34931 , \34744 );
and \U$34590 ( \34933 , \34930 , \34932 );
and \U$34591 ( \34934 , \34925 , \34930 );
or \U$34592 ( \34935 , \34928 , \34933 , \34934 );
and \U$34593 ( \34936 , \34923 , \34935 );
and \U$34594 ( \34937 , \34864 , \34922 );
or \U$34595 ( \34938 , \34936 , \34937 );
and \U$34596 ( \34939 , \34487 , \2263 );
not \U$34597 ( \34940 , \34487 );
and \U$34598 ( \34941 , \34940 , \2468 );
nor \U$34599 ( \34942 , \34939 , \34941 );
not \U$34600 ( \34943 , \34942 );
not \U$34601 ( \34944 , \34497 );
and \U$34602 ( \34945 , \34943 , \34944 );
and \U$34603 ( \34946 , \34942 , \34497 );
nor \U$34604 ( \34947 , \34945 , \34946 );
not \U$34605 ( \34948 , \34516 );
not \U$34606 ( \34949 , \34527 );
or \U$34607 ( \34950 , \34948 , \34949 );
or \U$34608 ( \34951 , \34516 , \34527 );
nand \U$34609 ( \34952 , \34950 , \34951 );
not \U$34610 ( \34953 , \34952 );
not \U$34611 ( \34954 , \34509 );
and \U$34612 ( \34955 , \34953 , \34954 );
and \U$34613 ( \34956 , \34952 , \34509 );
nor \U$34614 ( \34957 , \34955 , \34956 );
or \U$34615 ( \34958 , \34947 , \34957 );
and \U$34616 ( \34959 , \34947 , \34957 );
xor \U$34617 ( \34960 , \34764 , \34765 );
xor \U$34618 ( \34961 , \34960 , \34768 );
nor \U$34619 ( \34962 , \34959 , \34961 );
not \U$34620 ( \34963 , \34962 );
nand \U$34621 ( \34964 , \34958 , \34963 );
xor \U$34622 ( \34965 , \34938 , \34964 );
xor \U$34623 ( \34966 , \34604 , \34606 );
xor \U$34624 ( \34967 , \34966 , \34609 );
and \U$34625 ( \34968 , \34965 , \34967 );
and \U$34626 ( \34969 , \34938 , \34964 );
or \U$34627 ( \34970 , \34968 , \34969 );
not \U$34628 ( \34971 , \34595 );
not \U$34629 ( \34972 , \34598 );
or \U$34630 ( \34973 , \34971 , \34972 );
or \U$34631 ( \34974 , \34598 , \34595 );
nand \U$34632 ( \34975 , \34973 , \34974 );
xor \U$34633 ( \34976 , \34970 , \34975 );
not \U$34634 ( \34977 , \34615 );
xor \U$34635 ( \34978 , \34773 , \34612 );
not \U$34636 ( \34979 , \34978 );
or \U$34637 ( \34980 , \34977 , \34979 );
or \U$34638 ( \34981 , \34978 , \34615 );
nand \U$34639 ( \34982 , \34980 , \34981 );
xor \U$34640 ( \34983 , \34976 , \34982 );
xor \U$34641 ( \34984 , \34711 , \34718 );
xor \U$34642 ( \34985 , \34984 , \34747 );
not \U$34643 ( \34986 , \34985 );
not \U$34644 ( \34987 , \34871 );
not \U$34645 ( \34988 , \34884 );
or \U$34646 ( \34989 , \34987 , \34988 );
or \U$34647 ( \34990 , \34871 , \34884 );
nand \U$34648 ( \34991 , \34989 , \34990 );
not \U$34649 ( \34992 , \34991 );
not \U$34650 ( \34993 , \34872 );
and \U$34651 ( \34994 , \34992 , \34993 );
and \U$34652 ( \34995 , \34991 , \34872 );
nor \U$34653 ( \34996 , \34994 , \34995 );
and \U$34654 ( \34997 , \416 , RI986ee18_38);
and \U$34655 ( \34998 , RI986ec38_34, \414 );
nor \U$34656 ( \34999 , \34997 , \34998 );
and \U$34657 ( \35000 , \34999 , \421 );
not \U$34658 ( \35001 , \34999 );
and \U$34659 ( \35002 , \35001 , \422 );
nor \U$34660 ( \35003 , \35000 , \35002 );
nand \U$34661 ( \35004 , RI986ef08_40, RI9871fc8_144);
xor \U$34662 ( \35005 , \35003 , \35004 );
and \U$34663 ( \35006 , \354 , RI986ed28_36);
and \U$34664 ( \35007 , RI986f0e8_44, \352 );
nor \U$34665 ( \35008 , \35006 , \35007 );
not \U$34666 ( \35009 , \35008 );
not \U$34667 ( \35010 , \361 );
and \U$34668 ( \35011 , \35009 , \35010 );
and \U$34669 ( \35012 , \35008 , \361 );
nor \U$34670 ( \35013 , \35011 , \35012 );
and \U$34671 ( \35014 , \35005 , \35013 );
and \U$34672 ( \35015 , \35003 , \35004 );
or \U$34673 ( \35016 , \35014 , \35015 );
or \U$34674 ( \35017 , \34996 , \35016 );
not \U$34675 ( \35018 , \35016 );
not \U$34676 ( \35019 , \34996 );
or \U$34677 ( \35020 , \35018 , \35019 );
and \U$34678 ( \35021 , \376 , RI986f1d8_46);
and \U$34679 ( \35022 , RI986e5a8_20, \374 );
nor \U$34680 ( \35023 , \35021 , \35022 );
not \U$34681 ( \35024 , \35023 );
not \U$34682 ( \35025 , \365 );
and \U$34683 ( \35026 , \35024 , \35025 );
and \U$34684 ( \35027 , \35023 , \365 );
nor \U$34685 ( \35028 , \35026 , \35027 );
and \U$34686 ( \35029 , \395 , RI986eff8_42);
and \U$34687 ( \35030 , RI986f2c8_48, \393 );
nor \U$34688 ( \35031 , \35029 , \35030 );
not \U$34689 ( \35032 , \35031 );
not \U$34690 ( \35033 , \386 );
and \U$34691 ( \35034 , \35032 , \35033 );
and \U$34692 ( \35035 , \35031 , \487 );
nor \U$34693 ( \35036 , \35034 , \35035 );
or \U$34694 ( \35037 , \35028 , \35036 );
not \U$34695 ( \35038 , \35036 );
not \U$34696 ( \35039 , \35028 );
or \U$34697 ( \35040 , \35038 , \35039 );
not \U$34698 ( \35041 , \456 );
and \U$34699 ( \35042 , \465 , RI986e4b8_18);
and \U$34700 ( \35043 , RI986e788_24, \463 );
nor \U$34701 ( \35044 , \35042 , \35043 );
not \U$34702 ( \35045 , \35044 );
or \U$34703 ( \35046 , \35041 , \35045 );
or \U$34704 ( \35047 , \35044 , \454 );
nand \U$34705 ( \35048 , \35046 , \35047 );
nand \U$34706 ( \35049 , \35040 , \35048 );
nand \U$34707 ( \35050 , \35037 , \35049 );
nand \U$34708 ( \35051 , \35020 , \35050 );
nand \U$34709 ( \35052 , \35017 , \35051 );
and \U$34710 ( \35053 , \2274 , RI986dd38_2);
and \U$34711 ( \35054 , RI986e1e8_12, \2272 );
nor \U$34712 ( \35055 , \35053 , \35054 );
and \U$34713 ( \35056 , \35055 , \2031 );
not \U$34714 ( \35057 , \35055 );
and \U$34715 ( \35058 , \35057 , \2030 );
nor \U$34716 ( \35059 , \35056 , \35058 );
not \U$34717 ( \35060 , \35059 );
and \U$34718 ( \35061 , \2464 , RI986e0f8_10);
and \U$34719 ( \35062 , RI986e2d8_14, \2462 );
nor \U$34720 ( \35063 , \35061 , \35062 );
and \U$34721 ( \35064 , \35063 , \2263 );
not \U$34722 ( \35065 , \35063 );
and \U$34723 ( \35066 , \35065 , \2468 );
nor \U$34724 ( \35067 , \35064 , \35066 );
not \U$34725 ( \35068 , \35067 );
and \U$34726 ( \35069 , \35060 , \35068 );
and \U$34727 ( \35070 , \35067 , \35059 );
nand \U$34728 ( \35071 , RI986e3c8_16, \3254 );
not \U$34729 ( \35072 , \35071 );
not \U$34730 ( \35073 , \3406 );
and \U$34731 ( \35074 , \35072 , \35073 );
and \U$34732 ( \35075 , \35071 , \2935 );
nor \U$34733 ( \35076 , \35074 , \35075 );
nor \U$34734 ( \35077 , \35070 , \35076 );
nor \U$34735 ( \35078 , \35069 , \35077 );
and \U$34736 ( \35079 , \1329 , RI986f3b8_50);
and \U$34737 ( \35080 , RI986f598_54, \1327 );
nor \U$34738 ( \35081 , \35079 , \35080 );
and \U$34739 ( \35082 , \35081 , \1337 );
not \U$34740 ( \35083 , \35081 );
and \U$34741 ( \35084 , \35083 , \1336 );
nor \U$34742 ( \35085 , \35082 , \35084 );
not \U$34743 ( \35086 , \35085 );
and \U$34744 ( \35087 , \1311 , RI986f688_56);
and \U$34745 ( \35088 , RI986e008_8, \1309 );
nor \U$34746 ( \35089 , \35087 , \35088 );
and \U$34747 ( \35090 , \35089 , \1315 );
not \U$34748 ( \35091 , \35089 );
and \U$34749 ( \35092 , \35091 , \1458 );
nor \U$34750 ( \35093 , \35090 , \35092 );
not \U$34751 ( \35094 , \35093 );
and \U$34752 ( \35095 , \35086 , \35094 );
and \U$34753 ( \35096 , \35093 , \35085 );
and \U$34754 ( \35097 , \2042 , RI986df18_6);
and \U$34755 ( \35098 , RI986de28_4, \2040 );
nor \U$34756 ( \35099 , \35097 , \35098 );
not \U$34757 ( \35100 , \35099 );
not \U$34758 ( \35101 , \1462 );
and \U$34759 ( \35102 , \35100 , \35101 );
and \U$34760 ( \35103 , \35099 , \2034 );
nor \U$34761 ( \35104 , \35102 , \35103 );
nor \U$34762 ( \35105 , \35096 , \35104 );
nor \U$34763 ( \35106 , \35095 , \35105 );
xor \U$34764 ( \35107 , \35078 , \35106 );
and \U$34765 ( \35108 , \1293 , RI986f958_62);
and \U$34766 ( \35109 , RI986f4a8_52, \1291 );
nor \U$34767 ( \35110 , \35108 , \35109 );
not \U$34768 ( \35111 , \35110 );
not \U$34769 ( \35112 , \1128 );
and \U$34770 ( \35113 , \35111 , \35112 );
and \U$34771 ( \35114 , \35110 , \1128 );
nor \U$34772 ( \35115 , \35113 , \35114 );
and \U$34773 ( \35116 , \776 , RI986f778_58);
and \U$34774 ( \35117 , RI986fa48_64, \774 );
nor \U$34775 ( \35118 , \35116 , \35117 );
and \U$34776 ( \35119 , \35118 , \451 );
not \U$34777 ( \35120 , \35118 );
and \U$34778 ( \35121 , \35120 , \474 );
nor \U$34779 ( \35122 , \35119 , \35121 );
xor \U$34780 ( \35123 , \35115 , \35122 );
and \U$34781 ( \35124 , \438 , RI986e698_22);
and \U$34782 ( \35125 , RI986f868_60, \436 );
nor \U$34783 ( \35126 , \35124 , \35125 );
and \U$34784 ( \35127 , \35126 , \443 );
not \U$34785 ( \35128 , \35126 );
and \U$34786 ( \35129 , \35128 , \444 );
nor \U$34787 ( \35130 , \35127 , \35129 );
and \U$34788 ( \35131 , \35123 , \35130 );
and \U$34789 ( \35132 , \35115 , \35122 );
or \U$34790 ( \35133 , \35131 , \35132 );
and \U$34791 ( \35134 , \35107 , \35133 );
and \U$34792 ( \35135 , \35078 , \35106 );
nor \U$34793 ( \35136 , \35134 , \35135 );
xor \U$34794 ( \35137 , \35052 , \35136 );
not \U$34795 ( \35138 , \34917 );
not \U$34796 ( \35139 , \34897 );
or \U$34797 ( \35140 , \35138 , \35139 );
or \U$34798 ( \35141 , \34897 , \34917 );
nand \U$34799 ( \35142 , \35140 , \35141 );
not \U$34800 ( \35143 , \35142 );
not \U$34801 ( \35144 , \34905 );
and \U$34802 ( \35145 , \35143 , \35144 );
and \U$34803 ( \35146 , \35142 , \34905 );
nor \U$34804 ( \35147 , \35145 , \35146 );
xor \U$34805 ( \35148 , \34843 , \34850 );
xor \U$34806 ( \35149 , \35148 , \34858 );
or \U$34807 ( \35150 , \35147 , \35149 );
not \U$34808 ( \35151 , \35149 );
not \U$34809 ( \35152 , \35147 );
or \U$34810 ( \35153 , \35151 , \35152 );
not \U$34811 ( \35154 , \34813 );
xor \U$34812 ( \35155 , \34821 , \34832 );
not \U$34813 ( \35156 , \35155 );
or \U$34814 ( \35157 , \35154 , \35156 );
or \U$34815 ( \35158 , \35155 , \34813 );
nand \U$34816 ( \35159 , \35157 , \35158 );
nand \U$34817 ( \35160 , \35153 , \35159 );
nand \U$34818 ( \35161 , \35150 , \35160 );
and \U$34819 ( \35162 , \35137 , \35161 );
and \U$34820 ( \35163 , \35052 , \35136 );
or \U$34821 ( \35164 , \35162 , \35163 );
not \U$34822 ( \35165 , \35164 );
or \U$34823 ( \35166 , \34986 , \35165 );
or \U$34824 ( \35167 , \35164 , \34985 );
not \U$34825 ( \35168 , \34626 );
xor \U$34826 ( \35169 , \34642 , \34634 );
not \U$34827 ( \35170 , \35169 );
or \U$34828 ( \35171 , \35168 , \35170 );
or \U$34829 ( \35172 , \35169 , \34626 );
nand \U$34830 ( \35173 , \35171 , \35172 );
xor \U$34831 ( \35174 , \34886 , \34888 );
xor \U$34832 ( \35175 , \35174 , \34919 );
and \U$34833 ( \35176 , \35173 , \35175 );
xor \U$34834 ( \35177 , \34727 , \34735 );
xor \U$34835 ( \35178 , \35177 , \34744 );
xor \U$34836 ( \35179 , \34925 , \34930 );
xor \U$34837 ( \35180 , \35178 , \35179 );
xor \U$34838 ( \35181 , \34886 , \34888 );
xor \U$34839 ( \35182 , \35181 , \34919 );
and \U$34840 ( \35183 , \35180 , \35182 );
and \U$34841 ( \35184 , \35173 , \35180 );
or \U$34842 ( \35185 , \35176 , \35183 , \35184 );
nand \U$34843 ( \35186 , \35167 , \35185 );
nand \U$34844 ( \35187 , \35166 , \35186 );
not \U$34845 ( \35188 , \34771 );
xor \U$34846 ( \35189 , \34750 , \34702 );
not \U$34847 ( \35190 , \35189 );
or \U$34848 ( \35191 , \35188 , \35190 );
or \U$34849 ( \35192 , \35189 , \34771 );
nand \U$34850 ( \35193 , \35191 , \35192 );
xor \U$34851 ( \35194 , \35187 , \35193 );
not \U$34852 ( \35195 , \34961 );
xor \U$34853 ( \35196 , \34947 , \34957 );
not \U$34854 ( \35197 , \35196 );
and \U$34855 ( \35198 , \35195 , \35197 );
and \U$34856 ( \35199 , \34961 , \35196 );
nor \U$34857 ( \35200 , \35198 , \35199 );
not \U$34858 ( \35201 , \34700 );
not \U$34859 ( \35202 , \34670 );
or \U$34860 ( \35203 , \35201 , \35202 );
or \U$34861 ( \35204 , \34670 , \34700 );
nand \U$34862 ( \35205 , \35203 , \35204 );
not \U$34863 ( \35206 , \35205 );
not \U$34864 ( \35207 , \34644 );
and \U$34865 ( \35208 , \35206 , \35207 );
and \U$34866 ( \35209 , \35205 , \34644 );
nor \U$34867 ( \35210 , \35208 , \35209 );
or \U$34868 ( \35211 , \35200 , \35210 );
not \U$34869 ( \35212 , \35210 );
not \U$34870 ( \35213 , \35200 );
or \U$34871 ( \35214 , \35212 , \35213 );
xor \U$34872 ( \35215 , \34864 , \34922 );
xor \U$34873 ( \35216 , \35215 , \34935 );
nand \U$34874 ( \35217 , \35214 , \35216 );
nand \U$34875 ( \35218 , \35211 , \35217 );
and \U$34876 ( \35219 , \35194 , \35218 );
and \U$34877 ( \35220 , \35187 , \35193 );
or \U$34878 ( \35221 , \35219 , \35220 );
and \U$34879 ( \35222 , \34983 , \35221 );
not \U$34880 ( \35223 , \34983 );
not \U$34881 ( \35224 , \35221 );
and \U$34882 ( \35225 , \35223 , \35224 );
xor \U$34883 ( \35226 , \35187 , \35193 );
xor \U$34884 ( \35227 , \35226 , \35218 );
xor \U$34885 ( \35228 , \34938 , \34964 );
xor \U$34886 ( \35229 , \35228 , \34967 );
and \U$34887 ( \35230 , \35227 , \35229 );
not \U$34888 ( \35231 , \35227 );
not \U$34889 ( \35232 , \35229 );
and \U$34890 ( \35233 , \35231 , \35232 );
xnor \U$34891 ( \35234 , \35164 , \35185 );
not \U$34892 ( \35235 , \35234 );
not \U$34893 ( \35236 , \34985 );
and \U$34894 ( \35237 , \35235 , \35236 );
and \U$34895 ( \35238 , \35234 , \34985 );
nor \U$34896 ( \35239 , \35237 , \35238 );
not \U$34897 ( \35240 , \35050 );
not \U$34898 ( \35241 , \35016 );
or \U$34899 ( \35242 , \35240 , \35241 );
or \U$34900 ( \35243 , \35016 , \35050 );
nand \U$34901 ( \35244 , \35242 , \35243 );
not \U$34902 ( \35245 , \35244 );
not \U$34903 ( \35246 , \34996 );
and \U$34904 ( \35247 , \35245 , \35246 );
and \U$34905 ( \35248 , \35244 , \34996 );
nor \U$34906 ( \35249 , \35247 , \35248 );
xor \U$34907 ( \35250 , \34795 , \3406 );
xor \U$34908 ( \35251 , \35250 , \34803 );
xor \U$34909 ( \35252 , \35249 , \35251 );
not \U$34910 ( \35253 , \35147 );
not \U$34911 ( \35254 , \35159 );
or \U$34912 ( \35255 , \35253 , \35254 );
or \U$34913 ( \35256 , \35147 , \35159 );
nand \U$34914 ( \35257 , \35255 , \35256 );
not \U$34915 ( \35258 , \35257 );
not \U$34916 ( \35259 , \35149 );
and \U$34917 ( \35260 , \35258 , \35259 );
and \U$34918 ( \35261 , \35257 , \35149 );
nor \U$34919 ( \35262 , \35260 , \35261 );
and \U$34920 ( \35263 , \35252 , \35262 );
and \U$34921 ( \35264 , \35249 , \35251 );
or \U$34922 ( \35265 , \35263 , \35264 );
not \U$34923 ( \35266 , \35265 );
xor \U$34924 ( \35267 , \34806 , \34834 );
xor \U$34925 ( \35268 , \35267 , \34861 );
not \U$34926 ( \35269 , \35268 );
and \U$34927 ( \35270 , \35266 , \35269 );
and \U$34928 ( \35271 , \35265 , \35268 );
and \U$34929 ( \35272 , \1311 , RI986f598_54);
and \U$34930 ( \35273 , RI986f688_56, \1309 );
nor \U$34931 ( \35274 , \35272 , \35273 );
and \U$34932 ( \35275 , \35274 , \1315 );
not \U$34933 ( \35276 , \35274 );
and \U$34934 ( \35277 , \35276 , \1458 );
nor \U$34935 ( \35278 , \35275 , \35277 );
and \U$34936 ( \35279 , \2042 , RI986e008_8);
and \U$34937 ( \35280 , RI986df18_6, \2040 );
nor \U$34938 ( \35281 , \35279 , \35280 );
not \U$34939 ( \35282 , \35281 );
not \U$34940 ( \35283 , \2034 );
and \U$34941 ( \35284 , \35282 , \35283 );
and \U$34942 ( \35285 , \35281 , \1462 );
nor \U$34943 ( \35286 , \35284 , \35285 );
xor \U$34944 ( \35287 , \35278 , \35286 );
and \U$34945 ( \35288 , \2274 , RI986de28_4);
and \U$34946 ( \35289 , RI986dd38_2, \2272 );
nor \U$34947 ( \35290 , \35288 , \35289 );
and \U$34948 ( \35291 , \35290 , \2031 );
not \U$34949 ( \35292 , \35290 );
and \U$34950 ( \35293 , \35292 , \2030 );
nor \U$34951 ( \35294 , \35291 , \35293 );
and \U$34952 ( \35295 , \35287 , \35294 );
and \U$34953 ( \35296 , \35278 , \35286 );
or \U$34954 ( \35297 , \35295 , \35296 );
and \U$34955 ( \35298 , \3254 , RI986e2d8_14);
and \U$34956 ( \35299 , RI986e3c8_16, \3252 );
nor \U$34957 ( \35300 , \35298 , \35299 );
not \U$34958 ( \35301 , \35300 );
not \U$34959 ( \35302 , \2935 );
and \U$34960 ( \35303 , \35301 , \35302 );
and \U$34961 ( \35304 , \35300 , \3406 );
nor \U$34962 ( \35305 , \35303 , \35304 );
xor \U$34963 ( \35306 , \35305 , \3412 );
and \U$34964 ( \35307 , \2464 , RI986e1e8_12);
and \U$34965 ( \35308 , RI986e0f8_10, \2462 );
nor \U$34966 ( \35309 , \35307 , \35308 );
and \U$34967 ( \35310 , \35309 , \2263 );
not \U$34968 ( \35311 , \35309 );
and \U$34969 ( \35312 , \35311 , \2468 );
nor \U$34970 ( \35313 , \35310 , \35312 );
and \U$34971 ( \35314 , \35306 , \35313 );
and \U$34972 ( \35315 , \35305 , \3412 );
or \U$34973 ( \35316 , \35314 , \35315 );
xor \U$34974 ( \35317 , \35297 , \35316 );
and \U$34975 ( \35318 , \1293 , RI986fa48_64);
and \U$34976 ( \35319 , RI986f958_62, \1291 );
nor \U$34977 ( \35320 , \35318 , \35319 );
not \U$34978 ( \35321 , \35320 );
not \U$34979 ( \35322 , \1128 );
and \U$34980 ( \35323 , \35321 , \35322 );
and \U$34981 ( \35324 , \35320 , \1301 );
nor \U$34982 ( \35325 , \35323 , \35324 );
and \U$34983 ( \35326 , \776 , RI986f868_60);
and \U$34984 ( \35327 , RI986f778_58, \774 );
nor \U$34985 ( \35328 , \35326 , \35327 );
and \U$34986 ( \35329 , \35328 , \451 );
not \U$34987 ( \35330 , \35328 );
and \U$34988 ( \35331 , \35330 , \474 );
nor \U$34989 ( \35332 , \35329 , \35331 );
xor \U$34990 ( \35333 , \35325 , \35332 );
and \U$34991 ( \35334 , \1329 , RI986f4a8_52);
and \U$34992 ( \35335 , RI986f3b8_50, \1327 );
nor \U$34993 ( \35336 , \35334 , \35335 );
and \U$34994 ( \35337 , \35336 , \1337 );
not \U$34995 ( \35338 , \35336 );
and \U$34996 ( \35339 , \35338 , \1336 );
nor \U$34997 ( \35340 , \35337 , \35339 );
and \U$34998 ( \35341 , \35333 , \35340 );
and \U$34999 ( \35342 , \35325 , \35332 );
or \U$35000 ( \35343 , \35341 , \35342 );
and \U$35001 ( \35344 , \35317 , \35343 );
and \U$35002 ( \35345 , \35297 , \35316 );
or \U$35003 ( \35346 , \35344 , \35345 );
not \U$35004 ( \35347 , \456 );
and \U$35005 ( \35348 , \465 , RI986e5a8_20);
and \U$35006 ( \35349 , RI986e4b8_18, \463 );
nor \U$35007 ( \35350 , \35348 , \35349 );
not \U$35008 ( \35351 , \35350 );
or \U$35009 ( \35352 , \35347 , \35351 );
or \U$35010 ( \35353 , \35350 , \456 );
nand \U$35011 ( \35354 , \35352 , \35353 );
and \U$35012 ( \35355 , \438 , RI986e788_24);
and \U$35013 ( \35356 , RI986e698_22, \436 );
nor \U$35014 ( \35357 , \35355 , \35356 );
and \U$35015 ( \35358 , \35357 , \444 );
not \U$35016 ( \35359 , \35357 );
and \U$35017 ( \35360 , \35359 , \443 );
nor \U$35018 ( \35361 , \35358 , \35360 );
xor \U$35019 ( \35362 , \35354 , \35361 );
not \U$35020 ( \35363 , \367 );
and \U$35021 ( \35364 , \376 , RI986f2c8_48);
and \U$35022 ( \35365 , RI986f1d8_46, \374 );
nor \U$35023 ( \35366 , \35364 , \35365 );
not \U$35024 ( \35367 , \35366 );
or \U$35025 ( \35368 , \35363 , \35367 );
or \U$35026 ( \35369 , \35366 , \367 );
nand \U$35027 ( \35370 , \35368 , \35369 );
and \U$35028 ( \35371 , \35362 , \35370 );
and \U$35029 ( \35372 , \35354 , \35361 );
or \U$35030 ( \35373 , \35371 , \35372 );
not \U$35031 ( \35374 , \386 );
and \U$35032 ( \35375 , \395 , RI986f0e8_44);
and \U$35033 ( \35376 , RI986eff8_42, \393 );
nor \U$35034 ( \35377 , \35375 , \35376 );
not \U$35035 ( \35378 , \35377 );
or \U$35036 ( \35379 , \35374 , \35378 );
or \U$35037 ( \35380 , \35377 , \487 );
nand \U$35038 ( \35381 , \35379 , \35380 );
not \U$35039 ( \35382 , \345 );
and \U$35040 ( \35383 , \354 , RI986ec38_34);
and \U$35041 ( \35384 , RI986ed28_36, \352 );
nor \U$35042 ( \35385 , \35383 , \35384 );
not \U$35043 ( \35386 , \35385 );
or \U$35044 ( \35387 , \35382 , \35386 );
or \U$35045 ( \35388 , \35385 , \361 );
nand \U$35046 ( \35389 , \35387 , \35388 );
xor \U$35047 ( \35390 , \35381 , \35389 );
and \U$35048 ( \35391 , \416 , RI986ef08_40);
and \U$35049 ( \35392 , RI986ee18_38, \414 );
nor \U$35050 ( \35393 , \35391 , \35392 );
and \U$35051 ( \35394 , \35393 , \422 );
not \U$35052 ( \35395 , \35393 );
and \U$35053 ( \35396 , \35395 , \421 );
nor \U$35054 ( \35397 , \35394 , \35396 );
and \U$35055 ( \35398 , \35390 , \35397 );
and \U$35056 ( \35399 , \35381 , \35389 );
or \U$35057 ( \35400 , \35398 , \35399 );
nor \U$35058 ( \35401 , \35373 , \35400 );
xor \U$35059 ( \35402 , \35346 , \35401 );
not \U$35060 ( \35403 , \35028 );
not \U$35061 ( \35404 , \35048 );
or \U$35062 ( \35405 , \35403 , \35404 );
or \U$35063 ( \35406 , \35028 , \35048 );
nand \U$35064 ( \35407 , \35405 , \35406 );
not \U$35065 ( \35408 , \35407 );
not \U$35066 ( \35409 , \35036 );
and \U$35067 ( \35410 , \35408 , \35409 );
and \U$35068 ( \35411 , \35407 , \35036 );
nor \U$35069 ( \35412 , \35410 , \35411 );
xor \U$35070 ( \35413 , \35003 , \35004 );
xor \U$35071 ( \35414 , \35413 , \35013 );
and \U$35072 ( \35415 , \35412 , \35414 );
xor \U$35073 ( \35416 , \35115 , \35122 );
xor \U$35074 ( \35417 , \35416 , \35130 );
xor \U$35075 ( \35418 , \35003 , \35004 );
xor \U$35076 ( \35419 , \35418 , \35013 );
and \U$35077 ( \35420 , \35417 , \35419 );
and \U$35078 ( \35421 , \35412 , \35417 );
or \U$35079 ( \35422 , \35415 , \35420 , \35421 );
and \U$35080 ( \35423 , \35402 , \35422 );
and \U$35081 ( \35424 , \35346 , \35401 );
or \U$35082 ( \35425 , \35423 , \35424 );
nor \U$35083 ( \35426 , \35271 , \35425 );
nor \U$35084 ( \35427 , \35270 , \35426 );
xor \U$35085 ( \35428 , \35239 , \35427 );
not \U$35086 ( \35429 , \35210 );
not \U$35087 ( \35430 , \35216 );
or \U$35088 ( \35431 , \35429 , \35430 );
or \U$35089 ( \35432 , \35216 , \35210 );
nand \U$35090 ( \35433 , \35431 , \35432 );
not \U$35091 ( \35434 , \35433 );
not \U$35092 ( \35435 , \35200 );
and \U$35093 ( \35436 , \35434 , \35435 );
and \U$35094 ( \35437 , \35433 , \35200 );
nor \U$35095 ( \35438 , \35436 , \35437 );
and \U$35096 ( \35439 , \35428 , \35438 );
and \U$35097 ( \35440 , \35239 , \35427 );
or \U$35098 ( \35441 , \35439 , \35440 );
nor \U$35099 ( \35442 , \35233 , \35441 );
nor \U$35100 ( \35443 , \35230 , \35442 );
nor \U$35101 ( \35444 , \35225 , \35443 );
nor \U$35102 ( \35445 , \35222 , \35444 );
xor \U$35103 ( \35446 , \34599 , \34601 );
xor \U$35104 ( \35447 , \35446 , \34775 );
not \U$35105 ( \35448 , \35447 );
xor \U$35106 ( \35449 , \34970 , \34975 );
and \U$35107 ( \35450 , \35449 , \34982 );
and \U$35108 ( \35451 , \34970 , \34975 );
or \U$35109 ( \35452 , \35450 , \35451 );
not \U$35110 ( \35453 , \35452 );
and \U$35111 ( \35454 , \35448 , \35453 );
and \U$35112 ( \35455 , \35447 , \35452 );
nor \U$35113 ( \35456 , \35454 , \35455 );
not \U$35114 ( \35457 , \35456 );
xor \U$35115 ( \35458 , \34554 , \34571 );
xor \U$35116 ( \35459 , \35458 , \34576 );
not \U$35117 ( \35460 , \35459 );
and \U$35118 ( \35461 , \35457 , \35460 );
and \U$35119 ( \35462 , \35456 , \35459 );
nor \U$35120 ( \35463 , \35461 , \35462 );
or \U$35121 ( \35464 , \35445 , \35463 );
not \U$35122 ( \35465 , \34983 );
not \U$35123 ( \35466 , \35443 );
not \U$35124 ( \35467 , \35221 );
and \U$35125 ( \35468 , \35466 , \35467 );
and \U$35126 ( \35469 , \35443 , \35221 );
nor \U$35127 ( \35470 , \35468 , \35469 );
not \U$35128 ( \35471 , \35470 );
or \U$35129 ( \35472 , \35465 , \35471 );
or \U$35130 ( \35473 , \35470 , \34983 );
nand \U$35131 ( \35474 , \35472 , \35473 );
not \U$35132 ( \35475 , \35229 );
not \U$35133 ( \35476 , \35441 );
not \U$35134 ( \35477 , \35227 );
and \U$35135 ( \35478 , \35476 , \35477 );
and \U$35136 ( \35479 , \35441 , \35227 );
nor \U$35137 ( \35480 , \35478 , \35479 );
not \U$35138 ( \35481 , \35480 );
or \U$35139 ( \35482 , \35475 , \35481 );
or \U$35140 ( \35483 , \35480 , \35229 );
nand \U$35141 ( \35484 , \35482 , \35483 );
not \U$35142 ( \35485 , \35484 );
xor \U$35143 ( \35486 , \35239 , \35427 );
xor \U$35144 ( \35487 , \35486 , \35438 );
not \U$35145 ( \35488 , \35487 );
xor \U$35146 ( \35489 , \35052 , \35136 );
xor \U$35147 ( \35490 , \35489 , \35161 );
not \U$35148 ( \35491 , \35268 );
xor \U$35149 ( \35492 , \35425 , \35265 );
not \U$35150 ( \35493 , \35492 );
or \U$35151 ( \35494 , \35491 , \35493 );
or \U$35152 ( \35495 , \35492 , \35268 );
nand \U$35153 ( \35496 , \35494 , \35495 );
and \U$35154 ( \35497 , \35490 , \35496 );
and \U$35155 ( \35498 , \35488 , \35497 );
not \U$35156 ( \35499 , \35488 );
not \U$35157 ( \35500 , \35497 );
and \U$35158 ( \35501 , \35499 , \35500 );
xor \U$35159 ( \35502 , \35078 , \35106 );
xor \U$35160 ( \35503 , \35502 , \35133 );
xor \U$35161 ( \35504 , \35346 , \35401 );
xor \U$35162 ( \35505 , \35504 , \35422 );
xor \U$35163 ( \35506 , \35503 , \35505 );
xor \U$35164 ( \35507 , \35249 , \35251 );
xor \U$35165 ( \35508 , \35507 , \35262 );
and \U$35166 ( \35509 , \35506 , \35508 );
and \U$35167 ( \35510 , \35503 , \35505 );
nor \U$35168 ( \35511 , \35509 , \35510 );
xor \U$35169 ( \35512 , \34886 , \34888 );
xor \U$35170 ( \35513 , \35512 , \34919 );
xor \U$35171 ( \35514 , \35173 , \35180 );
xor \U$35172 ( \35515 , \35513 , \35514 );
and \U$35173 ( \35516 , \35511 , \35515 );
not \U$35174 ( \35517 , \35511 );
not \U$35175 ( \35518 , \35515 );
and \U$35176 ( \35519 , \35517 , \35518 );
and \U$35177 ( \35520 , \1311 , RI986f3b8_50);
and \U$35178 ( \35521 , RI986f598_54, \1309 );
nor \U$35179 ( \35522 , \35520 , \35521 );
and \U$35180 ( \35523 , \35522 , \1458 );
not \U$35181 ( \35524 , \35522 );
and \U$35182 ( \35525 , \35524 , \1315 );
nor \U$35183 ( \35526 , \35523 , \35525 );
not \U$35184 ( \35527 , \1462 );
and \U$35185 ( \35528 , \2042 , RI986f688_56);
and \U$35186 ( \35529 , RI986e008_8, \2040 );
nor \U$35187 ( \35530 , \35528 , \35529 );
not \U$35188 ( \35531 , \35530 );
or \U$35189 ( \35532 , \35527 , \35531 );
or \U$35190 ( \35533 , \35530 , \2034 );
nand \U$35191 ( \35534 , \35532 , \35533 );
xor \U$35192 ( \35535 , \35526 , \35534 );
and \U$35193 ( \35536 , \2274 , RI986df18_6);
and \U$35194 ( \35537 , RI986de28_4, \2272 );
nor \U$35195 ( \35538 , \35536 , \35537 );
and \U$35196 ( \35539 , \35538 , \2030 );
not \U$35197 ( \35540 , \35538 );
and \U$35198 ( \35541 , \35540 , \2031 );
nor \U$35199 ( \35542 , \35539 , \35541 );
and \U$35200 ( \35543 , \35535 , \35542 );
and \U$35201 ( \35544 , \35526 , \35534 );
or \U$35202 ( \35545 , \35543 , \35544 );
and \U$35203 ( \35546 , \2464 , RI986dd38_2);
and \U$35204 ( \35547 , RI986e1e8_12, \2462 );
nor \U$35205 ( \35548 , \35546 , \35547 );
and \U$35206 ( \35549 , \35548 , \2468 );
not \U$35207 ( \35550 , \35548 );
and \U$35208 ( \35551 , \35550 , \2263 );
nor \U$35209 ( \35552 , \35549 , \35551 );
not \U$35210 ( \35553 , \3918 );
nand \U$35211 ( \35554 , RI986e3c8_16, \3683 );
not \U$35212 ( \35555 , \35554 );
or \U$35213 ( \35556 , \35553 , \35555 );
or \U$35214 ( \35557 , \35554 , \3412 );
nand \U$35215 ( \35558 , \35556 , \35557 );
xor \U$35216 ( \35559 , \35552 , \35558 );
not \U$35217 ( \35560 , \3406 );
and \U$35218 ( \35561 , \3254 , RI986e0f8_10);
and \U$35219 ( \35562 , RI986e2d8_14, \3252 );
nor \U$35220 ( \35563 , \35561 , \35562 );
not \U$35221 ( \35564 , \35563 );
or \U$35222 ( \35565 , \35560 , \35564 );
or \U$35223 ( \35566 , \35563 , \2935 );
nand \U$35224 ( \35567 , \35565 , \35566 );
and \U$35225 ( \35568 , \35559 , \35567 );
and \U$35226 ( \35569 , \35552 , \35558 );
or \U$35227 ( \35570 , \35568 , \35569 );
xor \U$35228 ( \35571 , \35545 , \35570 );
and \U$35229 ( \35572 , \776 , RI986e698_22);
and \U$35230 ( \35573 , RI986f868_60, \774 );
nor \U$35231 ( \35574 , \35572 , \35573 );
and \U$35232 ( \35575 , \35574 , \474 );
not \U$35233 ( \35576 , \35574 );
and \U$35234 ( \35577 , \35576 , \451 );
nor \U$35235 ( \35578 , \35575 , \35577 );
not \U$35236 ( \35579 , \1301 );
and \U$35237 ( \35580 , \1293 , RI986f778_58);
and \U$35238 ( \35581 , RI986fa48_64, \1291 );
nor \U$35239 ( \35582 , \35580 , \35581 );
not \U$35240 ( \35583 , \35582 );
or \U$35241 ( \35584 , \35579 , \35583 );
or \U$35242 ( \35585 , \35582 , \1128 );
nand \U$35243 ( \35586 , \35584 , \35585 );
xor \U$35244 ( \35587 , \35578 , \35586 );
and \U$35245 ( \35588 , \1329 , RI986f958_62);
and \U$35246 ( \35589 , RI986f4a8_52, \1327 );
nor \U$35247 ( \35590 , \35588 , \35589 );
and \U$35248 ( \35591 , \35590 , \1336 );
not \U$35249 ( \35592 , \35590 );
and \U$35250 ( \35593 , \35592 , \1337 );
nor \U$35251 ( \35594 , \35591 , \35593 );
and \U$35252 ( \35595 , \35587 , \35594 );
and \U$35253 ( \35596 , \35578 , \35586 );
or \U$35254 ( \35597 , \35595 , \35596 );
and \U$35255 ( \35598 , \35571 , \35597 );
and \U$35256 ( \35599 , \35545 , \35570 );
or \U$35257 ( \35600 , \35598 , \35599 );
not \U$35258 ( \35601 , \361 );
and \U$35259 ( \35602 , \354 , RI986ee18_38);
and \U$35260 ( \35603 , RI986ec38_34, \352 );
nor \U$35261 ( \35604 , \35602 , \35603 );
not \U$35262 ( \35605 , \35604 );
or \U$35263 ( \35606 , \35601 , \35605 );
or \U$35264 ( \35607 , \35604 , \361 );
nand \U$35265 ( \35608 , \35606 , \35607 );
not \U$35266 ( \35609 , \386 );
and \U$35267 ( \35610 , \395 , RI986ed28_36);
and \U$35268 ( \35611 , RI986f0e8_44, \393 );
nor \U$35269 ( \35612 , \35610 , \35611 );
not \U$35270 ( \35613 , \35612 );
or \U$35271 ( \35614 , \35609 , \35613 );
or \U$35272 ( \35615 , \35612 , \386 );
nand \U$35273 ( \35616 , \35614 , \35615 );
xor \U$35274 ( \35617 , \35608 , \35616 );
and \U$35275 ( \35618 , \416 , RI986e878_26);
and \U$35276 ( \35619 , RI986ef08_40, \414 );
nor \U$35277 ( \35620 , \35618 , \35619 );
and \U$35278 ( \35621 , \35620 , \422 );
not \U$35279 ( \35622 , \35620 );
and \U$35280 ( \35623 , \35622 , \421 );
nor \U$35281 ( \35624 , \35621 , \35623 );
and \U$35282 ( \35625 , \35617 , \35624 );
and \U$35283 ( \35626 , \35608 , \35616 );
or \U$35284 ( \35627 , \35625 , \35626 );
nand \U$35285 ( \35628 , RI986e968_28, RI9871fc8_144);
not \U$35286 ( \35629 , \35628 );
xor \U$35287 ( \35630 , \35627 , \35629 );
not \U$35288 ( \35631 , \367 );
and \U$35289 ( \35632 , \376 , RI986eff8_42);
and \U$35290 ( \35633 , RI986f2c8_48, \374 );
nor \U$35291 ( \35634 , \35632 , \35633 );
not \U$35292 ( \35635 , \35634 );
or \U$35293 ( \35636 , \35631 , \35635 );
or \U$35294 ( \35637 , \35634 , \367 );
nand \U$35295 ( \35638 , \35636 , \35637 );
and \U$35296 ( \35639 , \438 , RI986e4b8_18);
and \U$35297 ( \35640 , RI986e788_24, \436 );
nor \U$35298 ( \35641 , \35639 , \35640 );
and \U$35299 ( \35642 , \35641 , \444 );
not \U$35300 ( \35643 , \35641 );
and \U$35301 ( \35644 , \35643 , \443 );
nor \U$35302 ( \35645 , \35642 , \35644 );
xor \U$35303 ( \35646 , \35638 , \35645 );
not \U$35304 ( \35647 , \456 );
and \U$35305 ( \35648 , \465 , RI986f1d8_46);
and \U$35306 ( \35649 , RI986e5a8_20, \463 );
nor \U$35307 ( \35650 , \35648 , \35649 );
not \U$35308 ( \35651 , \35650 );
or \U$35309 ( \35652 , \35647 , \35651 );
or \U$35310 ( \35653 , \35650 , \456 );
nand \U$35311 ( \35654 , \35652 , \35653 );
and \U$35312 ( \35655 , \35646 , \35654 );
and \U$35313 ( \35656 , \35638 , \35645 );
or \U$35314 ( \35657 , \35655 , \35656 );
and \U$35315 ( \35658 , \35630 , \35657 );
and \U$35316 ( \35659 , \35627 , \35629 );
or \U$35317 ( \35660 , \35658 , \35659 );
and \U$35318 ( \35661 , \35600 , \35660 );
not \U$35319 ( \35662 , \35600 );
not \U$35320 ( \35663 , \35660 );
and \U$35321 ( \35664 , \35662 , \35663 );
not \U$35322 ( \35665 , RI986e878_26);
nor \U$35323 ( \35666 , \35665 , \407 );
xor \U$35324 ( \35667 , \35381 , \35389 );
xor \U$35325 ( \35668 , \35667 , \35397 );
and \U$35326 ( \35669 , \35666 , \35668 );
xor \U$35327 ( \35670 , \35354 , \35361 );
xor \U$35328 ( \35671 , \35670 , \35370 );
xor \U$35329 ( \35672 , \35381 , \35389 );
xor \U$35330 ( \35673 , \35672 , \35397 );
and \U$35331 ( \35674 , \35671 , \35673 );
and \U$35332 ( \35675 , \35666 , \35671 );
or \U$35333 ( \35676 , \35669 , \35674 , \35675 );
not \U$35334 ( \35677 , \35676 );
nor \U$35335 ( \35678 , \35664 , \35677 );
nor \U$35336 ( \35679 , \35661 , \35678 );
not \U$35337 ( \35680 , \35059 );
xor \U$35338 ( \35681 , \35076 , \35067 );
not \U$35339 ( \35682 , \35681 );
or \U$35340 ( \35683 , \35680 , \35682 );
or \U$35341 ( \35684 , \35681 , \35059 );
nand \U$35342 ( \35685 , \35683 , \35684 );
not \U$35343 ( \35686 , \35085 );
xor \U$35344 ( \35687 , \35093 , \35104 );
not \U$35345 ( \35688 , \35687 );
or \U$35346 ( \35689 , \35686 , \35688 );
or \U$35347 ( \35690 , \35687 , \35085 );
nand \U$35348 ( \35691 , \35689 , \35690 );
and \U$35349 ( \35692 , \35685 , \35691 );
not \U$35350 ( \35693 , \35685 );
not \U$35351 ( \35694 , \35691 );
and \U$35352 ( \35695 , \35693 , \35694 );
xor \U$35353 ( \35696 , \35305 , \3412 );
xor \U$35354 ( \35697 , \35696 , \35313 );
not \U$35355 ( \35698 , \35697 );
xor \U$35356 ( \35699 , \35325 , \35332 );
xor \U$35357 ( \35700 , \35699 , \35340 );
not \U$35358 ( \35701 , \35700 );
and \U$35359 ( \35702 , \35698 , \35701 );
and \U$35360 ( \35703 , \35697 , \35700 );
xor \U$35361 ( \35704 , \35278 , \35286 );
xor \U$35362 ( \35705 , \35704 , \35294 );
nor \U$35363 ( \35706 , \35703 , \35705 );
nor \U$35364 ( \35707 , \35702 , \35706 );
nor \U$35365 ( \35708 , \35695 , \35707 );
nor \U$35366 ( \35709 , \35692 , \35708 );
xor \U$35367 ( \35710 , \35679 , \35709 );
and \U$35368 ( \35711 , \35373 , \35400 );
nor \U$35369 ( \35712 , \35711 , \35401 );
xor \U$35370 ( \35713 , \35297 , \35316 );
xor \U$35371 ( \35714 , \35713 , \35343 );
and \U$35372 ( \35715 , \35712 , \35714 );
xor \U$35373 ( \35716 , \35003 , \35004 );
xor \U$35374 ( \35717 , \35716 , \35013 );
xor \U$35375 ( \35718 , \35412 , \35417 );
xor \U$35376 ( \35719 , \35717 , \35718 );
xor \U$35377 ( \35720 , \35297 , \35316 );
xor \U$35378 ( \35721 , \35720 , \35343 );
and \U$35379 ( \35722 , \35719 , \35721 );
and \U$35380 ( \35723 , \35712 , \35719 );
or \U$35381 ( \35724 , \35715 , \35722 , \35723 );
and \U$35382 ( \35725 , \35710 , \35724 );
and \U$35383 ( \35726 , \35679 , \35709 );
or \U$35384 ( \35727 , \35725 , \35726 );
nor \U$35385 ( \35728 , \35519 , \35727 );
nor \U$35386 ( \35729 , \35516 , \35728 );
nor \U$35387 ( \35730 , \35501 , \35729 );
nor \U$35388 ( \35731 , \35498 , \35730 );
nor \U$35389 ( \35732 , \35485 , \35731 );
and \U$35390 ( \35733 , \35474 , \35732 );
xor \U$35391 ( \35734 , \35732 , \35474 );
not \U$35392 ( \35735 , \1128 );
and \U$35393 ( \35736 , \1293 , RI986f868_60);
and \U$35394 ( \35737 , RI986f778_58, \1291 );
nor \U$35395 ( \35738 , \35736 , \35737 );
not \U$35396 ( \35739 , \35738 );
or \U$35397 ( \35740 , \35735 , \35739 );
or \U$35398 ( \35741 , \35738 , \1128 );
nand \U$35399 ( \35742 , \35740 , \35741 );
and \U$35400 ( \35743 , \1329 , RI986fa48_64);
and \U$35401 ( \35744 , RI986f958_62, \1327 );
nor \U$35402 ( \35745 , \35743 , \35744 );
and \U$35403 ( \35746 , \35745 , \1336 );
not \U$35404 ( \35747 , \35745 );
and \U$35405 ( \35748 , \35747 , \1337 );
nor \U$35406 ( \35749 , \35746 , \35748 );
xor \U$35407 ( \35750 , \35742 , \35749 );
and \U$35408 ( \35751 , \1311 , RI986f4a8_52);
and \U$35409 ( \35752 , RI986f3b8_50, \1309 );
nor \U$35410 ( \35753 , \35751 , \35752 );
and \U$35411 ( \35754 , \35753 , \1458 );
not \U$35412 ( \35755 , \35753 );
and \U$35413 ( \35756 , \35755 , \1315 );
nor \U$35414 ( \35757 , \35754 , \35756 );
and \U$35415 ( \35758 , \35750 , \35757 );
and \U$35416 ( \35759 , \35742 , \35749 );
or \U$35417 ( \35760 , \35758 , \35759 );
and \U$35418 ( \35761 , \3683 , RI986e2d8_14);
and \U$35419 ( \35762 , RI986e3c8_16, \3681 );
nor \U$35420 ( \35763 , \35761 , \35762 );
not \U$35421 ( \35764 , \35763 );
not \U$35422 ( \35765 , \3412 );
and \U$35423 ( \35766 , \35764 , \35765 );
and \U$35424 ( \35767 , \35763 , \3918 );
nor \U$35425 ( \35768 , \35766 , \35767 );
or \U$35426 ( \35769 , \35768 , \3923 );
and \U$35427 ( \35770 , \35768 , \3923 );
and \U$35428 ( \35771 , \3254 , RI986e1e8_12);
and \U$35429 ( \35772 , RI986e0f8_10, \3252 );
nor \U$35430 ( \35773 , \35771 , \35772 );
not \U$35431 ( \35774 , \35773 );
not \U$35432 ( \35775 , \2935 );
and \U$35433 ( \35776 , \35774 , \35775 );
and \U$35434 ( \35777 , \35773 , \3406 );
nor \U$35435 ( \35778 , \35776 , \35777 );
nor \U$35436 ( \35779 , \35770 , \35778 );
not \U$35437 ( \35780 , \35779 );
nand \U$35438 ( \35781 , \35769 , \35780 );
xor \U$35439 ( \35782 , \35760 , \35781 );
and \U$35440 ( \35783 , \2042 , RI986f598_54);
and \U$35441 ( \35784 , RI986f688_56, \2040 );
nor \U$35442 ( \35785 , \35783 , \35784 );
not \U$35443 ( \35786 , \35785 );
not \U$35444 ( \35787 , \1462 );
and \U$35445 ( \35788 , \35786 , \35787 );
and \U$35446 ( \35789 , \35785 , \1462 );
nor \U$35447 ( \35790 , \35788 , \35789 );
and \U$35448 ( \35791 , \2274 , RI986e008_8);
and \U$35449 ( \35792 , RI986df18_6, \2272 );
nor \U$35450 ( \35793 , \35791 , \35792 );
and \U$35451 ( \35794 , \35793 , \2031 );
not \U$35452 ( \35795 , \35793 );
and \U$35453 ( \35796 , \35795 , \2030 );
nor \U$35454 ( \35797 , \35794 , \35796 );
or \U$35455 ( \35798 , \35790 , \35797 );
not \U$35456 ( \35799 , \35797 );
not \U$35457 ( \35800 , \35790 );
or \U$35458 ( \35801 , \35799 , \35800 );
and \U$35459 ( \35802 , \2464 , RI986de28_4);
and \U$35460 ( \35803 , RI986dd38_2, \2462 );
nor \U$35461 ( \35804 , \35802 , \35803 );
and \U$35462 ( \35805 , \35804 , \2468 );
not \U$35463 ( \35806 , \35804 );
and \U$35464 ( \35807 , \35806 , \2263 );
nor \U$35465 ( \35808 , \35805 , \35807 );
nand \U$35466 ( \35809 , \35801 , \35808 );
nand \U$35467 ( \35810 , \35798 , \35809 );
and \U$35468 ( \35811 , \35782 , \35810 );
and \U$35469 ( \35812 , \35760 , \35781 );
or \U$35470 ( \35813 , \35811 , \35812 );
not \U$35471 ( \35814 , \365 );
and \U$35472 ( \35815 , \376 , RI986f0e8_44);
and \U$35473 ( \35816 , RI986eff8_42, \374 );
nor \U$35474 ( \35817 , \35815 , \35816 );
not \U$35475 ( \35818 , \35817 );
or \U$35476 ( \35819 , \35814 , \35818 );
or \U$35477 ( \35820 , \35817 , \367 );
nand \U$35478 ( \35821 , \35819 , \35820 );
not \U$35479 ( \35822 , \487 );
and \U$35480 ( \35823 , \395 , RI986ec38_34);
and \U$35481 ( \35824 , RI986ed28_36, \393 );
nor \U$35482 ( \35825 , \35823 , \35824 );
not \U$35483 ( \35826 , \35825 );
or \U$35484 ( \35827 , \35822 , \35826 );
or \U$35485 ( \35828 , \35825 , \386 );
nand \U$35486 ( \35829 , \35827 , \35828 );
xor \U$35487 ( \35830 , \35821 , \35829 );
not \U$35488 ( \35831 , \345 );
and \U$35489 ( \35832 , \354 , RI986ef08_40);
and \U$35490 ( \35833 , RI986ee18_38, \352 );
nor \U$35491 ( \35834 , \35832 , \35833 );
not \U$35492 ( \35835 , \35834 );
or \U$35493 ( \35836 , \35831 , \35835 );
or \U$35494 ( \35837 , \35834 , \361 );
nand \U$35495 ( \35838 , \35836 , \35837 );
and \U$35496 ( \35839 , \35830 , \35838 );
and \U$35497 ( \35840 , \35821 , \35829 );
or \U$35498 ( \35841 , \35839 , \35840 );
not \U$35499 ( \35842 , RI986ea58_30);
nor \U$35500 ( \35843 , \35842 , \407 );
and \U$35501 ( \35844 , \416 , RI986e968_28);
and \U$35502 ( \35845 , RI986e878_26, \414 );
nor \U$35503 ( \35846 , \35844 , \35845 );
and \U$35504 ( \35847 , \35846 , \422 );
not \U$35505 ( \35848 , \35846 );
and \U$35506 ( \35849 , \35848 , \421 );
nor \U$35507 ( \35850 , \35847 , \35849 );
and \U$35508 ( \35851 , \35843 , \35850 );
xor \U$35509 ( \35852 , \35841 , \35851 );
not \U$35510 ( \35853 , \454 );
and \U$35511 ( \35854 , \465 , RI986f2c8_48);
and \U$35512 ( \35855 , RI986f1d8_46, \463 );
nor \U$35513 ( \35856 , \35854 , \35855 );
not \U$35514 ( \35857 , \35856 );
or \U$35515 ( \35858 , \35853 , \35857 );
or \U$35516 ( \35859 , \35856 , \456 );
nand \U$35517 ( \35860 , \35858 , \35859 );
and \U$35518 ( \35861 , \776 , RI986e788_24);
and \U$35519 ( \35862 , RI986e698_22, \774 );
nor \U$35520 ( \35863 , \35861 , \35862 );
and \U$35521 ( \35864 , \35863 , \474 );
not \U$35522 ( \35865 , \35863 );
and \U$35523 ( \35866 , \35865 , \451 );
nor \U$35524 ( \35867 , \35864 , \35866 );
xor \U$35525 ( \35868 , \35860 , \35867 );
and \U$35526 ( \35869 , \438 , RI986e5a8_20);
and \U$35527 ( \35870 , RI986e4b8_18, \436 );
nor \U$35528 ( \35871 , \35869 , \35870 );
and \U$35529 ( \35872 , \35871 , \444 );
not \U$35530 ( \35873 , \35871 );
and \U$35531 ( \35874 , \35873 , \443 );
nor \U$35532 ( \35875 , \35872 , \35874 );
and \U$35533 ( \35876 , \35868 , \35875 );
and \U$35534 ( \35877 , \35860 , \35867 );
or \U$35535 ( \35878 , \35876 , \35877 );
and \U$35536 ( \35879 , \35852 , \35878 );
and \U$35537 ( \35880 , \35841 , \35851 );
or \U$35538 ( \35881 , \35879 , \35880 );
xor \U$35539 ( \35882 , \35813 , \35881 );
xor \U$35540 ( \35883 , \35638 , \35645 );
xor \U$35541 ( \35884 , \35883 , \35654 );
xor \U$35542 ( \35885 , \35884 , \35628 );
xor \U$35543 ( \35886 , \35608 , \35616 );
xor \U$35544 ( \35887 , \35886 , \35624 );
and \U$35545 ( \35888 , \35885 , \35887 );
and \U$35546 ( \35889 , \35884 , \35628 );
or \U$35547 ( \35890 , \35888 , \35889 );
and \U$35548 ( \35891 , \35882 , \35890 );
and \U$35549 ( \35892 , \35813 , \35881 );
or \U$35550 ( \35893 , \35891 , \35892 );
xor \U$35551 ( \35894 , \35545 , \35570 );
xor \U$35552 ( \35895 , \35894 , \35597 );
xor \U$35553 ( \35896 , \35627 , \35629 );
xor \U$35554 ( \35897 , \35896 , \35657 );
and \U$35555 ( \35898 , \35895 , \35897 );
xor \U$35556 ( \35899 , \35893 , \35898 );
xor \U$35557 ( \35900 , \35381 , \35389 );
xor \U$35558 ( \35901 , \35900 , \35397 );
xor \U$35559 ( \35902 , \35666 , \35671 );
xor \U$35560 ( \35903 , \35901 , \35902 );
xor \U$35561 ( \35904 , \35552 , \35558 );
xor \U$35562 ( \35905 , \35904 , \35567 );
xor \U$35563 ( \35906 , \35526 , \35534 );
xor \U$35564 ( \35907 , \35906 , \35542 );
and \U$35565 ( \35908 , \35905 , \35907 );
xor \U$35566 ( \35909 , \35578 , \35586 );
xor \U$35567 ( \35910 , \35909 , \35594 );
xor \U$35568 ( \35911 , \35526 , \35534 );
xor \U$35569 ( \35912 , \35911 , \35542 );
and \U$35570 ( \35913 , \35910 , \35912 );
and \U$35571 ( \35914 , \35905 , \35910 );
or \U$35572 ( \35915 , \35908 , \35913 , \35914 );
xor \U$35573 ( \35916 , \35903 , \35915 );
not \U$35574 ( \35917 , \35700 );
xor \U$35575 ( \35918 , \35705 , \35697 );
not \U$35576 ( \35919 , \35918 );
or \U$35577 ( \35920 , \35917 , \35919 );
or \U$35578 ( \35921 , \35918 , \35700 );
nand \U$35579 ( \35922 , \35920 , \35921 );
and \U$35580 ( \35923 , \35916 , \35922 );
and \U$35581 ( \35924 , \35903 , \35915 );
or \U$35582 ( \35925 , \35923 , \35924 );
and \U$35583 ( \35926 , \35899 , \35925 );
and \U$35584 ( \35927 , \35893 , \35898 );
or \U$35585 ( \35928 , \35926 , \35927 );
not \U$35586 ( \35929 , \35928 );
not \U$35587 ( \35930 , \35685 );
not \U$35588 ( \35931 , \35707 );
or \U$35589 ( \35932 , \35930 , \35931 );
or \U$35590 ( \35933 , \35707 , \35685 );
nand \U$35591 ( \35934 , \35932 , \35933 );
xor \U$35592 ( \35935 , \35691 , \35934 );
not \U$35593 ( \35936 , \35677 );
xor \U$35594 ( \35937 , \35600 , \35660 );
not \U$35595 ( \35938 , \35937 );
or \U$35596 ( \35939 , \35936 , \35938 );
or \U$35597 ( \35940 , \35937 , \35677 );
nand \U$35598 ( \35941 , \35939 , \35940 );
and \U$35599 ( \35942 , \35935 , \35941 );
not \U$35600 ( \35943 , \35935 );
not \U$35601 ( \35944 , \35941 );
and \U$35602 ( \35945 , \35943 , \35944 );
xor \U$35603 ( \35946 , \35297 , \35316 );
xor \U$35604 ( \35947 , \35946 , \35343 );
xor \U$35605 ( \35948 , \35712 , \35719 );
xor \U$35606 ( \35949 , \35947 , \35948 );
nor \U$35607 ( \35950 , \35945 , \35949 );
nor \U$35608 ( \35951 , \35942 , \35950 );
not \U$35609 ( \35952 , \35951 );
or \U$35610 ( \35953 , \35929 , \35952 );
or \U$35611 ( \35954 , \35951 , \35928 );
nand \U$35612 ( \35955 , \35953 , \35954 );
not \U$35613 ( \35956 , \35955 );
xor \U$35614 ( \35957 , \35503 , \35505 );
xor \U$35615 ( \35958 , \35957 , \35508 );
not \U$35616 ( \35959 , \35958 );
and \U$35617 ( \35960 , \35956 , \35959 );
and \U$35618 ( \35961 , \35955 , \35958 );
nor \U$35619 ( \35962 , \35960 , \35961 );
xor \U$35620 ( \35963 , \35679 , \35709 );
xor \U$35621 ( \35964 , \35963 , \35724 );
or \U$35622 ( \35965 , \35962 , \35964 );
not \U$35623 ( \35966 , \35964 );
not \U$35624 ( \35967 , \35962 );
or \U$35625 ( \35968 , \35966 , \35967 );
xor \U$35626 ( \35969 , \35895 , \35897 );
xor \U$35627 ( \35970 , \35813 , \35881 );
xor \U$35628 ( \35971 , \35970 , \35890 );
and \U$35629 ( \35972 , \35969 , \35971 );
xor \U$35630 ( \35973 , \35903 , \35915 );
xor \U$35631 ( \35974 , \35973 , \35922 );
xor \U$35632 ( \35975 , \35813 , \35881 );
xor \U$35633 ( \35976 , \35975 , \35890 );
and \U$35634 ( \35977 , \35974 , \35976 );
and \U$35635 ( \35978 , \35969 , \35974 );
or \U$35636 ( \35979 , \35972 , \35977 , \35978 );
and \U$35637 ( \35980 , \3254 , RI986dd38_2);
and \U$35638 ( \35981 , RI986e1e8_12, \3252 );
nor \U$35639 ( \35982 , \35980 , \35981 );
not \U$35640 ( \35983 , \35982 );
not \U$35641 ( \35984 , \3406 );
and \U$35642 ( \35985 , \35983 , \35984 );
and \U$35643 ( \35986 , \35982 , \2935 );
nor \U$35644 ( \35987 , \35985 , \35986 );
not \U$35645 ( \35988 , \35987 );
and \U$35646 ( \35989 , \3683 , RI986e0f8_10);
and \U$35647 ( \35990 , RI986e2d8_14, \3681 );
nor \U$35648 ( \35991 , \35989 , \35990 );
not \U$35649 ( \35992 , \35991 );
not \U$35650 ( \35993 , \3412 );
and \U$35651 ( \35994 , \35992 , \35993 );
and \U$35652 ( \35995 , \35991 , \3412 );
nor \U$35653 ( \35996 , \35994 , \35995 );
not \U$35654 ( \35997 , \35996 );
and \U$35655 ( \35998 , \35988 , \35997 );
and \U$35656 ( \35999 , \35996 , \35987 );
nand \U$35657 ( \36000 , RI986e3c8_16, \4203 );
and \U$35658 ( \36001 , \36000 , \3922 );
not \U$35659 ( \36002 , \36000 );
and \U$35660 ( \36003 , \36002 , \4207 );
nor \U$35661 ( \36004 , \36001 , \36003 );
nor \U$35662 ( \36005 , \35999 , \36004 );
nor \U$35663 ( \36006 , \35998 , \36005 );
and \U$35664 ( \36007 , \2274 , RI986f688_56);
and \U$35665 ( \36008 , RI986e008_8, \2272 );
nor \U$35666 ( \36009 , \36007 , \36008 );
and \U$35667 ( \36010 , \36009 , \2030 );
not \U$35668 ( \36011 , \36009 );
and \U$35669 ( \36012 , \36011 , \2031 );
nor \U$35670 ( \36013 , \36010 , \36012 );
and \U$35671 ( \36014 , \2464 , RI986df18_6);
and \U$35672 ( \36015 , RI986de28_4, \2462 );
nor \U$35673 ( \36016 , \36014 , \36015 );
and \U$35674 ( \36017 , \36016 , \2468 );
not \U$35675 ( \36018 , \36016 );
and \U$35676 ( \36019 , \36018 , \2263 );
nor \U$35677 ( \36020 , \36017 , \36019 );
xor \U$35678 ( \36021 , \36013 , \36020 );
not \U$35679 ( \36022 , \1462 );
and \U$35680 ( \36023 , \2042 , RI986f3b8_50);
and \U$35681 ( \36024 , RI986f598_54, \2040 );
nor \U$35682 ( \36025 , \36023 , \36024 );
not \U$35683 ( \36026 , \36025 );
or \U$35684 ( \36027 , \36022 , \36026 );
or \U$35685 ( \36028 , \36025 , \1462 );
nand \U$35686 ( \36029 , \36027 , \36028 );
and \U$35687 ( \36030 , \36021 , \36029 );
and \U$35688 ( \36031 , \36013 , \36020 );
nor \U$35689 ( \36032 , \36030 , \36031 );
or \U$35690 ( \36033 , \36006 , \36032 );
not \U$35691 ( \36034 , \36006 );
not \U$35692 ( \36035 , \36032 );
or \U$35693 ( \36036 , \36034 , \36035 );
and \U$35694 ( \36037 , \1329 , RI986f778_58);
and \U$35695 ( \36038 , RI986fa48_64, \1327 );
nor \U$35696 ( \36039 , \36037 , \36038 );
and \U$35697 ( \36040 , \36039 , \1336 );
not \U$35698 ( \36041 , \36039 );
and \U$35699 ( \36042 , \36041 , \1337 );
nor \U$35700 ( \36043 , \36040 , \36042 );
not \U$35701 ( \36044 , \1128 );
and \U$35702 ( \36045 , \1293 , RI986e698_22);
and \U$35703 ( \36046 , RI986f868_60, \1291 );
nor \U$35704 ( \36047 , \36045 , \36046 );
not \U$35705 ( \36048 , \36047 );
or \U$35706 ( \36049 , \36044 , \36048 );
or \U$35707 ( \36050 , \36047 , \1301 );
nand \U$35708 ( \36051 , \36049 , \36050 );
xor \U$35709 ( \36052 , \36043 , \36051 );
and \U$35710 ( \36053 , \1311 , RI986f958_62);
and \U$35711 ( \36054 , RI986f4a8_52, \1309 );
nor \U$35712 ( \36055 , \36053 , \36054 );
and \U$35713 ( \36056 , \36055 , \1458 );
not \U$35714 ( \36057 , \36055 );
and \U$35715 ( \36058 , \36057 , \1318 );
nor \U$35716 ( \36059 , \36056 , \36058 );
and \U$35717 ( \36060 , \36052 , \36059 );
and \U$35718 ( \36061 , \36043 , \36051 );
or \U$35719 ( \36062 , \36060 , \36061 );
nand \U$35720 ( \36063 , \36036 , \36062 );
nand \U$35721 ( \36064 , \36033 , \36063 );
not \U$35722 ( \36065 , \345 );
and \U$35723 ( \36066 , \354 , RI986e878_26);
and \U$35724 ( \36067 , RI986ef08_40, \352 );
nor \U$35725 ( \36068 , \36066 , \36067 );
not \U$35726 ( \36069 , \36068 );
or \U$35727 ( \36070 , \36065 , \36069 );
or \U$35728 ( \36071 , \36068 , \361 );
nand \U$35729 ( \36072 , \36070 , \36071 );
not \U$35730 ( \36073 , \367 );
and \U$35731 ( \36074 , \376 , RI986ed28_36);
and \U$35732 ( \36075 , RI986f0e8_44, \374 );
nor \U$35733 ( \36076 , \36074 , \36075 );
not \U$35734 ( \36077 , \36076 );
or \U$35735 ( \36078 , \36073 , \36077 );
or \U$35736 ( \36079 , \36076 , \367 );
nand \U$35737 ( \36080 , \36078 , \36079 );
xor \U$35738 ( \36081 , \36072 , \36080 );
not \U$35739 ( \36082 , \487 );
and \U$35740 ( \36083 , \395 , RI986ee18_38);
and \U$35741 ( \36084 , RI986ec38_34, \393 );
nor \U$35742 ( \36085 , \36083 , \36084 );
not \U$35743 ( \36086 , \36085 );
or \U$35744 ( \36087 , \36082 , \36086 );
or \U$35745 ( \36088 , \36085 , \487 );
nand \U$35746 ( \36089 , \36087 , \36088 );
and \U$35747 ( \36090 , \36081 , \36089 );
and \U$35748 ( \36091 , \36072 , \36080 );
or \U$35749 ( \36092 , \36090 , \36091 );
nand \U$35750 ( \36093 , RI986eb48_32, RI9871fc8_144);
and \U$35751 ( \36094 , \416 , RI986ea58_30);
and \U$35752 ( \36095 , RI986e968_28, \414 );
nor \U$35753 ( \36096 , \36094 , \36095 );
and \U$35754 ( \36097 , \36096 , \421 );
not \U$35755 ( \36098 , \36096 );
and \U$35756 ( \36099 , \36098 , \422 );
nor \U$35757 ( \36100 , \36097 , \36099 );
nand \U$35758 ( \36101 , \36093 , \36100 );
xor \U$35759 ( \36102 , \36092 , \36101 );
not \U$35760 ( \36103 , \454 );
and \U$35761 ( \36104 , \465 , RI986eff8_42);
and \U$35762 ( \36105 , RI986f2c8_48, \463 );
nor \U$35763 ( \36106 , \36104 , \36105 );
not \U$35764 ( \36107 , \36106 );
or \U$35765 ( \36108 , \36103 , \36107 );
or \U$35766 ( \36109 , \36106 , \456 );
nand \U$35767 ( \36110 , \36108 , \36109 );
and \U$35768 ( \36111 , \776 , RI986e4b8_18);
and \U$35769 ( \36112 , RI986e788_24, \774 );
nor \U$35770 ( \36113 , \36111 , \36112 );
and \U$35771 ( \36114 , \36113 , \474 );
not \U$35772 ( \36115 , \36113 );
and \U$35773 ( \36116 , \36115 , \451 );
nor \U$35774 ( \36117 , \36114 , \36116 );
xor \U$35775 ( \36118 , \36110 , \36117 );
and \U$35776 ( \36119 , \438 , RI986f1d8_46);
and \U$35777 ( \36120 , RI986e5a8_20, \436 );
nor \U$35778 ( \36121 , \36119 , \36120 );
and \U$35779 ( \36122 , \36121 , \444 );
not \U$35780 ( \36123 , \36121 );
and \U$35781 ( \36124 , \36123 , \443 );
nor \U$35782 ( \36125 , \36122 , \36124 );
and \U$35783 ( \36126 , \36118 , \36125 );
and \U$35784 ( \36127 , \36110 , \36117 );
or \U$35785 ( \36128 , \36126 , \36127 );
and \U$35786 ( \36129 , \36102 , \36128 );
and \U$35787 ( \36130 , \36092 , \36101 );
or \U$35788 ( \36131 , \36129 , \36130 );
xor \U$35789 ( \36132 , \36064 , \36131 );
xor \U$35790 ( \36133 , \35843 , \35850 );
not \U$35791 ( \36134 , \36133 );
xor \U$35792 ( \36135 , \35860 , \35867 );
xor \U$35793 ( \36136 , \36135 , \35875 );
not \U$35794 ( \36137 , \36136 );
or \U$35795 ( \36138 , \36134 , \36137 );
or \U$35796 ( \36139 , \36136 , \36133 );
xor \U$35797 ( \36140 , \35821 , \35829 );
xor \U$35798 ( \36141 , \36140 , \35838 );
nand \U$35799 ( \36142 , \36139 , \36141 );
nand \U$35800 ( \36143 , \36138 , \36142 );
and \U$35801 ( \36144 , \36132 , \36143 );
and \U$35802 ( \36145 , \36064 , \36131 );
or \U$35803 ( \36146 , \36144 , \36145 );
xor \U$35804 ( \36147 , \35760 , \35781 );
xor \U$35805 ( \36148 , \36147 , \35810 );
xor \U$35806 ( \36149 , \35841 , \35851 );
xor \U$35807 ( \36150 , \36149 , \35878 );
and \U$35808 ( \36151 , \36148 , \36150 );
xor \U$35809 ( \36152 , \36146 , \36151 );
and \U$35810 ( \36153 , \35768 , \3922 );
not \U$35811 ( \36154 , \35768 );
and \U$35812 ( \36155 , \36154 , \4207 );
nor \U$35813 ( \36156 , \36153 , \36155 );
not \U$35814 ( \36157 , \36156 );
not \U$35815 ( \36158 , \35778 );
and \U$35816 ( \36159 , \36157 , \36158 );
and \U$35817 ( \36160 , \36156 , \35778 );
nor \U$35818 ( \36161 , \36159 , \36160 );
not \U$35819 ( \36162 , \35797 );
not \U$35820 ( \36163 , \35808 );
or \U$35821 ( \36164 , \36162 , \36163 );
or \U$35822 ( \36165 , \35797 , \35808 );
nand \U$35823 ( \36166 , \36164 , \36165 );
not \U$35824 ( \36167 , \36166 );
not \U$35825 ( \36168 , \35790 );
and \U$35826 ( \36169 , \36167 , \36168 );
and \U$35827 ( \36170 , \36166 , \35790 );
nor \U$35828 ( \36171 , \36169 , \36170 );
or \U$35829 ( \36172 , \36161 , \36171 );
not \U$35830 ( \36173 , \36171 );
not \U$35831 ( \36174 , \36161 );
or \U$35832 ( \36175 , \36173 , \36174 );
xor \U$35833 ( \36176 , \35742 , \35749 );
xor \U$35834 ( \36177 , \36176 , \35757 );
nand \U$35835 ( \36178 , \36175 , \36177 );
nand \U$35836 ( \36179 , \36172 , \36178 );
xor \U$35837 ( \36180 , \35884 , \35628 );
xor \U$35838 ( \36181 , \36180 , \35887 );
and \U$35839 ( \36182 , \36179 , \36181 );
xor \U$35840 ( \36183 , \35526 , \35534 );
xor \U$35841 ( \36184 , \36183 , \35542 );
xor \U$35842 ( \36185 , \35905 , \35910 );
xor \U$35843 ( \36186 , \36184 , \36185 );
xor \U$35844 ( \36187 , \35884 , \35628 );
xor \U$35845 ( \36188 , \36187 , \35887 );
and \U$35846 ( \36189 , \36186 , \36188 );
and \U$35847 ( \36190 , \36179 , \36186 );
or \U$35848 ( \36191 , \36182 , \36189 , \36190 );
and \U$35849 ( \36192 , \36152 , \36191 );
and \U$35850 ( \36193 , \36146 , \36151 );
or \U$35851 ( \36194 , \36192 , \36193 );
xor \U$35852 ( \36195 , \35979 , \36194 );
not \U$35853 ( \36196 , \35949 );
xor \U$35854 ( \36197 , \35941 , \35935 );
not \U$35855 ( \36198 , \36197 );
or \U$35856 ( \36199 , \36196 , \36198 );
or \U$35857 ( \36200 , \36197 , \35949 );
nand \U$35858 ( \36201 , \36199 , \36200 );
and \U$35859 ( \36202 , \36195 , \36201 );
and \U$35860 ( \36203 , \35979 , \36194 );
or \U$35861 ( \36204 , \36202 , \36203 );
nand \U$35862 ( \36205 , \35968 , \36204 );
nand \U$35863 ( \36206 , \35965 , \36205 );
xor \U$35864 ( \36207 , \35490 , \35496 );
not \U$35865 ( \36208 , \35515 );
not \U$35866 ( \36209 , \35511 );
not \U$35867 ( \36210 , \35727 );
and \U$35868 ( \36211 , \36209 , \36210 );
and \U$35869 ( \36212 , \35511 , \35727 );
nor \U$35870 ( \36213 , \36211 , \36212 );
not \U$35871 ( \36214 , \36213 );
or \U$35872 ( \36215 , \36208 , \36214 );
or \U$35873 ( \36216 , \36213 , \35515 );
nand \U$35874 ( \36217 , \36215 , \36216 );
xor \U$35875 ( \36218 , \36207 , \36217 );
or \U$35876 ( \36219 , \35958 , \35951 );
not \U$35877 ( \36220 , \35951 );
not \U$35878 ( \36221 , \35958 );
or \U$35879 ( \36222 , \36220 , \36221 );
nand \U$35880 ( \36223 , \36222 , \35928 );
nand \U$35881 ( \36224 , \36219 , \36223 );
xor \U$35882 ( \36225 , \36218 , \36224 );
xor \U$35883 ( \36226 , \36206 , \36225 );
xor \U$35884 ( \36227 , \35893 , \35898 );
xor \U$35885 ( \36228 , \36227 , \35925 );
xor \U$35886 ( \36229 , \35979 , \36194 );
xor \U$35887 ( \36230 , \36229 , \36201 );
and \U$35888 ( \36231 , \36228 , \36230 );
xor \U$35889 ( \36232 , \36148 , \36150 );
xor \U$35890 ( \36233 , \36064 , \36131 );
xor \U$35891 ( \36234 , \36233 , \36143 );
and \U$35892 ( \36235 , \36232 , \36234 );
xor \U$35893 ( \36236 , \35884 , \35628 );
xor \U$35894 ( \36237 , \36236 , \35887 );
xor \U$35895 ( \36238 , \36179 , \36186 );
xor \U$35896 ( \36239 , \36237 , \36238 );
xor \U$35897 ( \36240 , \36064 , \36131 );
xor \U$35898 ( \36241 , \36240 , \36143 );
and \U$35899 ( \36242 , \36239 , \36241 );
and \U$35900 ( \36243 , \36232 , \36239 );
or \U$35901 ( \36244 , \36235 , \36242 , \36243 );
and \U$35902 ( \36245 , \1329 , RI986f868_60);
and \U$35903 ( \36246 , RI986f778_58, \1327 );
nor \U$35904 ( \36247 , \36245 , \36246 );
and \U$35905 ( \36248 , \36247 , \1337 );
not \U$35906 ( \36249 , \36247 );
and \U$35907 ( \36250 , \36249 , \1336 );
nor \U$35908 ( \36251 , \36248 , \36250 );
and \U$35909 ( \36252 , \1311 , RI986fa48_64);
and \U$35910 ( \36253 , RI986f958_62, \1309 );
nor \U$35911 ( \36254 , \36252 , \36253 );
and \U$35912 ( \36255 , \36254 , \1315 );
not \U$35913 ( \36256 , \36254 );
and \U$35914 ( \36257 , \36256 , \1458 );
nor \U$35915 ( \36258 , \36255 , \36257 );
or \U$35916 ( \36259 , \36251 , \36258 );
not \U$35917 ( \36260 , \36258 );
not \U$35918 ( \36261 , \36251 );
or \U$35919 ( \36262 , \36260 , \36261 );
not \U$35920 ( \36263 , \1462 );
and \U$35921 ( \36264 , \2042 , RI986f4a8_52);
and \U$35922 ( \36265 , RI986f3b8_50, \2040 );
nor \U$35923 ( \36266 , \36264 , \36265 );
not \U$35924 ( \36267 , \36266 );
or \U$35925 ( \36268 , \36263 , \36267 );
or \U$35926 ( \36269 , \36266 , \2034 );
nand \U$35927 ( \36270 , \36268 , \36269 );
nand \U$35928 ( \36271 , \36262 , \36270 );
nand \U$35929 ( \36272 , \36259 , \36271 );
and \U$35930 ( \36273 , \3683 , RI986e1e8_12);
and \U$35931 ( \36274 , RI986e0f8_10, \3681 );
nor \U$35932 ( \36275 , \36273 , \36274 );
not \U$35933 ( \36276 , \36275 );
not \U$35934 ( \36277 , \3918 );
and \U$35935 ( \36278 , \36276 , \36277 );
and \U$35936 ( \36279 , \36275 , \3918 );
nor \U$35937 ( \36280 , \36278 , \36279 );
or \U$35938 ( \36281 , \36280 , \4521 );
not \U$35939 ( \36282 , \4519 );
not \U$35940 ( \36283 , \36280 );
or \U$35941 ( \36284 , \36282 , \36283 );
and \U$35942 ( \36285 , \4203 , RI986e2d8_14);
and \U$35943 ( \36286 , RI986e3c8_16, \4201 );
nor \U$35944 ( \36287 , \36285 , \36286 );
and \U$35945 ( \36288 , \36287 , \4207 );
not \U$35946 ( \36289 , \36287 );
and \U$35947 ( \36290 , \36289 , \3923 );
nor \U$35948 ( \36291 , \36288 , \36290 );
nand \U$35949 ( \36292 , \36284 , \36291 );
nand \U$35950 ( \36293 , \36281 , \36292 );
xor \U$35951 ( \36294 , \36272 , \36293 );
and \U$35952 ( \36295 , \2274 , RI986f598_54);
and \U$35953 ( \36296 , RI986f688_56, \2272 );
nor \U$35954 ( \36297 , \36295 , \36296 );
and \U$35955 ( \36298 , \36297 , \2031 );
not \U$35956 ( \36299 , \36297 );
and \U$35957 ( \36300 , \36299 , \2030 );
nor \U$35958 ( \36301 , \36298 , \36300 );
and \U$35959 ( \36302 , \2464 , RI986e008_8);
and \U$35960 ( \36303 , RI986df18_6, \2462 );
nor \U$35961 ( \36304 , \36302 , \36303 );
and \U$35962 ( \36305 , \36304 , \2263 );
not \U$35963 ( \36306 , \36304 );
and \U$35964 ( \36307 , \36306 , \2468 );
nor \U$35965 ( \36308 , \36305 , \36307 );
or \U$35966 ( \36309 , \36301 , \36308 );
not \U$35967 ( \36310 , \36308 );
not \U$35968 ( \36311 , \36301 );
or \U$35969 ( \36312 , \36310 , \36311 );
not \U$35970 ( \36313 , \2935 );
and \U$35971 ( \36314 , \3254 , RI986de28_4);
and \U$35972 ( \36315 , RI986dd38_2, \3252 );
nor \U$35973 ( \36316 , \36314 , \36315 );
not \U$35974 ( \36317 , \36316 );
or \U$35975 ( \36318 , \36313 , \36317 );
or \U$35976 ( \36319 , \36316 , \3406 );
nand \U$35977 ( \36320 , \36318 , \36319 );
nand \U$35978 ( \36321 , \36312 , \36320 );
nand \U$35979 ( \36322 , \36309 , \36321 );
and \U$35980 ( \36323 , \36294 , \36322 );
and \U$35981 ( \36324 , \36272 , \36293 );
or \U$35982 ( \36325 , \36323 , \36324 );
and \U$35983 ( \36326 , \416 , RI986eb48_32);
and \U$35984 ( \36327 , RI986ea58_30, \414 );
nor \U$35985 ( \36328 , \36326 , \36327 );
and \U$35986 ( \36329 , \36328 , \421 );
not \U$35987 ( \36330 , \36328 );
and \U$35988 ( \36331 , \36330 , \422 );
nor \U$35989 ( \36332 , \36329 , \36331 );
nand \U$35990 ( \36333 , RI9871668_124, RI9871fc8_144);
xor \U$35991 ( \36334 , \36332 , \36333 );
and \U$35992 ( \36335 , \354 , RI986e968_28);
and \U$35993 ( \36336 , RI986e878_26, \352 );
nor \U$35994 ( \36337 , \36335 , \36336 );
not \U$35995 ( \36338 , \36337 );
not \U$35996 ( \36339 , \361 );
and \U$35997 ( \36340 , \36338 , \36339 );
and \U$35998 ( \36341 , \36337 , \361 );
nor \U$35999 ( \36342 , \36340 , \36341 );
and \U$36000 ( \36343 , \36334 , \36342 );
and \U$36001 ( \36344 , \36332 , \36333 );
or \U$36002 ( \36345 , \36343 , \36344 );
and \U$36003 ( \36346 , \376 , RI986ec38_34);
and \U$36004 ( \36347 , RI986ed28_36, \374 );
nor \U$36005 ( \36348 , \36346 , \36347 );
not \U$36006 ( \36349 , \36348 );
not \U$36007 ( \36350 , \367 );
and \U$36008 ( \36351 , \36349 , \36350 );
and \U$36009 ( \36352 , \36348 , \367 );
nor \U$36010 ( \36353 , \36351 , \36352 );
not \U$36011 ( \36354 , \36353 );
and \U$36012 ( \36355 , \395 , RI986ef08_40);
and \U$36013 ( \36356 , RI986ee18_38, \393 );
nor \U$36014 ( \36357 , \36355 , \36356 );
not \U$36015 ( \36358 , \36357 );
not \U$36016 ( \36359 , \386 );
and \U$36017 ( \36360 , \36358 , \36359 );
and \U$36018 ( \36361 , \36357 , \487 );
nor \U$36019 ( \36362 , \36360 , \36361 );
not \U$36020 ( \36363 , \36362 );
and \U$36021 ( \36364 , \36354 , \36363 );
and \U$36022 ( \36365 , \36362 , \36353 );
and \U$36023 ( \36366 , \465 , RI986f0e8_44);
and \U$36024 ( \36367 , RI986eff8_42, \463 );
nor \U$36025 ( \36368 , \36366 , \36367 );
not \U$36026 ( \36369 , \36368 );
not \U$36027 ( \36370 , \454 );
and \U$36028 ( \36371 , \36369 , \36370 );
and \U$36029 ( \36372 , \36368 , \454 );
nor \U$36030 ( \36373 , \36371 , \36372 );
nor \U$36031 ( \36374 , \36365 , \36373 );
nor \U$36032 ( \36375 , \36364 , \36374 );
xor \U$36033 ( \36376 , \36345 , \36375 );
and \U$36034 ( \36377 , \776 , RI986e5a8_20);
and \U$36035 ( \36378 , RI986e4b8_18, \774 );
nor \U$36036 ( \36379 , \36377 , \36378 );
and \U$36037 ( \36380 , \36379 , \474 );
not \U$36038 ( \36381 , \36379 );
and \U$36039 ( \36382 , \36381 , \451 );
nor \U$36040 ( \36383 , \36380 , \36382 );
not \U$36041 ( \36384 , \1301 );
and \U$36042 ( \36385 , \1293 , RI986e788_24);
and \U$36043 ( \36386 , RI986e698_22, \1291 );
nor \U$36044 ( \36387 , \36385 , \36386 );
not \U$36045 ( \36388 , \36387 );
or \U$36046 ( \36389 , \36384 , \36388 );
or \U$36047 ( \36390 , \36387 , \1128 );
nand \U$36048 ( \36391 , \36389 , \36390 );
xor \U$36049 ( \36392 , \36383 , \36391 );
and \U$36050 ( \36393 , \438 , RI986f2c8_48);
and \U$36051 ( \36394 , RI986f1d8_46, \436 );
nor \U$36052 ( \36395 , \36393 , \36394 );
and \U$36053 ( \36396 , \36395 , \444 );
not \U$36054 ( \36397 , \36395 );
and \U$36055 ( \36398 , \36397 , \443 );
nor \U$36056 ( \36399 , \36396 , \36398 );
and \U$36057 ( \36400 , \36392 , \36399 );
and \U$36058 ( \36401 , \36383 , \36391 );
nor \U$36059 ( \36402 , \36400 , \36401 );
and \U$36060 ( \36403 , \36376 , \36402 );
and \U$36061 ( \36404 , \36345 , \36375 );
nor \U$36062 ( \36405 , \36403 , \36404 );
xor \U$36063 ( \36406 , \36325 , \36405 );
or \U$36064 ( \36407 , \36100 , \36093 );
nand \U$36065 ( \36408 , \36407 , \36101 );
xor \U$36066 ( \36409 , \36110 , \36117 );
xor \U$36067 ( \36410 , \36409 , \36125 );
and \U$36068 ( \36411 , \36408 , \36410 );
xor \U$36069 ( \36412 , \36072 , \36080 );
xor \U$36070 ( \36413 , \36412 , \36089 );
xor \U$36071 ( \36414 , \36110 , \36117 );
xor \U$36072 ( \36415 , \36414 , \36125 );
and \U$36073 ( \36416 , \36413 , \36415 );
and \U$36074 ( \36417 , \36408 , \36413 );
or \U$36075 ( \36418 , \36411 , \36416 , \36417 );
and \U$36076 ( \36419 , \36406 , \36418 );
and \U$36077 ( \36420 , \36325 , \36405 );
nor \U$36078 ( \36421 , \36419 , \36420 );
not \U$36079 ( \36422 , \36062 );
not \U$36080 ( \36423 , \36006 );
or \U$36081 ( \36424 , \36422 , \36423 );
or \U$36082 ( \36425 , \36006 , \36062 );
nand \U$36083 ( \36426 , \36424 , \36425 );
not \U$36084 ( \36427 , \36426 );
not \U$36085 ( \36428 , \36032 );
and \U$36086 ( \36429 , \36427 , \36428 );
and \U$36087 ( \36430 , \36426 , \36032 );
nor \U$36088 ( \36431 , \36429 , \36430 );
not \U$36089 ( \36432 , \36431 );
xor \U$36090 ( \36433 , \36092 , \36101 );
xor \U$36091 ( \36434 , \36433 , \36128 );
nand \U$36092 ( \36435 , \36432 , \36434 );
or \U$36093 ( \36436 , \36421 , \36435 );
not \U$36094 ( \36437 , \36435 );
not \U$36095 ( \36438 , \36421 );
or \U$36096 ( \36439 , \36437 , \36438 );
xnor \U$36097 ( \36440 , \36141 , \36136 );
not \U$36098 ( \36441 , \36440 );
not \U$36099 ( \36442 , \36133 );
and \U$36100 ( \36443 , \36441 , \36442 );
and \U$36101 ( \36444 , \36440 , \36133 );
nor \U$36102 ( \36445 , \36443 , \36444 );
not \U$36103 ( \36446 , \36177 );
not \U$36104 ( \36447 , \36161 );
or \U$36105 ( \36448 , \36446 , \36447 );
or \U$36106 ( \36449 , \36161 , \36177 );
nand \U$36107 ( \36450 , \36448 , \36449 );
not \U$36108 ( \36451 , \36450 );
not \U$36109 ( \36452 , \36171 );
and \U$36110 ( \36453 , \36451 , \36452 );
and \U$36111 ( \36454 , \36450 , \36171 );
nor \U$36112 ( \36455 , \36453 , \36454 );
or \U$36113 ( \36456 , \36445 , \36455 );
not \U$36114 ( \36457 , \36445 );
not \U$36115 ( \36458 , \36455 );
or \U$36116 ( \36459 , \36457 , \36458 );
not \U$36117 ( \36460 , \35987 );
xor \U$36118 ( \36461 , \36004 , \35996 );
not \U$36119 ( \36462 , \36461 );
or \U$36120 ( \36463 , \36460 , \36462 );
or \U$36121 ( \36464 , \36461 , \35987 );
nand \U$36122 ( \36465 , \36463 , \36464 );
xor \U$36123 ( \36466 , \36043 , \36051 );
xor \U$36124 ( \36467 , \36466 , \36059 );
xor \U$36125 ( \36468 , \36465 , \36467 );
xor \U$36126 ( \36469 , \36013 , \36020 );
xor \U$36127 ( \36470 , \36469 , \36029 );
and \U$36128 ( \36471 , \36468 , \36470 );
and \U$36129 ( \36472 , \36465 , \36467 );
or \U$36130 ( \36473 , \36471 , \36472 );
nand \U$36131 ( \36474 , \36459 , \36473 );
nand \U$36132 ( \36475 , \36456 , \36474 );
nand \U$36133 ( \36476 , \36439 , \36475 );
nand \U$36134 ( \36477 , \36436 , \36476 );
xor \U$36135 ( \36478 , \36244 , \36477 );
xor \U$36136 ( \36479 , \35813 , \35881 );
xor \U$36137 ( \36480 , \36479 , \35890 );
xor \U$36138 ( \36481 , \35969 , \35974 );
xor \U$36139 ( \36482 , \36480 , \36481 );
and \U$36140 ( \36483 , \36478 , \36482 );
and \U$36141 ( \36484 , \36244 , \36477 );
or \U$36142 ( \36485 , \36483 , \36484 );
xor \U$36143 ( \36486 , \35979 , \36194 );
xor \U$36144 ( \36487 , \36486 , \36201 );
and \U$36145 ( \36488 , \36485 , \36487 );
and \U$36146 ( \36489 , \36228 , \36485 );
or \U$36147 ( \36490 , \36231 , \36488 , \36489 );
not \U$36148 ( \36491 , \36490 );
not \U$36149 ( \36492 , \35964 );
not \U$36150 ( \36493 , \36204 );
or \U$36151 ( \36494 , \36492 , \36493 );
or \U$36152 ( \36495 , \36204 , \35964 );
nand \U$36153 ( \36496 , \36494 , \36495 );
not \U$36154 ( \36497 , \36496 );
not \U$36155 ( \36498 , \35962 );
and \U$36156 ( \36499 , \36497 , \36498 );
and \U$36157 ( \36500 , \36496 , \35962 );
nor \U$36158 ( \36501 , \36499 , \36500 );
nor \U$36159 ( \36502 , \36491 , \36501 );
and \U$36160 ( \36503 , \36226 , \36502 );
xor \U$36161 ( \36504 , \36502 , \36226 );
not \U$36162 ( \36505 , \36501 );
not \U$36163 ( \36506 , \36490 );
and \U$36164 ( \36507 , \36505 , \36506 );
and \U$36165 ( \36508 , \36501 , \36490 );
nor \U$36166 ( \36509 , \36507 , \36508 );
xor \U$36167 ( \36510 , \36325 , \36405 );
xor \U$36168 ( \36511 , \36510 , \36418 );
not \U$36169 ( \36512 , \36431 );
not \U$36170 ( \36513 , \36434 );
or \U$36171 ( \36514 , \36512 , \36513 );
or \U$36172 ( \36515 , \36434 , \36431 );
nand \U$36173 ( \36516 , \36514 , \36515 );
and \U$36174 ( \36517 , \36511 , \36516 );
not \U$36175 ( \36518 , \36511 );
not \U$36176 ( \36519 , \36516 );
and \U$36177 ( \36520 , \36518 , \36519 );
not \U$36178 ( \36521 , \36473 );
not \U$36179 ( \36522 , \36455 );
or \U$36180 ( \36523 , \36521 , \36522 );
or \U$36181 ( \36524 , \36455 , \36473 );
nand \U$36182 ( \36525 , \36523 , \36524 );
not \U$36183 ( \36526 , \36525 );
not \U$36184 ( \36527 , \36445 );
and \U$36185 ( \36528 , \36526 , \36527 );
and \U$36186 ( \36529 , \36525 , \36445 );
nor \U$36187 ( \36530 , \36528 , \36529 );
nor \U$36188 ( \36531 , \36520 , \36530 );
nor \U$36189 ( \36532 , \36517 , \36531 );
and \U$36190 ( \36533 , \2274 , RI986f3b8_50);
and \U$36191 ( \36534 , RI986f598_54, \2272 );
nor \U$36192 ( \36535 , \36533 , \36534 );
and \U$36193 ( \36536 , \36535 , \2030 );
not \U$36194 ( \36537 , \36535 );
and \U$36195 ( \36538 , \36537 , \2031 );
nor \U$36196 ( \36539 , \36536 , \36538 );
and \U$36197 ( \36540 , \2464 , RI986f688_56);
and \U$36198 ( \36541 , RI986e008_8, \2462 );
nor \U$36199 ( \36542 , \36540 , \36541 );
and \U$36200 ( \36543 , \36542 , \2468 );
not \U$36201 ( \36544 , \36542 );
and \U$36202 ( \36545 , \36544 , \2263 );
nor \U$36203 ( \36546 , \36543 , \36545 );
xor \U$36204 ( \36547 , \36539 , \36546 );
not \U$36205 ( \36548 , \2935 );
and \U$36206 ( \36549 , \3254 , RI986df18_6);
and \U$36207 ( \36550 , RI986de28_4, \3252 );
nor \U$36208 ( \36551 , \36549 , \36550 );
not \U$36209 ( \36552 , \36551 );
or \U$36210 ( \36553 , \36548 , \36552 );
or \U$36211 ( \36554 , \36551 , \3406 );
nand \U$36212 ( \36555 , \36553 , \36554 );
and \U$36213 ( \36556 , \36547 , \36555 );
and \U$36214 ( \36557 , \36539 , \36546 );
or \U$36215 ( \36558 , \36556 , \36557 );
not \U$36216 ( \36559 , \3918 );
and \U$36217 ( \36560 , \3683 , RI986dd38_2);
and \U$36218 ( \36561 , RI986e1e8_12, \3681 );
nor \U$36219 ( \36562 , \36560 , \36561 );
not \U$36220 ( \36563 , \36562 );
or \U$36221 ( \36564 , \36559 , \36563 );
or \U$36222 ( \36565 , \36562 , \3412 );
nand \U$36223 ( \36566 , \36564 , \36565 );
not \U$36224 ( \36567 , \4519 );
nand \U$36225 ( \36568 , RI986e3c8_16, \4710 );
not \U$36226 ( \36569 , \36568 );
or \U$36227 ( \36570 , \36567 , \36569 );
or \U$36228 ( \36571 , \36568 , \4519 );
nand \U$36229 ( \36572 , \36570 , \36571 );
xor \U$36230 ( \36573 , \36566 , \36572 );
and \U$36231 ( \36574 , \4203 , RI986e0f8_10);
and \U$36232 ( \36575 , RI986e2d8_14, \4201 );
nor \U$36233 ( \36576 , \36574 , \36575 );
and \U$36234 ( \36577 , \36576 , \4207 );
not \U$36235 ( \36578 , \36576 );
and \U$36236 ( \36579 , \36578 , \3922 );
nor \U$36237 ( \36580 , \36577 , \36579 );
and \U$36238 ( \36581 , \36573 , \36580 );
and \U$36239 ( \36582 , \36566 , \36572 );
or \U$36240 ( \36583 , \36581 , \36582 );
xor \U$36241 ( \36584 , \36558 , \36583 );
and \U$36242 ( \36585 , \1329 , RI986e698_22);
and \U$36243 ( \36586 , RI986f868_60, \1327 );
nor \U$36244 ( \36587 , \36585 , \36586 );
and \U$36245 ( \36588 , \36587 , \1336 );
not \U$36246 ( \36589 , \36587 );
and \U$36247 ( \36590 , \36589 , \1337 );
nor \U$36248 ( \36591 , \36588 , \36590 );
and \U$36249 ( \36592 , \1311 , RI986f778_58);
and \U$36250 ( \36593 , RI986fa48_64, \1309 );
nor \U$36251 ( \36594 , \36592 , \36593 );
and \U$36252 ( \36595 , \36594 , \1319 );
not \U$36253 ( \36596 , \36594 );
and \U$36254 ( \36597 , \36596 , \1318 );
nor \U$36255 ( \36598 , \36595 , \36597 );
xor \U$36256 ( \36599 , \36591 , \36598 );
not \U$36257 ( \36600 , \2034 );
and \U$36258 ( \36601 , \2042 , RI986f958_62);
and \U$36259 ( \36602 , RI986f4a8_52, \2040 );
nor \U$36260 ( \36603 , \36601 , \36602 );
not \U$36261 ( \36604 , \36603 );
or \U$36262 ( \36605 , \36600 , \36604 );
or \U$36263 ( \36606 , \36603 , \1462 );
nand \U$36264 ( \36607 , \36605 , \36606 );
and \U$36265 ( \36608 , \36599 , \36607 );
and \U$36266 ( \36609 , \36591 , \36598 );
or \U$36267 ( \36610 , \36608 , \36609 );
and \U$36268 ( \36611 , \36584 , \36610 );
and \U$36269 ( \36612 , \36558 , \36583 );
or \U$36270 ( \36613 , \36611 , \36612 );
and \U$36271 ( \36614 , \376 , RI986ee18_38);
and \U$36272 ( \36615 , RI986ec38_34, \374 );
nor \U$36273 ( \36616 , \36614 , \36615 );
not \U$36274 ( \36617 , \36616 );
not \U$36275 ( \36618 , \367 );
and \U$36276 ( \36619 , \36617 , \36618 );
and \U$36277 ( \36620 , \36616 , \365 );
nor \U$36278 ( \36621 , \36619 , \36620 );
and \U$36279 ( \36622 , \395 , RI986e878_26);
and \U$36280 ( \36623 , RI986ef08_40, \393 );
nor \U$36281 ( \36624 , \36622 , \36623 );
not \U$36282 ( \36625 , \36624 );
not \U$36283 ( \36626 , \386 );
and \U$36284 ( \36627 , \36625 , \36626 );
and \U$36285 ( \36628 , \36624 , \487 );
nor \U$36286 ( \36629 , \36627 , \36628 );
or \U$36287 ( \36630 , \36621 , \36629 );
not \U$36288 ( \36631 , \36629 );
not \U$36289 ( \36632 , \36621 );
or \U$36290 ( \36633 , \36631 , \36632 );
not \U$36291 ( \36634 , \456 );
and \U$36292 ( \36635 , \465 , RI986ed28_36);
and \U$36293 ( \36636 , RI986f0e8_44, \463 );
nor \U$36294 ( \36637 , \36635 , \36636 );
not \U$36295 ( \36638 , \36637 );
or \U$36296 ( \36639 , \36634 , \36638 );
or \U$36297 ( \36640 , \36637 , \456 );
nand \U$36298 ( \36641 , \36639 , \36640 );
nand \U$36299 ( \36642 , \36633 , \36641 );
nand \U$36300 ( \36643 , \36630 , \36642 );
and \U$36301 ( \36644 , \354 , RI986ea58_30);
and \U$36302 ( \36645 , RI986e968_28, \352 );
nor \U$36303 ( \36646 , \36644 , \36645 );
not \U$36304 ( \36647 , \36646 );
not \U$36305 ( \36648 , \361 );
and \U$36306 ( \36649 , \36647 , \36648 );
and \U$36307 ( \36650 , \36646 , \345 );
nor \U$36308 ( \36651 , \36649 , \36650 );
nand \U$36309 ( \36652 , RI9871578_122, RI9871fc8_144);
or \U$36310 ( \36653 , \36651 , \36652 );
not \U$36311 ( \36654 , \36652 );
not \U$36312 ( \36655 , \36651 );
or \U$36313 ( \36656 , \36654 , \36655 );
and \U$36314 ( \36657 , \416 , RI9871668_124);
and \U$36315 ( \36658 , RI986eb48_32, \414 );
nor \U$36316 ( \36659 , \36657 , \36658 );
and \U$36317 ( \36660 , \36659 , \422 );
not \U$36318 ( \36661 , \36659 );
and \U$36319 ( \36662 , \36661 , \421 );
nor \U$36320 ( \36663 , \36660 , \36662 );
nand \U$36321 ( \36664 , \36656 , \36663 );
nand \U$36322 ( \36665 , \36653 , \36664 );
xor \U$36323 ( \36666 , \36643 , \36665 );
and \U$36324 ( \36667 , \438 , RI986eff8_42);
and \U$36325 ( \36668 , RI986f2c8_48, \436 );
nor \U$36326 ( \36669 , \36667 , \36668 );
and \U$36327 ( \36670 , \36669 , \444 );
not \U$36328 ( \36671 , \36669 );
and \U$36329 ( \36672 , \36671 , \443 );
nor \U$36330 ( \36673 , \36670 , \36672 );
and \U$36331 ( \36674 , \776 , RI986f1d8_46);
and \U$36332 ( \36675 , RI986e5a8_20, \774 );
nor \U$36333 ( \36676 , \36674 , \36675 );
and \U$36334 ( \36677 , \36676 , \474 );
not \U$36335 ( \36678 , \36676 );
and \U$36336 ( \36679 , \36678 , \451 );
nor \U$36337 ( \36680 , \36677 , \36679 );
xor \U$36338 ( \36681 , \36673 , \36680 );
not \U$36339 ( \36682 , \1301 );
and \U$36340 ( \36683 , \1293 , RI986e4b8_18);
and \U$36341 ( \36684 , RI986e788_24, \1291 );
nor \U$36342 ( \36685 , \36683 , \36684 );
not \U$36343 ( \36686 , \36685 );
or \U$36344 ( \36687 , \36682 , \36686 );
or \U$36345 ( \36688 , \36685 , \1301 );
nand \U$36346 ( \36689 , \36687 , \36688 );
and \U$36347 ( \36690 , \36681 , \36689 );
and \U$36348 ( \36691 , \36673 , \36680 );
or \U$36349 ( \36692 , \36690 , \36691 );
and \U$36350 ( \36693 , \36666 , \36692 );
and \U$36351 ( \36694 , \36643 , \36665 );
or \U$36352 ( \36695 , \36693 , \36694 );
and \U$36353 ( \36696 , \36613 , \36695 );
not \U$36354 ( \36697 , \36613 );
not \U$36355 ( \36698 , \36695 );
and \U$36356 ( \36699 , \36697 , \36698 );
xor \U$36357 ( \36700 , \36383 , \36391 );
xor \U$36358 ( \36701 , \36700 , \36399 );
not \U$36359 ( \36702 , \36362 );
xor \U$36360 ( \36703 , \36373 , \36353 );
not \U$36361 ( \36704 , \36703 );
or \U$36362 ( \36705 , \36702 , \36704 );
or \U$36363 ( \36706 , \36703 , \36362 );
nand \U$36364 ( \36707 , \36705 , \36706 );
and \U$36365 ( \36708 , \36701 , \36707 );
not \U$36366 ( \36709 , \36707 );
not \U$36367 ( \36710 , \36701 );
and \U$36368 ( \36711 , \36709 , \36710 );
xor \U$36369 ( \36712 , \36332 , \36333 );
xor \U$36370 ( \36713 , \36712 , \36342 );
nor \U$36371 ( \36714 , \36711 , \36713 );
nor \U$36372 ( \36715 , \36708 , \36714 );
nor \U$36373 ( \36716 , \36699 , \36715 );
nor \U$36374 ( \36717 , \36696 , \36716 );
xor \U$36375 ( \36718 , \36345 , \36375 );
xor \U$36376 ( \36719 , \36718 , \36402 );
not \U$36377 ( \36720 , \36719 );
xor \U$36378 ( \36721 , \36272 , \36293 );
xor \U$36379 ( \36722 , \36721 , \36322 );
nand \U$36380 ( \36723 , \36720 , \36722 );
xor \U$36381 ( \36724 , \36717 , \36723 );
xor \U$36382 ( \36725 , \36465 , \36467 );
xor \U$36383 ( \36726 , \36725 , \36470 );
xor \U$36384 ( \36727 , \36110 , \36117 );
xor \U$36385 ( \36728 , \36727 , \36125 );
xor \U$36386 ( \36729 , \36408 , \36413 );
xor \U$36387 ( \36730 , \36728 , \36729 );
and \U$36388 ( \36731 , \36726 , \36730 );
not \U$36389 ( \36732 , \36726 );
not \U$36390 ( \36733 , \36730 );
and \U$36391 ( \36734 , \36732 , \36733 );
not \U$36392 ( \36735 , \4519 );
not \U$36393 ( \36736 , \36291 );
or \U$36394 ( \36737 , \36735 , \36736 );
or \U$36395 ( \36738 , \36291 , \4519 );
nand \U$36396 ( \36739 , \36737 , \36738 );
not \U$36397 ( \36740 , \36739 );
not \U$36398 ( \36741 , \36280 );
and \U$36399 ( \36742 , \36740 , \36741 );
and \U$36400 ( \36743 , \36739 , \36280 );
nor \U$36401 ( \36744 , \36742 , \36743 );
not \U$36402 ( \36745 , \36744 );
not \U$36403 ( \36746 , \36308 );
not \U$36404 ( \36747 , \36320 );
or \U$36405 ( \36748 , \36746 , \36747 );
or \U$36406 ( \36749 , \36308 , \36320 );
nand \U$36407 ( \36750 , \36748 , \36749 );
not \U$36408 ( \36751 , \36750 );
not \U$36409 ( \36752 , \36301 );
and \U$36410 ( \36753 , \36751 , \36752 );
and \U$36411 ( \36754 , \36750 , \36301 );
nor \U$36412 ( \36755 , \36753 , \36754 );
not \U$36413 ( \36756 , \36755 );
and \U$36414 ( \36757 , \36745 , \36756 );
and \U$36415 ( \36758 , \36744 , \36755 );
not \U$36416 ( \36759 , \36258 );
not \U$36417 ( \36760 , \36270 );
or \U$36418 ( \36761 , \36759 , \36760 );
or \U$36419 ( \36762 , \36258 , \36270 );
nand \U$36420 ( \36763 , \36761 , \36762 );
not \U$36421 ( \36764 , \36763 );
not \U$36422 ( \36765 , \36251 );
and \U$36423 ( \36766 , \36764 , \36765 );
and \U$36424 ( \36767 , \36763 , \36251 );
nor \U$36425 ( \36768 , \36766 , \36767 );
nor \U$36426 ( \36769 , \36758 , \36768 );
nor \U$36427 ( \36770 , \36757 , \36769 );
nor \U$36428 ( \36771 , \36734 , \36770 );
nor \U$36429 ( \36772 , \36731 , \36771 );
and \U$36430 ( \36773 , \36724 , \36772 );
and \U$36431 ( \36774 , \36717 , \36723 );
or \U$36432 ( \36775 , \36773 , \36774 );
or \U$36433 ( \36776 , \36532 , \36775 );
not \U$36434 ( \36777 , \36775 );
not \U$36435 ( \36778 , \36532 );
or \U$36436 ( \36779 , \36777 , \36778 );
xor \U$36437 ( \36780 , \36064 , \36131 );
xor \U$36438 ( \36781 , \36780 , \36143 );
xor \U$36439 ( \36782 , \36232 , \36239 );
xor \U$36440 ( \36783 , \36781 , \36782 );
nand \U$36441 ( \36784 , \36779 , \36783 );
nand \U$36442 ( \36785 , \36776 , \36784 );
xor \U$36443 ( \36786 , \36146 , \36151 );
xor \U$36444 ( \36787 , \36786 , \36191 );
xor \U$36445 ( \36788 , \36785 , \36787 );
xor \U$36446 ( \36789 , \36244 , \36477 );
xor \U$36447 ( \36790 , \36789 , \36482 );
and \U$36448 ( \36791 , \36788 , \36790 );
and \U$36449 ( \36792 , \36785 , \36787 );
or \U$36450 ( \36793 , \36791 , \36792 );
xor \U$36451 ( \36794 , \35979 , \36194 );
xor \U$36452 ( \36795 , \36794 , \36201 );
xor \U$36453 ( \36796 , \36228 , \36485 );
xor \U$36454 ( \36797 , \36795 , \36796 );
nand \U$36455 ( \36798 , \36793 , \36797 );
xor \U$36456 ( \36799 , \36509 , \36798 );
xor \U$36457 ( \36800 , \36793 , \36797 );
xor \U$36458 ( \36801 , \36785 , \36787 );
xor \U$36459 ( \36802 , \36801 , \36790 );
not \U$36460 ( \36803 , \36802 );
xnor \U$36461 ( \36804 , \36775 , \36532 );
not \U$36462 ( \36805 , \36804 );
not \U$36463 ( \36806 , \36783 );
and \U$36464 ( \36807 , \36805 , \36806 );
and \U$36465 ( \36808 , \36804 , \36783 );
nor \U$36466 ( \36809 , \36807 , \36808 );
not \U$36467 ( \36810 , \36421 );
not \U$36468 ( \36811 , \36475 );
or \U$36469 ( \36812 , \36810 , \36811 );
or \U$36470 ( \36813 , \36475 , \36421 );
nand \U$36471 ( \36814 , \36812 , \36813 );
not \U$36472 ( \36815 , \36814 );
not \U$36473 ( \36816 , \36435 );
and \U$36474 ( \36817 , \36815 , \36816 );
and \U$36475 ( \36818 , \36814 , \36435 );
nor \U$36476 ( \36819 , \36817 , \36818 );
xor \U$36477 ( \36820 , \36809 , \36819 );
not \U$36478 ( \36821 , \36516 );
not \U$36479 ( \36822 , \36530 );
not \U$36480 ( \36823 , \36511 );
and \U$36481 ( \36824 , \36822 , \36823 );
and \U$36482 ( \36825 , \36530 , \36511 );
nor \U$36483 ( \36826 , \36824 , \36825 );
not \U$36484 ( \36827 , \36826 );
or \U$36485 ( \36828 , \36821 , \36827 );
or \U$36486 ( \36829 , \36826 , \36516 );
nand \U$36487 ( \36830 , \36828 , \36829 );
not \U$36488 ( \36831 , \454 );
and \U$36489 ( \36832 , \465 , RI986ec38_34);
and \U$36490 ( \36833 , RI986ed28_36, \463 );
nor \U$36491 ( \36834 , \36832 , \36833 );
not \U$36492 ( \36835 , \36834 );
or \U$36493 ( \36836 , \36831 , \36835 );
or \U$36494 ( \36837 , \36834 , \454 );
nand \U$36495 ( \36838 , \36836 , \36837 );
and \U$36496 ( \36839 , \438 , RI986f0e8_44);
and \U$36497 ( \36840 , RI986eff8_42, \436 );
nor \U$36498 ( \36841 , \36839 , \36840 );
and \U$36499 ( \36842 , \36841 , \444 );
not \U$36500 ( \36843 , \36841 );
and \U$36501 ( \36844 , \36843 , \443 );
nor \U$36502 ( \36845 , \36842 , \36844 );
xor \U$36503 ( \36846 , \36838 , \36845 );
not \U$36504 ( \36847 , \367 );
and \U$36505 ( \36848 , \376 , RI986ef08_40);
and \U$36506 ( \36849 , RI986ee18_38, \374 );
nor \U$36507 ( \36850 , \36848 , \36849 );
not \U$36508 ( \36851 , \36850 );
or \U$36509 ( \36852 , \36847 , \36851 );
or \U$36510 ( \36853 , \36850 , \365 );
nand \U$36511 ( \36854 , \36852 , \36853 );
and \U$36512 ( \36855 , \36846 , \36854 );
and \U$36513 ( \36856 , \36838 , \36845 );
or \U$36514 ( \36857 , \36855 , \36856 );
not \U$36515 ( \36858 , \345 );
and \U$36516 ( \36859 , \354 , RI986eb48_32);
and \U$36517 ( \36860 , RI986ea58_30, \352 );
nor \U$36518 ( \36861 , \36859 , \36860 );
not \U$36519 ( \36862 , \36861 );
or \U$36520 ( \36863 , \36858 , \36862 );
or \U$36521 ( \36864 , \36861 , \361 );
nand \U$36522 ( \36865 , \36863 , \36864 );
not \U$36523 ( \36866 , \487 );
and \U$36524 ( \36867 , \395 , RI986e968_28);
and \U$36525 ( \36868 , RI986e878_26, \393 );
nor \U$36526 ( \36869 , \36867 , \36868 );
not \U$36527 ( \36870 , \36869 );
or \U$36528 ( \36871 , \36866 , \36870 );
or \U$36529 ( \36872 , \36869 , \386 );
nand \U$36530 ( \36873 , \36871 , \36872 );
xor \U$36531 ( \36874 , \36865 , \36873 );
and \U$36532 ( \36875 , \416 , RI9871578_122);
and \U$36533 ( \36876 , RI9871668_124, \414 );
nor \U$36534 ( \36877 , \36875 , \36876 );
and \U$36535 ( \36878 , \36877 , \422 );
not \U$36536 ( \36879 , \36877 );
and \U$36537 ( \36880 , \36879 , \421 );
nor \U$36538 ( \36881 , \36878 , \36880 );
and \U$36539 ( \36882 , \36874 , \36881 );
and \U$36540 ( \36883 , \36865 , \36873 );
or \U$36541 ( \36884 , \36882 , \36883 );
xor \U$36542 ( \36885 , \36857 , \36884 );
and \U$36543 ( \36886 , \1329 , RI986e788_24);
and \U$36544 ( \36887 , RI986e698_22, \1327 );
nor \U$36545 ( \36888 , \36886 , \36887 );
and \U$36546 ( \36889 , \36888 , \1336 );
not \U$36547 ( \36890 , \36888 );
and \U$36548 ( \36891 , \36890 , \1337 );
nor \U$36549 ( \36892 , \36889 , \36891 );
and \U$36550 ( \36893 , \776 , RI986f2c8_48);
and \U$36551 ( \36894 , RI986f1d8_46, \774 );
nor \U$36552 ( \36895 , \36893 , \36894 );
and \U$36553 ( \36896 , \36895 , \474 );
not \U$36554 ( \36897 , \36895 );
and \U$36555 ( \36898 , \36897 , \451 );
nor \U$36556 ( \36899 , \36896 , \36898 );
xor \U$36557 ( \36900 , \36892 , \36899 );
not \U$36558 ( \36901 , \1128 );
and \U$36559 ( \36902 , \1293 , RI986e5a8_20);
and \U$36560 ( \36903 , RI986e4b8_18, \1291 );
nor \U$36561 ( \36904 , \36902 , \36903 );
not \U$36562 ( \36905 , \36904 );
or \U$36563 ( \36906 , \36901 , \36905 );
or \U$36564 ( \36907 , \36904 , \1301 );
nand \U$36565 ( \36908 , \36906 , \36907 );
and \U$36566 ( \36909 , \36900 , \36908 );
and \U$36567 ( \36910 , \36892 , \36899 );
or \U$36568 ( \36911 , \36909 , \36910 );
and \U$36569 ( \36912 , \36885 , \36911 );
and \U$36570 ( \36913 , \36857 , \36884 );
or \U$36571 ( \36914 , \36912 , \36913 );
not \U$36572 ( \36915 , \36651 );
not \U$36573 ( \36916 , \36663 );
or \U$36574 ( \36917 , \36915 , \36916 );
or \U$36575 ( \36918 , \36651 , \36663 );
nand \U$36576 ( \36919 , \36917 , \36918 );
not \U$36577 ( \36920 , \36919 );
not \U$36578 ( \36921 , \36652 );
and \U$36579 ( \36922 , \36920 , \36921 );
and \U$36580 ( \36923 , \36919 , \36652 );
nor \U$36581 ( \36924 , \36922 , \36923 );
not \U$36582 ( \36925 , \36621 );
not \U$36583 ( \36926 , \36641 );
or \U$36584 ( \36927 , \36925 , \36926 );
or \U$36585 ( \36928 , \36621 , \36641 );
nand \U$36586 ( \36929 , \36927 , \36928 );
not \U$36587 ( \36930 , \36929 );
not \U$36588 ( \36931 , \36629 );
and \U$36589 ( \36932 , \36930 , \36931 );
and \U$36590 ( \36933 , \36929 , \36629 );
nor \U$36591 ( \36934 , \36932 , \36933 );
nand \U$36592 ( \36935 , \36924 , \36934 );
xor \U$36593 ( \36936 , \36914 , \36935 );
and \U$36594 ( \36937 , \2274 , RI986f4a8_52);
and \U$36595 ( \36938 , RI986f3b8_50, \2272 );
nor \U$36596 ( \36939 , \36937 , \36938 );
and \U$36597 ( \36940 , \36939 , \2030 );
not \U$36598 ( \36941 , \36939 );
and \U$36599 ( \36942 , \36941 , \2031 );
nor \U$36600 ( \36943 , \36940 , \36942 );
and \U$36601 ( \36944 , \1311 , RI986f868_60);
and \U$36602 ( \36945 , RI986f778_58, \1309 );
nor \U$36603 ( \36946 , \36944 , \36945 );
and \U$36604 ( \36947 , \36946 , \1458 );
not \U$36605 ( \36948 , \36946 );
and \U$36606 ( \36949 , \36948 , \1318 );
nor \U$36607 ( \36950 , \36947 , \36949 );
xor \U$36608 ( \36951 , \36943 , \36950 );
not \U$36609 ( \36952 , \2034 );
and \U$36610 ( \36953 , \2042 , RI986fa48_64);
and \U$36611 ( \36954 , RI986f958_62, \2040 );
nor \U$36612 ( \36955 , \36953 , \36954 );
not \U$36613 ( \36956 , \36955 );
or \U$36614 ( \36957 , \36952 , \36956 );
or \U$36615 ( \36958 , \36955 , \2034 );
nand \U$36616 ( \36959 , \36957 , \36958 );
and \U$36617 ( \36960 , \36951 , \36959 );
and \U$36618 ( \36961 , \36943 , \36950 );
or \U$36619 ( \36962 , \36960 , \36961 );
and \U$36620 ( \36963 , \4203 , RI986e1e8_12);
and \U$36621 ( \36964 , RI986e0f8_10, \4201 );
nor \U$36622 ( \36965 , \36963 , \36964 );
and \U$36623 ( \36966 , \36965 , \4207 );
not \U$36624 ( \36967 , \36965 );
and \U$36625 ( \36968 , \36967 , \3922 );
nor \U$36626 ( \36969 , \36966 , \36968 );
xor \U$36627 ( \36970 , \36969 , \5052 );
not \U$36628 ( \36971 , \4521 );
and \U$36629 ( \36972 , \4710 , RI986e2d8_14);
and \U$36630 ( \36973 , RI986e3c8_16, \4708 );
nor \U$36631 ( \36974 , \36972 , \36973 );
not \U$36632 ( \36975 , \36974 );
or \U$36633 ( \36976 , \36971 , \36975 );
or \U$36634 ( \36977 , \36974 , \4521 );
nand \U$36635 ( \36978 , \36976 , \36977 );
and \U$36636 ( \36979 , \36970 , \36978 );
and \U$36637 ( \36980 , \36969 , \5052 );
or \U$36638 ( \36981 , \36979 , \36980 );
xor \U$36639 ( \36982 , \36962 , \36981 );
and \U$36640 ( \36983 , \2464 , RI986f598_54);
and \U$36641 ( \36984 , RI986f688_56, \2462 );
nor \U$36642 ( \36985 , \36983 , \36984 );
and \U$36643 ( \36986 , \36985 , \2468 );
not \U$36644 ( \36987 , \36985 );
and \U$36645 ( \36988 , \36987 , \2263 );
nor \U$36646 ( \36989 , \36986 , \36988 );
not \U$36647 ( \36990 , \3406 );
and \U$36648 ( \36991 , \3254 , RI986e008_8);
and \U$36649 ( \36992 , RI986df18_6, \3252 );
nor \U$36650 ( \36993 , \36991 , \36992 );
not \U$36651 ( \36994 , \36993 );
or \U$36652 ( \36995 , \36990 , \36994 );
or \U$36653 ( \36996 , \36993 , \2935 );
nand \U$36654 ( \36997 , \36995 , \36996 );
xor \U$36655 ( \36998 , \36989 , \36997 );
not \U$36656 ( \36999 , \3412 );
and \U$36657 ( \37000 , \3683 , RI986de28_4);
and \U$36658 ( \37001 , RI986dd38_2, \3681 );
nor \U$36659 ( \37002 , \37000 , \37001 );
not \U$36660 ( \37003 , \37002 );
or \U$36661 ( \37004 , \36999 , \37003 );
or \U$36662 ( \37005 , \37002 , \3412 );
nand \U$36663 ( \37006 , \37004 , \37005 );
and \U$36664 ( \37007 , \36998 , \37006 );
and \U$36665 ( \37008 , \36989 , \36997 );
or \U$36666 ( \37009 , \37007 , \37008 );
and \U$36667 ( \37010 , \36982 , \37009 );
and \U$36668 ( \37011 , \36962 , \36981 );
or \U$36669 ( \37012 , \37010 , \37011 );
and \U$36670 ( \37013 , \36936 , \37012 );
and \U$36671 ( \37014 , \36914 , \36935 );
or \U$36672 ( \37015 , \37013 , \37014 );
xor \U$36673 ( \37016 , \36558 , \36583 );
xor \U$36674 ( \37017 , \37016 , \36610 );
xor \U$36675 ( \37018 , \36643 , \36665 );
xor \U$36676 ( \37019 , \37018 , \36692 );
and \U$36677 ( \37020 , \37017 , \37019 );
xor \U$36678 ( \37021 , \37015 , \37020 );
not \U$36679 ( \37022 , \36701 );
not \U$36680 ( \37023 , \36707 );
not \U$36681 ( \37024 , \36713 );
and \U$36682 ( \37025 , \37023 , \37024 );
and \U$36683 ( \37026 , \36707 , \36713 );
nor \U$36684 ( \37027 , \37025 , \37026 );
not \U$36685 ( \37028 , \37027 );
or \U$36686 ( \37029 , \37022 , \37028 );
or \U$36687 ( \37030 , \37027 , \36701 );
nand \U$36688 ( \37031 , \37029 , \37030 );
xor \U$36689 ( \37032 , \36591 , \36598 );
xor \U$36690 ( \37033 , \37032 , \36607 );
xor \U$36691 ( \37034 , \36673 , \36680 );
xor \U$36692 ( \37035 , \37034 , \36689 );
and \U$36693 ( \37036 , \37033 , \37035 );
xor \U$36694 ( \37037 , \36539 , \36546 );
xor \U$36695 ( \37038 , \37037 , \36555 );
xor \U$36696 ( \37039 , \36673 , \36680 );
xor \U$36697 ( \37040 , \37039 , \36689 );
and \U$36698 ( \37041 , \37038 , \37040 );
and \U$36699 ( \37042 , \37033 , \37038 );
or \U$36700 ( \37043 , \37036 , \37041 , \37042 );
xor \U$36701 ( \37044 , \37031 , \37043 );
not \U$36702 ( \37045 , \36744 );
xor \U$36703 ( \37046 , \36768 , \36755 );
not \U$36704 ( \37047 , \37046 );
or \U$36705 ( \37048 , \37045 , \37047 );
or \U$36706 ( \37049 , \37046 , \36744 );
nand \U$36707 ( \37050 , \37048 , \37049 );
and \U$36708 ( \37051 , \37044 , \37050 );
and \U$36709 ( \37052 , \37031 , \37043 );
or \U$36710 ( \37053 , \37051 , \37052 );
and \U$36711 ( \37054 , \37021 , \37053 );
and \U$36712 ( \37055 , \37015 , \37020 );
or \U$36713 ( \37056 , \37054 , \37055 );
xor \U$36714 ( \37057 , \36830 , \37056 );
not \U$36715 ( \37058 , \36715 );
xor \U$36716 ( \37059 , \36613 , \36695 );
not \U$36717 ( \37060 , \37059 );
or \U$36718 ( \37061 , \37058 , \37060 );
or \U$36719 ( \37062 , \37059 , \36715 );
nand \U$36720 ( \37063 , \37061 , \37062 );
not \U$36721 ( \37064 , \36722 );
not \U$36722 ( \37065 , \36719 );
or \U$36723 ( \37066 , \37064 , \37065 );
or \U$36724 ( \37067 , \36719 , \36722 );
nand \U$36725 ( \37068 , \37066 , \37067 );
xor \U$36726 ( \37069 , \37063 , \37068 );
not \U$36727 ( \37070 , \36730 );
not \U$36728 ( \37071 , \36726 );
not \U$36729 ( \37072 , \36770 );
and \U$36730 ( \37073 , \37071 , \37072 );
and \U$36731 ( \37074 , \36726 , \36770 );
nor \U$36732 ( \37075 , \37073 , \37074 );
not \U$36733 ( \37076 , \37075 );
or \U$36734 ( \37077 , \37070 , \37076 );
or \U$36735 ( \37078 , \37075 , \36730 );
nand \U$36736 ( \37079 , \37077 , \37078 );
and \U$36737 ( \37080 , \37069 , \37079 );
and \U$36738 ( \37081 , \37063 , \37068 );
or \U$36739 ( \37082 , \37080 , \37081 );
and \U$36740 ( \37083 , \37057 , \37082 );
and \U$36741 ( \37084 , \36830 , \37056 );
nor \U$36742 ( \37085 , \37083 , \37084 );
and \U$36743 ( \37086 , \36820 , \37085 );
and \U$36744 ( \37087 , \36809 , \36819 );
or \U$36745 ( \37088 , \37086 , \37087 );
nor \U$36746 ( \37089 , \36803 , \37088 );
and \U$36747 ( \37090 , \36800 , \37089 );
xor \U$36748 ( \37091 , \37089 , \36800 );
and \U$36749 ( \37092 , \416 , RI9871758_126);
and \U$36750 ( \37093 , RI9871848_128, \414 );
nor \U$36751 ( \37094 , \37092 , \37093 );
and \U$36752 ( \37095 , \37094 , \422 );
not \U$36753 ( \37096 , \37094 );
and \U$36754 ( \37097 , \37096 , \421 );
nor \U$36755 ( \37098 , \37095 , \37097 );
not \U$36756 ( \37099 , RI9871488_120);
nor \U$36757 ( \37100 , \37099 , \407 );
xor \U$36758 ( \37101 , \37098 , \37100 );
nand \U$36759 ( \37102 , RI9871398_118, RI9871fc8_144);
and \U$36760 ( \37103 , \416 , RI9871488_120);
and \U$36761 ( \37104 , RI9871758_126, \414 );
nor \U$36762 ( \37105 , \37103 , \37104 );
and \U$36763 ( \37106 , \37105 , \421 );
not \U$36764 ( \37107 , \37105 );
and \U$36765 ( \37108 , \37107 , \422 );
nor \U$36766 ( \37109 , \37106 , \37108 );
nand \U$36767 ( \37110 , \37102 , \37109 );
xor \U$36768 ( \37111 , \37101 , \37110 );
not \U$36769 ( \37112 , \454 );
and \U$36770 ( \37113 , \465 , RI986e878_26);
and \U$36771 ( \37114 , RI986ef08_40, \463 );
nor \U$36772 ( \37115 , \37113 , \37114 );
not \U$36773 ( \37116 , \37115 );
or \U$36774 ( \37117 , \37112 , \37116 );
or \U$36775 ( \37118 , \37115 , \456 );
nand \U$36776 ( \37119 , \37117 , \37118 );
and \U$36777 ( \37120 , \776 , RI986ed28_36);
and \U$36778 ( \37121 , RI986f0e8_44, \774 );
nor \U$36779 ( \37122 , \37120 , \37121 );
and \U$36780 ( \37123 , \37122 , \474 );
not \U$36781 ( \37124 , \37122 );
and \U$36782 ( \37125 , \37124 , \451 );
nor \U$36783 ( \37126 , \37123 , \37125 );
xor \U$36784 ( \37127 , \37119 , \37126 );
and \U$36785 ( \37128 , \438 , RI986ee18_38);
and \U$36786 ( \37129 , RI986ec38_34, \436 );
nor \U$36787 ( \37130 , \37128 , \37129 );
and \U$36788 ( \37131 , \37130 , \444 );
not \U$36789 ( \37132 , \37130 );
and \U$36790 ( \37133 , \37132 , \443 );
nor \U$36791 ( \37134 , \37131 , \37133 );
and \U$36792 ( \37135 , \37127 , \37134 );
and \U$36793 ( \37136 , \37119 , \37126 );
or \U$36794 ( \37137 , \37135 , \37136 );
not \U$36795 ( \37138 , \487 );
and \U$36796 ( \37139 , \395 , RI9871668_124);
and \U$36797 ( \37140 , RI986eb48_32, \393 );
nor \U$36798 ( \37141 , \37139 , \37140 );
not \U$36799 ( \37142 , \37141 );
or \U$36800 ( \37143 , \37138 , \37142 );
or \U$36801 ( \37144 , \37141 , \487 );
nand \U$36802 ( \37145 , \37143 , \37144 );
not \U$36803 ( \37146 , \367 );
and \U$36804 ( \37147 , \376 , RI986ea58_30);
and \U$36805 ( \37148 , RI986e968_28, \374 );
nor \U$36806 ( \37149 , \37147 , \37148 );
not \U$36807 ( \37150 , \37149 );
or \U$36808 ( \37151 , \37146 , \37150 );
or \U$36809 ( \37152 , \37149 , \365 );
nand \U$36810 ( \37153 , \37151 , \37152 );
xor \U$36811 ( \37154 , \37145 , \37153 );
not \U$36812 ( \37155 , \361 );
and \U$36813 ( \37156 , \354 , RI9871848_128);
and \U$36814 ( \37157 , RI9871578_122, \352 );
nor \U$36815 ( \37158 , \37156 , \37157 );
not \U$36816 ( \37159 , \37158 );
or \U$36817 ( \37160 , \37155 , \37159 );
or \U$36818 ( \37161 , \37158 , \361 );
nand \U$36819 ( \37162 , \37160 , \37161 );
and \U$36820 ( \37163 , \37154 , \37162 );
and \U$36821 ( \37164 , \37145 , \37153 );
or \U$36822 ( \37165 , \37163 , \37164 );
xor \U$36823 ( \37166 , \37137 , \37165 );
not \U$36824 ( \37167 , \1301 );
and \U$36825 ( \37168 , \1293 , RI986eff8_42);
and \U$36826 ( \37169 , RI986f2c8_48, \1291 );
nor \U$36827 ( \37170 , \37168 , \37169 );
not \U$36828 ( \37171 , \37170 );
or \U$36829 ( \37172 , \37167 , \37171 );
or \U$36830 ( \37173 , \37170 , \1301 );
nand \U$36831 ( \37174 , \37172 , \37173 );
and \U$36832 ( \37175 , \1329 , RI986f1d8_46);
and \U$36833 ( \37176 , RI986e5a8_20, \1327 );
nor \U$36834 ( \37177 , \37175 , \37176 );
and \U$36835 ( \37178 , \37177 , \1336 );
not \U$36836 ( \37179 , \37177 );
and \U$36837 ( \37180 , \37179 , \1337 );
nor \U$36838 ( \37181 , \37178 , \37180 );
xor \U$36839 ( \37182 , \37174 , \37181 );
and \U$36840 ( \37183 , \1311 , RI986e4b8_18);
and \U$36841 ( \37184 , RI986e788_24, \1309 );
nor \U$36842 ( \37185 , \37183 , \37184 );
and \U$36843 ( \37186 , \37185 , \1458 );
not \U$36844 ( \37187 , \37185 );
and \U$36845 ( \37188 , \37187 , \1318 );
nor \U$36846 ( \37189 , \37186 , \37188 );
and \U$36847 ( \37190 , \37182 , \37189 );
and \U$36848 ( \37191 , \37174 , \37181 );
or \U$36849 ( \37192 , \37190 , \37191 );
xor \U$36850 ( \37193 , \37166 , \37192 );
and \U$36851 ( \37194 , \37111 , \37193 );
not \U$36852 ( \37195 , \361 );
and \U$36853 ( \37196 , \354 , RI9871578_122);
and \U$36854 ( \37197 , RI9871668_124, \352 );
nor \U$36855 ( \37198 , \37196 , \37197 );
not \U$36856 ( \37199 , \37198 );
or \U$36857 ( \37200 , \37195 , \37199 );
or \U$36858 ( \37201 , \37198 , \345 );
nand \U$36859 ( \37202 , \37200 , \37201 );
not \U$36860 ( \37203 , \365 );
and \U$36861 ( \37204 , \376 , RI986e968_28);
and \U$36862 ( \37205 , RI986e878_26, \374 );
nor \U$36863 ( \37206 , \37204 , \37205 );
not \U$36864 ( \37207 , \37206 );
or \U$36865 ( \37208 , \37203 , \37207 );
or \U$36866 ( \37209 , \37206 , \367 );
nand \U$36867 ( \37210 , \37208 , \37209 );
xor \U$36868 ( \37211 , \37202 , \37210 );
not \U$36869 ( \37212 , \487 );
and \U$36870 ( \37213 , \395 , RI986eb48_32);
and \U$36871 ( \37214 , RI986ea58_30, \393 );
nor \U$36872 ( \37215 , \37213 , \37214 );
not \U$36873 ( \37216 , \37215 );
or \U$36874 ( \37217 , \37212 , \37216 );
or \U$36875 ( \37218 , \37215 , \487 );
nand \U$36876 ( \37219 , \37217 , \37218 );
xor \U$36877 ( \37220 , \37211 , \37219 );
not \U$36878 ( \37221 , \456 );
and \U$36879 ( \37222 , \465 , RI986ef08_40);
and \U$36880 ( \37223 , RI986ee18_38, \463 );
nor \U$36881 ( \37224 , \37222 , \37223 );
not \U$36882 ( \37225 , \37224 );
or \U$36883 ( \37226 , \37221 , \37225 );
or \U$36884 ( \37227 , \37224 , \456 );
nand \U$36885 ( \37228 , \37226 , \37227 );
and \U$36886 ( \37229 , \776 , RI986f0e8_44);
and \U$36887 ( \37230 , RI986eff8_42, \774 );
nor \U$36888 ( \37231 , \37229 , \37230 );
and \U$36889 ( \37232 , \37231 , \474 );
not \U$36890 ( \37233 , \37231 );
and \U$36891 ( \37234 , \37233 , \451 );
nor \U$36892 ( \37235 , \37232 , \37234 );
xor \U$36893 ( \37236 , \37228 , \37235 );
and \U$36894 ( \37237 , \438 , RI986ec38_34);
and \U$36895 ( \37238 , RI986ed28_36, \436 );
nor \U$36896 ( \37239 , \37237 , \37238 );
and \U$36897 ( \37240 , \37239 , \444 );
not \U$36898 ( \37241 , \37239 );
and \U$36899 ( \37242 , \37241 , \443 );
nor \U$36900 ( \37243 , \37240 , \37242 );
xor \U$36901 ( \37244 , \37236 , \37243 );
not \U$36902 ( \37245 , \1128 );
and \U$36903 ( \37246 , \1293 , RI986f2c8_48);
and \U$36904 ( \37247 , RI986f1d8_46, \1291 );
nor \U$36905 ( \37248 , \37246 , \37247 );
not \U$36906 ( \37249 , \37248 );
or \U$36907 ( \37250 , \37245 , \37249 );
or \U$36908 ( \37251 , \37248 , \1301 );
nand \U$36909 ( \37252 , \37250 , \37251 );
and \U$36910 ( \37253 , \1329 , RI986e5a8_20);
and \U$36911 ( \37254 , RI986e4b8_18, \1327 );
nor \U$36912 ( \37255 , \37253 , \37254 );
and \U$36913 ( \37256 , \37255 , \1336 );
not \U$36914 ( \37257 , \37255 );
and \U$36915 ( \37258 , \37257 , \1337 );
nor \U$36916 ( \37259 , \37256 , \37258 );
xor \U$36917 ( \37260 , \37252 , \37259 );
and \U$36918 ( \37261 , \1311 , RI986e788_24);
and \U$36919 ( \37262 , RI986e698_22, \1309 );
nor \U$36920 ( \37263 , \37261 , \37262 );
and \U$36921 ( \37264 , \37263 , \1458 );
not \U$36922 ( \37265 , \37263 );
and \U$36923 ( \37266 , \37265 , \1318 );
nor \U$36924 ( \37267 , \37264 , \37266 );
xor \U$36925 ( \37268 , \37260 , \37267 );
xor \U$36926 ( \37269 , \37244 , \37268 );
xor \U$36927 ( \37270 , \37220 , \37269 );
xor \U$36928 ( \37271 , \37137 , \37165 );
xor \U$36929 ( \37272 , \37271 , \37192 );
and \U$36930 ( \37273 , \37270 , \37272 );
and \U$36931 ( \37274 , \37111 , \37270 );
or \U$36932 ( \37275 , \37194 , \37273 , \37274 );
and \U$36933 ( \37276 , \776 , RI986ec38_34);
and \U$36934 ( \37277 , RI986ed28_36, \774 );
nor \U$36935 ( \37278 , \37276 , \37277 );
and \U$36936 ( \37279 , \37278 , \474 );
not \U$36937 ( \37280 , \37278 );
and \U$36938 ( \37281 , \37280 , \451 );
nor \U$36939 ( \37282 , \37279 , \37281 );
and \U$36940 ( \37283 , \438 , RI986ef08_40);
and \U$36941 ( \37284 , RI986ee18_38, \436 );
nor \U$36942 ( \37285 , \37283 , \37284 );
and \U$36943 ( \37286 , \37285 , \444 );
not \U$36944 ( \37287 , \37285 );
and \U$36945 ( \37288 , \37287 , \443 );
nor \U$36946 ( \37289 , \37286 , \37288 );
xor \U$36947 ( \37290 , \37282 , \37289 );
not \U$36948 ( \37291 , \1128 );
and \U$36949 ( \37292 , \1293 , RI986f0e8_44);
and \U$36950 ( \37293 , RI986eff8_42, \1291 );
nor \U$36951 ( \37294 , \37292 , \37293 );
not \U$36952 ( \37295 , \37294 );
or \U$36953 ( \37296 , \37291 , \37295 );
or \U$36954 ( \37297 , \37294 , \1301 );
nand \U$36955 ( \37298 , \37296 , \37297 );
and \U$36956 ( \37299 , \37290 , \37298 );
and \U$36957 ( \37300 , \37282 , \37289 );
or \U$36958 ( \37301 , \37299 , \37300 );
not \U$36959 ( \37302 , \487 );
and \U$36960 ( \37303 , \395 , RI9871578_122);
and \U$36961 ( \37304 , RI9871668_124, \393 );
nor \U$36962 ( \37305 , \37303 , \37304 );
not \U$36963 ( \37306 , \37305 );
or \U$36964 ( \37307 , \37302 , \37306 );
or \U$36965 ( \37308 , \37305 , \386 );
nand \U$36966 ( \37309 , \37307 , \37308 );
not \U$36967 ( \37310 , \454 );
and \U$36968 ( \37311 , \465 , RI986e968_28);
and \U$36969 ( \37312 , RI986e878_26, \463 );
nor \U$36970 ( \37313 , \37311 , \37312 );
not \U$36971 ( \37314 , \37313 );
or \U$36972 ( \37315 , \37310 , \37314 );
or \U$36973 ( \37316 , \37313 , \456 );
nand \U$36974 ( \37317 , \37315 , \37316 );
xor \U$36975 ( \37318 , \37309 , \37317 );
not \U$36976 ( \37319 , \365 );
and \U$36977 ( \37320 , \376 , RI986eb48_32);
and \U$36978 ( \37321 , RI986ea58_30, \374 );
nor \U$36979 ( \37322 , \37320 , \37321 );
not \U$36980 ( \37323 , \37322 );
or \U$36981 ( \37324 , \37319 , \37323 );
or \U$36982 ( \37325 , \37322 , \365 );
nand \U$36983 ( \37326 , \37324 , \37325 );
and \U$36984 ( \37327 , \37318 , \37326 );
and \U$36985 ( \37328 , \37309 , \37317 );
or \U$36986 ( \37329 , \37327 , \37328 );
xor \U$36987 ( \37330 , \37301 , \37329 );
and \U$36988 ( \37331 , \1311 , RI986e5a8_20);
and \U$36989 ( \37332 , RI986e4b8_18, \1309 );
nor \U$36990 ( \37333 , \37331 , \37332 );
and \U$36991 ( \37334 , \37333 , \1458 );
not \U$36992 ( \37335 , \37333 );
and \U$36993 ( \37336 , \37335 , \1318 );
nor \U$36994 ( \37337 , \37334 , \37336 );
and \U$36995 ( \37338 , \1329 , RI986f2c8_48);
and \U$36996 ( \37339 , RI986f1d8_46, \1327 );
nor \U$36997 ( \37340 , \37338 , \37339 );
and \U$36998 ( \37341 , \37340 , \1336 );
not \U$36999 ( \37342 , \37340 );
and \U$37000 ( \37343 , \37342 , \1337 );
nor \U$37001 ( \37344 , \37341 , \37343 );
xor \U$37002 ( \37345 , \37337 , \37344 );
not \U$37003 ( \37346 , \2034 );
and \U$37004 ( \37347 , \2042 , RI986e788_24);
and \U$37005 ( \37348 , RI986e698_22, \2040 );
nor \U$37006 ( \37349 , \37347 , \37348 );
not \U$37007 ( \37350 , \37349 );
or \U$37008 ( \37351 , \37346 , \37350 );
or \U$37009 ( \37352 , \37349 , \2034 );
nand \U$37010 ( \37353 , \37351 , \37352 );
and \U$37011 ( \37354 , \37345 , \37353 );
and \U$37012 ( \37355 , \37337 , \37344 );
or \U$37013 ( \37356 , \37354 , \37355 );
and \U$37014 ( \37357 , \37330 , \37356 );
and \U$37015 ( \37358 , \37301 , \37329 );
or \U$37016 ( \37359 , \37357 , \37358 );
not \U$37017 ( \37360 , \3918 );
and \U$37018 ( \37361 , \3683 , RI986f598_54);
and \U$37019 ( \37362 , RI986f688_56, \3681 );
nor \U$37020 ( \37363 , \37361 , \37362 );
not \U$37021 ( \37364 , \37363 );
or \U$37022 ( \37365 , \37360 , \37364 );
or \U$37023 ( \37366 , \37363 , \3918 );
nand \U$37024 ( \37367 , \37365 , \37366 );
and \U$37025 ( \37368 , \4203 , RI986e008_8);
and \U$37026 ( \37369 , RI986df18_6, \4201 );
nor \U$37027 ( \37370 , \37368 , \37369 );
and \U$37028 ( \37371 , \37370 , \4207 );
not \U$37029 ( \37372 , \37370 );
and \U$37030 ( \37373 , \37372 , \3923 );
nor \U$37031 ( \37374 , \37371 , \37373 );
xor \U$37032 ( \37375 , \37367 , \37374 );
not \U$37033 ( \37376 , \4521 );
and \U$37034 ( \37377 , \4710 , RI986de28_4);
and \U$37035 ( \37378 , RI986dd38_2, \4708 );
nor \U$37036 ( \37379 , \37377 , \37378 );
not \U$37037 ( \37380 , \37379 );
or \U$37038 ( \37381 , \37376 , \37380 );
or \U$37039 ( \37382 , \37379 , \4519 );
nand \U$37040 ( \37383 , \37381 , \37382 );
and \U$37041 ( \37384 , \37375 , \37383 );
and \U$37042 ( \37385 , \37367 , \37374 );
or \U$37043 ( \37386 , \37384 , \37385 );
and \U$37044 ( \37387 , \5318 , RI986e1e8_12);
and \U$37045 ( \37388 , RI986e0f8_10, \5316 );
nor \U$37046 ( \37389 , \37387 , \37388 );
and \U$37047 ( \37390 , \37389 , \5052 );
not \U$37048 ( \37391 , \37389 );
and \U$37049 ( \37392 , \37391 , \5322 );
nor \U$37050 ( \37393 , \37390 , \37392 );
xor \U$37051 ( \37394 , \37393 , \6190 );
and \U$37052 ( \37395 , \5881 , RI986e2d8_14);
and \U$37053 ( \37396 , RI986e3c8_16, \5879 );
nor \U$37054 ( \37397 , \37395 , \37396 );
and \U$37055 ( \37398 , \37397 , \5594 );
not \U$37056 ( \37399 , \37397 );
and \U$37057 ( \37400 , \37399 , \5885 );
nor \U$37058 ( \37401 , \37398 , \37400 );
and \U$37059 ( \37402 , \37394 , \37401 );
and \U$37060 ( \37403 , \37393 , \6190 );
or \U$37061 ( \37404 , \37402 , \37403 );
xor \U$37062 ( \37405 , \37386 , \37404 );
and \U$37063 ( \37406 , \2274 , RI986f868_60);
and \U$37064 ( \37407 , RI986f778_58, \2272 );
nor \U$37065 ( \37408 , \37406 , \37407 );
and \U$37066 ( \37409 , \37408 , \2030 );
not \U$37067 ( \37410 , \37408 );
and \U$37068 ( \37411 , \37410 , \2031 );
nor \U$37069 ( \37412 , \37409 , \37411 );
and \U$37070 ( \37413 , \2464 , RI986fa48_64);
and \U$37071 ( \37414 , RI986f958_62, \2462 );
nor \U$37072 ( \37415 , \37413 , \37414 );
and \U$37073 ( \37416 , \37415 , \2468 );
not \U$37074 ( \37417 , \37415 );
and \U$37075 ( \37418 , \37417 , \2263 );
nor \U$37076 ( \37419 , \37416 , \37418 );
xor \U$37077 ( \37420 , \37412 , \37419 );
not \U$37078 ( \37421 , \3406 );
and \U$37079 ( \37422 , \3254 , RI986f4a8_52);
and \U$37080 ( \37423 , RI986f3b8_50, \3252 );
nor \U$37081 ( \37424 , \37422 , \37423 );
not \U$37082 ( \37425 , \37424 );
or \U$37083 ( \37426 , \37421 , \37425 );
or \U$37084 ( \37427 , \37424 , \3406 );
nand \U$37085 ( \37428 , \37426 , \37427 );
and \U$37086 ( \37429 , \37420 , \37428 );
and \U$37087 ( \37430 , \37412 , \37419 );
or \U$37088 ( \37431 , \37429 , \37430 );
and \U$37089 ( \37432 , \37405 , \37431 );
and \U$37090 ( \37433 , \37386 , \37404 );
or \U$37091 ( \37434 , \37432 , \37433 );
xor \U$37092 ( \37435 , \37359 , \37434 );
and \U$37093 ( \37436 , \416 , RI9871398_118);
and \U$37094 ( \37437 , RI9871488_120, \414 );
nor \U$37095 ( \37438 , \37436 , \37437 );
and \U$37096 ( \37439 , \37438 , \422 );
not \U$37097 ( \37440 , \37438 );
and \U$37098 ( \37441 , \37440 , \421 );
nor \U$37099 ( \37442 , \37439 , \37441 );
not \U$37100 ( \37443 , RI98711b8_114);
nor \U$37101 ( \37444 , \37443 , \407 );
xor \U$37102 ( \37445 , \37442 , \37444 );
not \U$37103 ( \37446 , \361 );
and \U$37104 ( \37447 , \354 , RI9871758_126);
and \U$37105 ( \37448 , RI9871848_128, \352 );
nor \U$37106 ( \37449 , \37447 , \37448 );
not \U$37107 ( \37450 , \37449 );
or \U$37108 ( \37451 , \37446 , \37450 );
or \U$37109 ( \37452 , \37449 , \361 );
nand \U$37110 ( \37453 , \37451 , \37452 );
and \U$37111 ( \37454 , \37445 , \37453 );
and \U$37112 ( \37455 , \37442 , \37444 );
or \U$37113 ( \37456 , \37454 , \37455 );
or \U$37114 ( \37457 , \37109 , \37102 );
nand \U$37115 ( \37458 , \37457 , \37110 );
xor \U$37116 ( \37459 , \37456 , \37458 );
xor \U$37117 ( \37460 , \37145 , \37153 );
xor \U$37118 ( \37461 , \37460 , \37162 );
and \U$37119 ( \37462 , \37459 , \37461 );
and \U$37120 ( \37463 , \37456 , \37458 );
or \U$37121 ( \37464 , \37462 , \37463 );
and \U$37122 ( \37465 , \37435 , \37464 );
and \U$37123 ( \37466 , \37359 , \37434 );
or \U$37124 ( \37467 , \37465 , \37466 );
xor \U$37125 ( \37468 , \37275 , \37467 );
xor \U$37126 ( \37469 , \37174 , \37181 );
xor \U$37127 ( \37470 , \37469 , \37189 );
xor \U$37128 ( \37471 , \37119 , \37126 );
xor \U$37129 ( \37472 , \37471 , \37134 );
and \U$37130 ( \37473 , \37470 , \37472 );
not \U$37131 ( \37474 , \1462 );
and \U$37132 ( \37475 , \2042 , RI986e698_22);
and \U$37133 ( \37476 , RI986f868_60, \2040 );
nor \U$37134 ( \37477 , \37475 , \37476 );
not \U$37135 ( \37478 , \37477 );
or \U$37136 ( \37479 , \37474 , \37478 );
or \U$37137 ( \37480 , \37477 , \1462 );
nand \U$37138 ( \37481 , \37479 , \37480 );
and \U$37139 ( \37482 , \2274 , RI986f778_58);
and \U$37140 ( \37483 , RI986fa48_64, \2272 );
nor \U$37141 ( \37484 , \37482 , \37483 );
and \U$37142 ( \37485 , \37484 , \2030 );
not \U$37143 ( \37486 , \37484 );
and \U$37144 ( \37487 , \37486 , \2031 );
nor \U$37145 ( \37488 , \37485 , \37487 );
xor \U$37146 ( \37489 , \37481 , \37488 );
and \U$37147 ( \37490 , \2464 , RI986f958_62);
and \U$37148 ( \37491 , RI986f4a8_52, \2462 );
nor \U$37149 ( \37492 , \37490 , \37491 );
and \U$37150 ( \37493 , \37492 , \2468 );
not \U$37151 ( \37494 , \37492 );
and \U$37152 ( \37495 , \37494 , \2263 );
nor \U$37153 ( \37496 , \37493 , \37495 );
xor \U$37154 ( \37497 , \37489 , \37496 );
xor \U$37155 ( \37498 , \37119 , \37126 );
xor \U$37156 ( \37499 , \37498 , \37134 );
and \U$37157 ( \37500 , \37497 , \37499 );
and \U$37158 ( \37501 , \37470 , \37497 );
or \U$37159 ( \37502 , \37473 , \37500 , \37501 );
not \U$37160 ( \37503 , \3412 );
and \U$37161 ( \37504 , \3683 , RI986f688_56);
and \U$37162 ( \37505 , RI986e008_8, \3681 );
nor \U$37163 ( \37506 , \37504 , \37505 );
not \U$37164 ( \37507 , \37506 );
or \U$37165 ( \37508 , \37503 , \37507 );
or \U$37166 ( \37509 , \37506 , \3918 );
nand \U$37167 ( \37510 , \37508 , \37509 );
not \U$37168 ( \37511 , \2935 );
and \U$37169 ( \37512 , \3254 , RI986f3b8_50);
and \U$37170 ( \37513 , RI986f598_54, \3252 );
nor \U$37171 ( \37514 , \37512 , \37513 );
not \U$37172 ( \37515 , \37514 );
or \U$37173 ( \37516 , \37511 , \37515 );
or \U$37174 ( \37517 , \37514 , \2935 );
nand \U$37175 ( \37518 , \37516 , \37517 );
xor \U$37176 ( \37519 , \37510 , \37518 );
and \U$37177 ( \37520 , \4203 , RI986df18_6);
and \U$37178 ( \37521 , RI986de28_4, \4201 );
nor \U$37179 ( \37522 , \37520 , \37521 );
and \U$37180 ( \37523 , \37522 , \4207 );
not \U$37181 ( \37524 , \37522 );
and \U$37182 ( \37525 , \37524 , \3922 );
nor \U$37183 ( \37526 , \37523 , \37525 );
xor \U$37184 ( \37527 , \37519 , \37526 );
not \U$37185 ( \37528 , \4521 );
and \U$37186 ( \37529 , \4710 , RI986dd38_2);
and \U$37187 ( \37530 , RI986e1e8_12, \4708 );
nor \U$37188 ( \37531 , \37529 , \37530 );
not \U$37189 ( \37532 , \37531 );
or \U$37190 ( \37533 , \37528 , \37532 );
or \U$37191 ( \37534 , \37531 , \4521 );
nand \U$37192 ( \37535 , \37533 , \37534 );
nand \U$37193 ( \37536 , RI986e3c8_16, \5881 );
and \U$37194 ( \37537 , \37536 , \5594 );
not \U$37195 ( \37538 , \37536 );
and \U$37196 ( \37539 , \37538 , \5885 );
nor \U$37197 ( \37540 , \37537 , \37539 );
xor \U$37198 ( \37541 , \37535 , \37540 );
and \U$37199 ( \37542 , \5318 , RI986e0f8_10);
and \U$37200 ( \37543 , RI986e2d8_14, \5316 );
nor \U$37201 ( \37544 , \37542 , \37543 );
and \U$37202 ( \37545 , \37544 , \5052 );
not \U$37203 ( \37546 , \37544 );
and \U$37204 ( \37547 , \37546 , \5322 );
nor \U$37205 ( \37548 , \37545 , \37547 );
xor \U$37206 ( \37549 , \37541 , \37548 );
and \U$37207 ( \37550 , \37527 , \37549 );
xor \U$37208 ( \37551 , \37502 , \37550 );
not \U$37209 ( \37552 , \2935 );
and \U$37210 ( \37553 , \3254 , RI986f598_54);
and \U$37211 ( \37554 , RI986f688_56, \3252 );
nor \U$37212 ( \37555 , \37553 , \37554 );
not \U$37213 ( \37556 , \37555 );
or \U$37214 ( \37557 , \37552 , \37556 );
or \U$37215 ( \37558 , \37555 , \2935 );
nand \U$37216 ( \37559 , \37557 , \37558 );
not \U$37217 ( \37560 , \3918 );
and \U$37218 ( \37561 , \3683 , RI986e008_8);
and \U$37219 ( \37562 , RI986df18_6, \3681 );
nor \U$37220 ( \37563 , \37561 , \37562 );
not \U$37221 ( \37564 , \37563 );
or \U$37222 ( \37565 , \37560 , \37564 );
or \U$37223 ( \37566 , \37563 , \3412 );
nand \U$37224 ( \37567 , \37565 , \37566 );
xor \U$37225 ( \37568 , \37559 , \37567 );
and \U$37226 ( \37569 , \4203 , RI986de28_4);
and \U$37227 ( \37570 , RI986dd38_2, \4201 );
nor \U$37228 ( \37571 , \37569 , \37570 );
and \U$37229 ( \37572 , \37571 , \4207 );
not \U$37230 ( \37573 , \37571 );
and \U$37231 ( \37574 , \37573 , \3922 );
nor \U$37232 ( \37575 , \37572 , \37574 );
xor \U$37233 ( \37576 , \37568 , \37575 );
not \U$37234 ( \37577 , \4519 );
and \U$37235 ( \37578 , \4710 , RI986e1e8_12);
and \U$37236 ( \37579 , RI986e0f8_10, \4708 );
nor \U$37237 ( \37580 , \37578 , \37579 );
not \U$37238 ( \37581 , \37580 );
or \U$37239 ( \37582 , \37577 , \37581 );
or \U$37240 ( \37583 , \37580 , \4521 );
nand \U$37241 ( \37584 , \37582 , \37583 );
xor \U$37242 ( \37585 , \37584 , \5594 );
and \U$37243 ( \37586 , \5318 , RI986e2d8_14);
and \U$37244 ( \37587 , RI986e3c8_16, \5316 );
nor \U$37245 ( \37588 , \37586 , \37587 );
and \U$37246 ( \37589 , \37588 , \5052 );
not \U$37247 ( \37590 , \37588 );
and \U$37248 ( \37591 , \37590 , \5322 );
nor \U$37249 ( \37592 , \37589 , \37591 );
xor \U$37250 ( \37593 , \37585 , \37592 );
not \U$37251 ( \37594 , \1462 );
and \U$37252 ( \37595 , \2042 , RI986f868_60);
and \U$37253 ( \37596 , RI986f778_58, \2040 );
nor \U$37254 ( \37597 , \37595 , \37596 );
not \U$37255 ( \37598 , \37597 );
or \U$37256 ( \37599 , \37594 , \37598 );
or \U$37257 ( \37600 , \37597 , \2034 );
nand \U$37258 ( \37601 , \37599 , \37600 );
and \U$37259 ( \37602 , \2274 , RI986fa48_64);
and \U$37260 ( \37603 , RI986f958_62, \2272 );
nor \U$37261 ( \37604 , \37602 , \37603 );
and \U$37262 ( \37605 , \37604 , \2030 );
not \U$37263 ( \37606 , \37604 );
and \U$37264 ( \37607 , \37606 , \2031 );
nor \U$37265 ( \37608 , \37605 , \37607 );
xor \U$37266 ( \37609 , \37601 , \37608 );
and \U$37267 ( \37610 , \2464 , RI986f4a8_52);
and \U$37268 ( \37611 , RI986f3b8_50, \2462 );
nor \U$37269 ( \37612 , \37610 , \37611 );
and \U$37270 ( \37613 , \37612 , \2468 );
not \U$37271 ( \37614 , \37612 );
and \U$37272 ( \37615 , \37614 , \2263 );
nor \U$37273 ( \37616 , \37613 , \37615 );
xor \U$37274 ( \37617 , \37609 , \37616 );
xor \U$37275 ( \37618 , \37593 , \37617 );
xor \U$37276 ( \37619 , \37576 , \37618 );
and \U$37277 ( \37620 , \37551 , \37619 );
and \U$37278 ( \37621 , \37502 , \37550 );
or \U$37279 ( \37622 , \37620 , \37621 );
and \U$37280 ( \37623 , \37468 , \37622 );
and \U$37281 ( \37624 , \37275 , \37467 );
or \U$37282 ( \37625 , \37623 , \37624 );
xor \U$37283 ( \37626 , \37601 , \37608 );
and \U$37284 ( \37627 , \37626 , \37616 );
and \U$37285 ( \37628 , \37601 , \37608 );
or \U$37286 ( \37629 , \37627 , \37628 );
xor \U$37287 ( \37630 , \37584 , \5594 );
and \U$37288 ( \37631 , \37630 , \37592 );
and \U$37289 ( \37632 , \37584 , \5594 );
or \U$37290 ( \37633 , \37631 , \37632 );
xor \U$37291 ( \37634 , \37629 , \37633 );
xor \U$37292 ( \37635 , \37559 , \37567 );
and \U$37293 ( \37636 , \37635 , \37575 );
and \U$37294 ( \37637 , \37559 , \37567 );
or \U$37295 ( \37638 , \37636 , \37637 );
xor \U$37296 ( \37639 , \37634 , \37638 );
xor \U$37297 ( \37640 , \37228 , \37235 );
and \U$37298 ( \37641 , \37640 , \37243 );
and \U$37299 ( \37642 , \37228 , \37235 );
or \U$37300 ( \37643 , \37641 , \37642 );
xor \U$37301 ( \37644 , \37202 , \37210 );
and \U$37302 ( \37645 , \37644 , \37219 );
and \U$37303 ( \37646 , \37202 , \37210 );
or \U$37304 ( \37647 , \37645 , \37646 );
xor \U$37305 ( \37648 , \37643 , \37647 );
xor \U$37306 ( \37649 , \37252 , \37259 );
and \U$37307 ( \37650 , \37649 , \37267 );
and \U$37308 ( \37651 , \37252 , \37259 );
or \U$37309 ( \37652 , \37650 , \37651 );
xor \U$37310 ( \37653 , \37648 , \37652 );
xor \U$37311 ( \37654 , \37639 , \37653 );
and \U$37312 ( \37655 , \395 , RI986ea58_30);
and \U$37313 ( \37656 , RI986e968_28, \393 );
nor \U$37314 ( \37657 , \37655 , \37656 );
not \U$37315 ( \37658 , \37657 );
not \U$37316 ( \37659 , \487 );
and \U$37317 ( \37660 , \37658 , \37659 );
and \U$37318 ( \37661 , \37657 , \487 );
nor \U$37319 ( \37662 , \37660 , \37661 );
and \U$37320 ( \37663 , \354 , RI9871668_124);
and \U$37321 ( \37664 , RI986eb48_32, \352 );
nor \U$37322 ( \37665 , \37663 , \37664 );
not \U$37323 ( \37666 , \37665 );
not \U$37324 ( \37667 , \345 );
and \U$37325 ( \37668 , \37666 , \37667 );
and \U$37326 ( \37669 , \37665 , \345 );
nor \U$37327 ( \37670 , \37668 , \37669 );
xor \U$37328 ( \37671 , \37662 , \37670 );
and \U$37329 ( \37672 , \416 , RI9871848_128);
and \U$37330 ( \37673 , RI9871578_122, \414 );
nor \U$37331 ( \37674 , \37672 , \37673 );
and \U$37332 ( \37675 , \37674 , \421 );
not \U$37333 ( \37676 , \37674 );
and \U$37334 ( \37677 , \37676 , \422 );
nor \U$37335 ( \37678 , \37675 , \37677 );
xor \U$37336 ( \37679 , \37671 , \37678 );
nand \U$37337 ( \37680 , RI9871758_126, RI9871fc8_144);
or \U$37338 ( \37681 , \37679 , \37680 );
nand \U$37339 ( \37682 , \37680 , \37679 );
nand \U$37340 ( \37683 , \37681 , \37682 );
and \U$37341 ( \37684 , \4203 , RI986dd38_2);
and \U$37342 ( \37685 , RI986e1e8_12, \4201 );
nor \U$37343 ( \37686 , \37684 , \37685 );
and \U$37344 ( \37687 , \37686 , \4207 );
not \U$37345 ( \37688 , \37686 );
and \U$37346 ( \37689 , \37688 , \3923 );
nor \U$37347 ( \37690 , \37687 , \37689 );
nand \U$37348 ( \37691 , RI986e3c8_16, \5318 );
and \U$37349 ( \37692 , \37691 , \5052 );
not \U$37350 ( \37693 , \37691 );
and \U$37351 ( \37694 , \37693 , \5322 );
nor \U$37352 ( \37695 , \37692 , \37694 );
xor \U$37353 ( \37696 , \37690 , \37695 );
not \U$37354 ( \37697 , \4519 );
and \U$37355 ( \37698 , \4710 , RI986e0f8_10);
and \U$37356 ( \37699 , RI986e2d8_14, \4708 );
nor \U$37357 ( \37700 , \37698 , \37699 );
not \U$37358 ( \37701 , \37700 );
or \U$37359 ( \37702 , \37697 , \37701 );
or \U$37360 ( \37703 , \37700 , \4521 );
nand \U$37361 ( \37704 , \37702 , \37703 );
xor \U$37362 ( \37705 , \37696 , \37704 );
xor \U$37363 ( \37706 , \37683 , \37705 );
and \U$37364 ( \37707 , \1311 , RI986e698_22);
and \U$37365 ( \37708 , RI986f868_60, \1309 );
nor \U$37366 ( \37709 , \37707 , \37708 );
and \U$37367 ( \37710 , \37709 , \1458 );
not \U$37368 ( \37711 , \37709 );
and \U$37369 ( \37712 , \37711 , \1315 );
nor \U$37370 ( \37713 , \37710 , \37712 );
not \U$37371 ( \37714 , \2034 );
and \U$37372 ( \37715 , \2042 , RI986f778_58);
and \U$37373 ( \37716 , RI986fa48_64, \2040 );
nor \U$37374 ( \37717 , \37715 , \37716 );
not \U$37375 ( \37718 , \37717 );
or \U$37376 ( \37719 , \37714 , \37718 );
or \U$37377 ( \37720 , \37717 , \2034 );
nand \U$37378 ( \37721 , \37719 , \37720 );
xor \U$37379 ( \37722 , \37713 , \37721 );
and \U$37380 ( \37723 , \2274 , RI986f958_62);
and \U$37381 ( \37724 , RI986f4a8_52, \2272 );
nor \U$37382 ( \37725 , \37723 , \37724 );
and \U$37383 ( \37726 , \37725 , \2030 );
not \U$37384 ( \37727 , \37725 );
and \U$37385 ( \37728 , \37727 , \2031 );
nor \U$37386 ( \37729 , \37726 , \37728 );
xor \U$37387 ( \37730 , \37722 , \37729 );
not \U$37388 ( \37731 , \456 );
and \U$37389 ( \37732 , \465 , RI986ee18_38);
and \U$37390 ( \37733 , RI986ec38_34, \463 );
nor \U$37391 ( \37734 , \37732 , \37733 );
not \U$37392 ( \37735 , \37734 );
or \U$37393 ( \37736 , \37731 , \37735 );
or \U$37394 ( \37737 , \37734 , \456 );
nand \U$37395 ( \37738 , \37736 , \37737 );
and \U$37396 ( \37739 , \438 , RI986ed28_36);
and \U$37397 ( \37740 , RI986f0e8_44, \436 );
nor \U$37398 ( \37741 , \37739 , \37740 );
and \U$37399 ( \37742 , \37741 , \444 );
not \U$37400 ( \37743 , \37741 );
and \U$37401 ( \37744 , \37743 , \443 );
nor \U$37402 ( \37745 , \37742 , \37744 );
xor \U$37403 ( \37746 , \37738 , \37745 );
not \U$37404 ( \37747 , \367 );
and \U$37405 ( \37748 , \376 , RI986e878_26);
and \U$37406 ( \37749 , RI986ef08_40, \374 );
nor \U$37407 ( \37750 , \37748 , \37749 );
not \U$37408 ( \37751 , \37750 );
or \U$37409 ( \37752 , \37747 , \37751 );
or \U$37410 ( \37753 , \37750 , \365 );
nand \U$37411 ( \37754 , \37752 , \37753 );
xor \U$37412 ( \37755 , \37746 , \37754 );
and \U$37413 ( \37756 , \776 , RI986eff8_42);
and \U$37414 ( \37757 , RI986f2c8_48, \774 );
nor \U$37415 ( \37758 , \37756 , \37757 );
and \U$37416 ( \37759 , \37758 , \474 );
not \U$37417 ( \37760 , \37758 );
and \U$37418 ( \37761 , \37760 , \451 );
nor \U$37419 ( \37762 , \37759 , \37761 );
not \U$37420 ( \37763 , \1301 );
and \U$37421 ( \37764 , \1293 , RI986f1d8_46);
and \U$37422 ( \37765 , RI986e5a8_20, \1291 );
nor \U$37423 ( \37766 , \37764 , \37765 );
not \U$37424 ( \37767 , \37766 );
or \U$37425 ( \37768 , \37763 , \37767 );
or \U$37426 ( \37769 , \37766 , \1301 );
nand \U$37427 ( \37770 , \37768 , \37769 );
xor \U$37428 ( \37771 , \37762 , \37770 );
and \U$37429 ( \37772 , \1329 , RI986e4b8_18);
and \U$37430 ( \37773 , RI986e788_24, \1327 );
nor \U$37431 ( \37774 , \37772 , \37773 );
and \U$37432 ( \37775 , \37774 , \1336 );
not \U$37433 ( \37776 , \37774 );
and \U$37434 ( \37777 , \37776 , \1337 );
nor \U$37435 ( \37778 , \37775 , \37777 );
xor \U$37436 ( \37779 , \37771 , \37778 );
xor \U$37437 ( \37780 , \37755 , \37779 );
xor \U$37438 ( \37781 , \37730 , \37780 );
xor \U$37439 ( \37782 , \37706 , \37781 );
and \U$37440 ( \37783 , \37654 , \37782 );
and \U$37441 ( \37784 , \37639 , \37653 );
or \U$37442 ( \37785 , \37783 , \37784 );
xor \U$37443 ( \37786 , \37625 , \37785 );
xor \U$37444 ( \37787 , \37713 , \37721 );
xor \U$37445 ( \37788 , \37787 , \37729 );
and \U$37446 ( \37789 , \37755 , \37788 );
xor \U$37447 ( \37790 , \37713 , \37721 );
xor \U$37448 ( \37791 , \37790 , \37729 );
and \U$37449 ( \37792 , \37779 , \37791 );
and \U$37450 ( \37793 , \37755 , \37779 );
or \U$37451 ( \37794 , \37789 , \37792 , \37793 );
xor \U$37452 ( \37795 , \36969 , \5052 );
xor \U$37453 ( \37796 , \37795 , \36978 );
xor \U$37454 ( \37797 , \37794 , \37796 );
xor \U$37455 ( \37798 , \36943 , \36950 );
xor \U$37456 ( \37799 , \37798 , \36959 );
xor \U$37457 ( \37800 , \36892 , \36899 );
xor \U$37458 ( \37801 , \37800 , \36908 );
xor \U$37459 ( \37802 , \36989 , \36997 );
xor \U$37460 ( \37803 , \37802 , \37006 );
xor \U$37461 ( \37804 , \37801 , \37803 );
xor \U$37462 ( \37805 , \37799 , \37804 );
xor \U$37463 ( \37806 , \37797 , \37805 );
xor \U$37464 ( \37807 , \37629 , \37633 );
and \U$37465 ( \37808 , \37807 , \37638 );
and \U$37466 ( \37809 , \37629 , \37633 );
or \U$37467 ( \37810 , \37808 , \37809 );
xor \U$37468 ( \37811 , \37810 , \37682 );
xor \U$37469 ( \37812 , \37643 , \37647 );
and \U$37470 ( \37813 , \37812 , \37652 );
and \U$37471 ( \37814 , \37643 , \37647 );
or \U$37472 ( \37815 , \37813 , \37814 );
xor \U$37473 ( \37816 , \37811 , \37815 );
xor \U$37474 ( \37817 , \37738 , \37745 );
and \U$37475 ( \37818 , \37817 , \37754 );
and \U$37476 ( \37819 , \37738 , \37745 );
or \U$37477 ( \37820 , \37818 , \37819 );
xor \U$37478 ( \37821 , \37662 , \37670 );
and \U$37479 ( \37822 , \37821 , \37678 );
and \U$37480 ( \37823 , \37662 , \37670 );
nor \U$37481 ( \37824 , \37822 , \37823 );
xor \U$37482 ( \37825 , \37820 , \37824 );
xor \U$37483 ( \37826 , \37762 , \37770 );
and \U$37484 ( \37827 , \37826 , \37778 );
and \U$37485 ( \37828 , \37762 , \37770 );
or \U$37486 ( \37829 , \37827 , \37828 );
xor \U$37487 ( \37830 , \37825 , \37829 );
and \U$37488 ( \37831 , \2464 , RI986f3b8_50);
and \U$37489 ( \37832 , RI986f598_54, \2462 );
nor \U$37490 ( \37833 , \37831 , \37832 );
and \U$37491 ( \37834 , \37833 , \2468 );
not \U$37492 ( \37835 , \37833 );
and \U$37493 ( \37836 , \37835 , \2263 );
nor \U$37494 ( \37837 , \37834 , \37836 );
not \U$37495 ( \37838 , \3406 );
and \U$37496 ( \37839 , \3254 , RI986f688_56);
and \U$37497 ( \37840 , RI986e008_8, \3252 );
nor \U$37498 ( \37841 , \37839 , \37840 );
not \U$37499 ( \37842 , \37841 );
or \U$37500 ( \37843 , \37838 , \37842 );
or \U$37501 ( \37844 , \37841 , \2935 );
nand \U$37502 ( \37845 , \37843 , \37844 );
xor \U$37503 ( \37846 , \37837 , \37845 );
not \U$37504 ( \37847 , \3412 );
and \U$37505 ( \37848 , \3683 , RI986df18_6);
and \U$37506 ( \37849 , RI986de28_4, \3681 );
nor \U$37507 ( \37850 , \37848 , \37849 );
not \U$37508 ( \37851 , \37850 );
or \U$37509 ( \37852 , \37847 , \37851 );
or \U$37510 ( \37853 , \37850 , \3918 );
nand \U$37511 ( \37854 , \37852 , \37853 );
and \U$37512 ( \37855 , \37846 , \37854 );
and \U$37513 ( \37856 , \37837 , \37845 );
or \U$37514 ( \37857 , \37855 , \37856 );
xor \U$37515 ( \37858 , \37690 , \37695 );
and \U$37516 ( \37859 , \37858 , \37704 );
and \U$37517 ( \37860 , \37690 , \37695 );
or \U$37518 ( \37861 , \37859 , \37860 );
xor \U$37519 ( \37862 , \37857 , \37861 );
xor \U$37520 ( \37863 , \37713 , \37721 );
and \U$37521 ( \37864 , \37863 , \37729 );
and \U$37522 ( \37865 , \37713 , \37721 );
or \U$37523 ( \37866 , \37864 , \37865 );
xor \U$37524 ( \37867 , \37862 , \37866 );
xor \U$37525 ( \37868 , \36865 , \36873 );
xor \U$37526 ( \37869 , \37868 , \36881 );
not \U$37527 ( \37870 , RI9871848_128);
nor \U$37528 ( \37871 , \37870 , \407 );
xor \U$37529 ( \37872 , \36838 , \36845 );
xor \U$37530 ( \37873 , \37872 , \36854 );
xor \U$37531 ( \37874 , \37871 , \37873 );
xor \U$37532 ( \37875 , \37869 , \37874 );
xor \U$37533 ( \37876 , \37867 , \37875 );
xor \U$37534 ( \37877 , \37830 , \37876 );
xor \U$37535 ( \37878 , \37816 , \37877 );
xor \U$37536 ( \37879 , \37806 , \37878 );
and \U$37537 ( \37880 , \37786 , \37879 );
and \U$37538 ( \37881 , \37625 , \37785 );
or \U$37539 ( \37882 , \37880 , \37881 );
xor \U$37540 ( \37883 , \37820 , \37824 );
xor \U$37541 ( \37884 , \37883 , \37829 );
and \U$37542 ( \37885 , \37867 , \37884 );
xor \U$37543 ( \37886 , \37820 , \37824 );
xor \U$37544 ( \37887 , \37886 , \37829 );
and \U$37545 ( \37888 , \37875 , \37887 );
and \U$37546 ( \37889 , \37867 , \37875 );
or \U$37547 ( \37890 , \37885 , \37888 , \37889 );
xor \U$37548 ( \37891 , \37810 , \37682 );
and \U$37549 ( \37892 , \37891 , \37815 );
and \U$37550 ( \37893 , \37810 , \37682 );
or \U$37551 ( \37894 , \37892 , \37893 );
xor \U$37552 ( \37895 , \37890 , \37894 );
xor \U$37553 ( \37896 , \37794 , \37796 );
and \U$37554 ( \37897 , \37896 , \37805 );
and \U$37555 ( \37898 , \37794 , \37796 );
or \U$37556 ( \37899 , \37897 , \37898 );
xor \U$37557 ( \37900 , \37895 , \37899 );
xor \U$37558 ( \37901 , \37882 , \37900 );
xor \U$37559 ( \37902 , \37794 , \37796 );
xor \U$37560 ( \37903 , \37902 , \37805 );
and \U$37561 ( \37904 , \37816 , \37903 );
xor \U$37562 ( \37905 , \37794 , \37796 );
xor \U$37563 ( \37906 , \37905 , \37805 );
and \U$37564 ( \37907 , \37877 , \37906 );
and \U$37565 ( \37908 , \37816 , \37877 );
or \U$37566 ( \37909 , \37904 , \37907 , \37908 );
xor \U$37567 ( \37910 , \37559 , \37567 );
xor \U$37568 ( \37911 , \37910 , \37575 );
and \U$37569 ( \37912 , \37593 , \37911 );
xor \U$37570 ( \37913 , \37559 , \37567 );
xor \U$37571 ( \37914 , \37913 , \37575 );
and \U$37572 ( \37915 , \37617 , \37914 );
and \U$37573 ( \37916 , \37593 , \37617 );
or \U$37574 ( \37917 , \37912 , \37915 , \37916 );
xor \U$37575 ( \37918 , \37837 , \37845 );
xor \U$37576 ( \37919 , \37918 , \37854 );
xor \U$37577 ( \37920 , \37917 , \37919 );
xor \U$37578 ( \37921 , \37202 , \37210 );
xor \U$37579 ( \37922 , \37921 , \37219 );
and \U$37580 ( \37923 , \37244 , \37922 );
xor \U$37581 ( \37924 , \37202 , \37210 );
xor \U$37582 ( \37925 , \37924 , \37219 );
and \U$37583 ( \37926 , \37268 , \37925 );
and \U$37584 ( \37927 , \37244 , \37268 );
or \U$37585 ( \37928 , \37923 , \37926 , \37927 );
and \U$37586 ( \37929 , \37920 , \37928 );
and \U$37587 ( \37930 , \37917 , \37919 );
or \U$37588 ( \37931 , \37929 , \37930 );
xor \U$37589 ( \37932 , \37481 , \37488 );
and \U$37590 ( \37933 , \37932 , \37496 );
and \U$37591 ( \37934 , \37481 , \37488 );
or \U$37592 ( \37935 , \37933 , \37934 );
xor \U$37593 ( \37936 , \37535 , \37540 );
and \U$37594 ( \37937 , \37936 , \37548 );
and \U$37595 ( \37938 , \37535 , \37540 );
or \U$37596 ( \37939 , \37937 , \37938 );
xor \U$37597 ( \37940 , \37935 , \37939 );
xor \U$37598 ( \37941 , \37510 , \37518 );
and \U$37599 ( \37942 , \37941 , \37526 );
and \U$37600 ( \37943 , \37510 , \37518 );
or \U$37601 ( \37944 , \37942 , \37943 );
and \U$37602 ( \37945 , \37940 , \37944 );
and \U$37603 ( \37946 , \37935 , \37939 );
or \U$37604 ( \37947 , \37945 , \37946 );
xor \U$37605 ( \37948 , \37098 , \37100 );
and \U$37606 ( \37949 , \37948 , \37110 );
and \U$37607 ( \37950 , \37098 , \37100 );
or \U$37608 ( \37951 , \37949 , \37950 );
xor \U$37609 ( \37952 , \37947 , \37951 );
xor \U$37610 ( \37953 , \37137 , \37165 );
and \U$37611 ( \37954 , \37953 , \37192 );
and \U$37612 ( \37955 , \37137 , \37165 );
or \U$37613 ( \37956 , \37954 , \37955 );
and \U$37614 ( \37957 , \37952 , \37956 );
and \U$37615 ( \37958 , \37947 , \37951 );
or \U$37616 ( \37959 , \37957 , \37958 );
xor \U$37617 ( \37960 , \37931 , \37959 );
xor \U$37618 ( \37961 , \37683 , \37705 );
and \U$37619 ( \37962 , \37961 , \37781 );
and \U$37620 ( \37963 , \37683 , \37705 );
or \U$37621 ( \37964 , \37962 , \37963 );
and \U$37622 ( \37965 , \37960 , \37964 );
and \U$37623 ( \37966 , \37931 , \37959 );
or \U$37624 ( \37967 , \37965 , \37966 );
xor \U$37625 ( \37968 , \37909 , \37967 );
xor \U$37626 ( \37969 , \36943 , \36950 );
xor \U$37627 ( \37970 , \37969 , \36959 );
and \U$37628 ( \37971 , \37801 , \37970 );
xor \U$37629 ( \37972 , \36943 , \36950 );
xor \U$37630 ( \37973 , \37972 , \36959 );
and \U$37631 ( \37974 , \37803 , \37973 );
and \U$37632 ( \37975 , \37801 , \37803 );
or \U$37633 ( \37976 , \37971 , \37974 , \37975 );
xor \U$37634 ( \37977 , \36566 , \36572 );
xor \U$37635 ( \37978 , \37977 , \36580 );
xor \U$37636 ( \37979 , \37976 , \37978 );
xor \U$37637 ( \37980 , \36673 , \36680 );
xor \U$37638 ( \37981 , \37980 , \36689 );
xor \U$37639 ( \37982 , \37033 , \37038 );
xor \U$37640 ( \37983 , \37981 , \37982 );
xor \U$37641 ( \37984 , \37979 , \37983 );
xor \U$37642 ( \37985 , \37857 , \37861 );
and \U$37643 ( \37986 , \37985 , \37866 );
and \U$37644 ( \37987 , \37857 , \37861 );
or \U$37645 ( \37988 , \37986 , \37987 );
xor \U$37646 ( \37989 , \37820 , \37824 );
and \U$37647 ( \37990 , \37989 , \37829 );
and \U$37648 ( \37991 , \37820 , \37824 );
or \U$37649 ( \37992 , \37990 , \37991 );
xor \U$37650 ( \37993 , \37988 , \37992 );
xor \U$37651 ( \37994 , \36865 , \36873 );
xor \U$37652 ( \37995 , \37994 , \36881 );
and \U$37653 ( \37996 , \37871 , \37995 );
xor \U$37654 ( \37997 , \36865 , \36873 );
xor \U$37655 ( \37998 , \37997 , \36881 );
and \U$37656 ( \37999 , \37873 , \37998 );
and \U$37657 ( \38000 , \37871 , \37873 );
or \U$37658 ( \38001 , \37996 , \37999 , \38000 );
xor \U$37659 ( \38002 , \37993 , \38001 );
xor \U$37660 ( \38003 , \36962 , \36981 );
xor \U$37661 ( \38004 , \38003 , \37009 );
or \U$37662 ( \38005 , \36924 , \36934 );
nand \U$37663 ( \38006 , \38005 , \36935 );
xor \U$37664 ( \38007 , \36857 , \36884 );
xor \U$37665 ( \38008 , \38007 , \36911 );
xor \U$37666 ( \38009 , \38006 , \38008 );
xor \U$37667 ( \38010 , \38004 , \38009 );
xor \U$37668 ( \38011 , \38002 , \38010 );
xor \U$37669 ( \38012 , \37984 , \38011 );
xor \U$37670 ( \38013 , \37968 , \38012 );
and \U$37671 ( \38014 , \37901 , \38013 );
and \U$37672 ( \38015 , \37882 , \37900 );
or \U$37673 ( \38016 , \38014 , \38015 );
xor \U$37674 ( \38017 , \37909 , \37967 );
and \U$37675 ( \38018 , \38017 , \38012 );
and \U$37676 ( \38019 , \37909 , \37967 );
or \U$37677 ( \38020 , \38018 , \38019 );
xor \U$37678 ( \38021 , \36962 , \36981 );
xor \U$37679 ( \38022 , \38021 , \37009 );
and \U$37680 ( \38023 , \38006 , \38022 );
xor \U$37681 ( \38024 , \36962 , \36981 );
xor \U$37682 ( \38025 , \38024 , \37009 );
and \U$37683 ( \38026 , \38008 , \38025 );
and \U$37684 ( \38027 , \38006 , \38008 );
or \U$37685 ( \38028 , \38023 , \38026 , \38027 );
xor \U$37686 ( \38029 , \37988 , \37992 );
and \U$37687 ( \38030 , \38029 , \38001 );
and \U$37688 ( \38031 , \37988 , \37992 );
or \U$37689 ( \38032 , \38030 , \38031 );
xor \U$37690 ( \38033 , \38028 , \38032 );
xor \U$37691 ( \38034 , \37976 , \37978 );
and \U$37692 ( \38035 , \38034 , \37983 );
and \U$37693 ( \38036 , \37976 , \37978 );
or \U$37694 ( \38037 , \38035 , \38036 );
xor \U$37695 ( \38038 , \38033 , \38037 );
xor \U$37696 ( \38039 , \38020 , \38038 );
xor \U$37697 ( \38040 , \37976 , \37978 );
xor \U$37698 ( \38041 , \38040 , \37983 );
and \U$37699 ( \38042 , \38002 , \38041 );
xor \U$37700 ( \38043 , \37976 , \37978 );
xor \U$37701 ( \38044 , \38043 , \37983 );
and \U$37702 ( \38045 , \38010 , \38044 );
and \U$37703 ( \38046 , \38002 , \38010 );
or \U$37704 ( \38047 , \38042 , \38045 , \38046 );
xor \U$37705 ( \38048 , \37890 , \37894 );
and \U$37706 ( \38049 , \38048 , \37899 );
and \U$37707 ( \38050 , \37890 , \37894 );
or \U$37708 ( \38051 , \38049 , \38050 );
xor \U$37709 ( \38052 , \38047 , \38051 );
xor \U$37710 ( \38053 , \36914 , \36935 );
xor \U$37711 ( \38054 , \38053 , \37012 );
xor \U$37712 ( \38055 , \37017 , \37019 );
xor \U$37713 ( \38056 , \37031 , \37043 );
xor \U$37714 ( \38057 , \38056 , \37050 );
xor \U$37715 ( \38058 , \38055 , \38057 );
xor \U$37716 ( \38059 , \38054 , \38058 );
xor \U$37717 ( \38060 , \38052 , \38059 );
xor \U$37718 ( \38061 , \38039 , \38060 );
xor \U$37719 ( \38062 , \38016 , \38061 );
not \U$37720 ( \38063 , \38062 );
xor \U$37721 ( \38064 , \37931 , \37959 );
xor \U$37722 ( \38065 , \38064 , \37964 );
xor \U$37723 ( \38066 , \37947 , \37951 );
xor \U$37724 ( \38067 , \38066 , \37956 );
xor \U$37725 ( \38068 , \37639 , \37653 );
xor \U$37726 ( \38069 , \38068 , \37782 );
and \U$37727 ( \38070 , \38067 , \38069 );
xor \U$37728 ( \38071 , \37275 , \37467 );
xor \U$37729 ( \38072 , \38071 , \37622 );
xor \U$37730 ( \38073 , \37639 , \37653 );
xor \U$37731 ( \38074 , \38073 , \37782 );
and \U$37732 ( \38075 , \38072 , \38074 );
and \U$37733 ( \38076 , \38067 , \38072 );
or \U$37734 ( \38077 , \38070 , \38075 , \38076 );
xor \U$37735 ( \38078 , \38065 , \38077 );
xor \U$37736 ( \38079 , \37386 , \37404 );
xor \U$37737 ( \38080 , \38079 , \37431 );
xor \U$37738 ( \38081 , \37301 , \37329 );
xor \U$37739 ( \38082 , \38081 , \37356 );
xor \U$37740 ( \38083 , \38080 , \38082 );
xor \U$37741 ( \38084 , \37456 , \37458 );
xor \U$37742 ( \38085 , \38084 , \37461 );
and \U$37743 ( \38086 , \38083 , \38085 );
and \U$37744 ( \38087 , \38080 , \38082 );
or \U$37745 ( \38088 , \38086 , \38087 );
not \U$37746 ( \38089 , \3918 );
and \U$37747 ( \38090 , \3683 , RI986f3b8_50);
and \U$37748 ( \38091 , RI986f598_54, \3681 );
nor \U$37749 ( \38092 , \38090 , \38091 );
not \U$37750 ( \38093 , \38092 );
or \U$37751 ( \38094 , \38089 , \38093 );
or \U$37752 ( \38095 , \38092 , \3918 );
nand \U$37753 ( \38096 , \38094 , \38095 );
and \U$37754 ( \38097 , \4203 , RI986f688_56);
and \U$37755 ( \38098 , RI986e008_8, \4201 );
nor \U$37756 ( \38099 , \38097 , \38098 );
and \U$37757 ( \38100 , \38099 , \4207 );
not \U$37758 ( \38101 , \38099 );
and \U$37759 ( \38102 , \38101 , \3923 );
nor \U$37760 ( \38103 , \38100 , \38102 );
xor \U$37761 ( \38104 , \38096 , \38103 );
not \U$37762 ( \38105 , \4519 );
and \U$37763 ( \38106 , \4710 , RI986df18_6);
and \U$37764 ( \38107 , RI986de28_4, \4708 );
nor \U$37765 ( \38108 , \38106 , \38107 );
not \U$37766 ( \38109 , \38108 );
or \U$37767 ( \38110 , \38105 , \38109 );
or \U$37768 ( \38111 , \38108 , \4519 );
nand \U$37769 ( \38112 , \38110 , \38111 );
and \U$37770 ( \38113 , \38104 , \38112 );
and \U$37771 ( \38114 , \38096 , \38103 );
or \U$37772 ( \38115 , \38113 , \38114 );
and \U$37773 ( \38116 , \5318 , RI986dd38_2);
and \U$37774 ( \38117 , RI986e1e8_12, \5316 );
nor \U$37775 ( \38118 , \38116 , \38117 );
and \U$37776 ( \38119 , \38118 , \5052 );
not \U$37777 ( \38120 , \38118 );
and \U$37778 ( \38121 , \38120 , \5322 );
nor \U$37779 ( \38122 , \38119 , \38121 );
nand \U$37780 ( \38123 , RI986e3c8_16, \6453 );
and \U$37781 ( \38124 , \38123 , \6190 );
not \U$37782 ( \38125 , \38123 );
and \U$37783 ( \38126 , \38125 , \6705 );
nor \U$37784 ( \38127 , \38124 , \38126 );
xor \U$37785 ( \38128 , \38122 , \38127 );
and \U$37786 ( \38129 , \5881 , RI986e0f8_10);
and \U$37787 ( \38130 , RI986e2d8_14, \5879 );
nor \U$37788 ( \38131 , \38129 , \38130 );
and \U$37789 ( \38132 , \38131 , \5594 );
not \U$37790 ( \38133 , \38131 );
and \U$37791 ( \38134 , \38133 , \5885 );
nor \U$37792 ( \38135 , \38132 , \38134 );
and \U$37793 ( \38136 , \38128 , \38135 );
and \U$37794 ( \38137 , \38122 , \38127 );
or \U$37795 ( \38138 , \38136 , \38137 );
xor \U$37796 ( \38139 , \38115 , \38138 );
not \U$37797 ( \38140 , \3406 );
and \U$37798 ( \38141 , \3254 , RI986f958_62);
and \U$37799 ( \38142 , RI986f4a8_52, \3252 );
nor \U$37800 ( \38143 , \38141 , \38142 );
not \U$37801 ( \38144 , \38143 );
or \U$37802 ( \38145 , \38140 , \38144 );
or \U$37803 ( \38146 , \38143 , \3406 );
nand \U$37804 ( \38147 , \38145 , \38146 );
and \U$37805 ( \38148 , \2274 , RI986e698_22);
and \U$37806 ( \38149 , RI986f868_60, \2272 );
nor \U$37807 ( \38150 , \38148 , \38149 );
and \U$37808 ( \38151 , \38150 , \2030 );
not \U$37809 ( \38152 , \38150 );
and \U$37810 ( \38153 , \38152 , \2031 );
nor \U$37811 ( \38154 , \38151 , \38153 );
xor \U$37812 ( \38155 , \38147 , \38154 );
and \U$37813 ( \38156 , \2464 , RI986f778_58);
and \U$37814 ( \38157 , RI986fa48_64, \2462 );
nor \U$37815 ( \38158 , \38156 , \38157 );
and \U$37816 ( \38159 , \38158 , \2468 );
not \U$37817 ( \38160 , \38158 );
and \U$37818 ( \38161 , \38160 , \2263 );
nor \U$37819 ( \38162 , \38159 , \38161 );
and \U$37820 ( \38163 , \38155 , \38162 );
and \U$37821 ( \38164 , \38147 , \38154 );
or \U$37822 ( \38165 , \38163 , \38164 );
and \U$37823 ( \38166 , \38139 , \38165 );
and \U$37824 ( \38167 , \38115 , \38138 );
or \U$37825 ( \38168 , \38166 , \38167 );
and \U$37826 ( \38169 , \438 , RI986e878_26);
and \U$37827 ( \38170 , RI986ef08_40, \436 );
nor \U$37828 ( \38171 , \38169 , \38170 );
and \U$37829 ( \38172 , \38171 , \444 );
not \U$37830 ( \38173 , \38171 );
and \U$37831 ( \38174 , \38173 , \443 );
nor \U$37832 ( \38175 , \38172 , \38174 );
and \U$37833 ( \38176 , \776 , RI986ee18_38);
and \U$37834 ( \38177 , RI986ec38_34, \774 );
nor \U$37835 ( \38178 , \38176 , \38177 );
and \U$37836 ( \38179 , \38178 , \474 );
not \U$37837 ( \38180 , \38178 );
and \U$37838 ( \38181 , \38180 , \451 );
nor \U$37839 ( \38182 , \38179 , \38181 );
xor \U$37840 ( \38183 , \38175 , \38182 );
not \U$37841 ( \38184 , \1128 );
and \U$37842 ( \38185 , \1293 , RI986ed28_36);
and \U$37843 ( \38186 , RI986f0e8_44, \1291 );
nor \U$37844 ( \38187 , \38185 , \38186 );
not \U$37845 ( \38188 , \38187 );
or \U$37846 ( \38189 , \38184 , \38188 );
or \U$37847 ( \38190 , \38187 , \1301 );
nand \U$37848 ( \38191 , \38189 , \38190 );
and \U$37849 ( \38192 , \38183 , \38191 );
and \U$37850 ( \38193 , \38175 , \38182 );
or \U$37851 ( \38194 , \38192 , \38193 );
not \U$37852 ( \38195 , \365 );
and \U$37853 ( \38196 , \376 , RI9871668_124);
and \U$37854 ( \38197 , RI986eb48_32, \374 );
nor \U$37855 ( \38198 , \38196 , \38197 );
not \U$37856 ( \38199 , \38198 );
or \U$37857 ( \38200 , \38195 , \38199 );
or \U$37858 ( \38201 , \38198 , \367 );
nand \U$37859 ( \38202 , \38200 , \38201 );
not \U$37860 ( \38203 , \454 );
and \U$37861 ( \38204 , \465 , RI986ea58_30);
and \U$37862 ( \38205 , RI986e968_28, \463 );
nor \U$37863 ( \38206 , \38204 , \38205 );
not \U$37864 ( \38207 , \38206 );
or \U$37865 ( \38208 , \38203 , \38207 );
or \U$37866 ( \38209 , \38206 , \454 );
nand \U$37867 ( \38210 , \38208 , \38209 );
xor \U$37868 ( \38211 , \38202 , \38210 );
not \U$37869 ( \38212 , \386 );
and \U$37870 ( \38213 , \395 , RI9871848_128);
and \U$37871 ( \38214 , RI9871578_122, \393 );
nor \U$37872 ( \38215 , \38213 , \38214 );
not \U$37873 ( \38216 , \38215 );
or \U$37874 ( \38217 , \38212 , \38216 );
or \U$37875 ( \38218 , \38215 , \386 );
nand \U$37876 ( \38219 , \38217 , \38218 );
and \U$37877 ( \38220 , \38211 , \38219 );
and \U$37878 ( \38221 , \38202 , \38210 );
or \U$37879 ( \38222 , \38220 , \38221 );
xor \U$37880 ( \38223 , \38194 , \38222 );
and \U$37881 ( \38224 , \1329 , RI986eff8_42);
and \U$37882 ( \38225 , RI986f2c8_48, \1327 );
nor \U$37883 ( \38226 , \38224 , \38225 );
and \U$37884 ( \38227 , \38226 , \1336 );
not \U$37885 ( \38228 , \38226 );
and \U$37886 ( \38229 , \38228 , \1337 );
nor \U$37887 ( \38230 , \38227 , \38229 );
and \U$37888 ( \38231 , \1311 , RI986f1d8_46);
and \U$37889 ( \38232 , RI986e5a8_20, \1309 );
nor \U$37890 ( \38233 , \38231 , \38232 );
and \U$37891 ( \38234 , \38233 , \1458 );
not \U$37892 ( \38235 , \38233 );
and \U$37893 ( \38236 , \38235 , \1315 );
nor \U$37894 ( \38237 , \38234 , \38236 );
xor \U$37895 ( \38238 , \38230 , \38237 );
not \U$37896 ( \38239 , \1462 );
and \U$37897 ( \38240 , \2042 , RI986e4b8_18);
and \U$37898 ( \38241 , RI986e788_24, \2040 );
nor \U$37899 ( \38242 , \38240 , \38241 );
not \U$37900 ( \38243 , \38242 );
or \U$37901 ( \38244 , \38239 , \38243 );
or \U$37902 ( \38245 , \38242 , \2034 );
nand \U$37903 ( \38246 , \38244 , \38245 );
and \U$37904 ( \38247 , \38238 , \38246 );
and \U$37905 ( \38248 , \38230 , \38237 );
or \U$37906 ( \38249 , \38247 , \38248 );
and \U$37907 ( \38250 , \38223 , \38249 );
and \U$37908 ( \38251 , \38194 , \38222 );
or \U$37909 ( \38252 , \38250 , \38251 );
xor \U$37910 ( \38253 , \38168 , \38252 );
xor \U$37911 ( \38254 , \37442 , \37444 );
xor \U$37912 ( \38255 , \38254 , \37453 );
and \U$37913 ( \38256 , \416 , RI98711b8_114);
and \U$37914 ( \38257 , RI9871398_118, \414 );
nor \U$37915 ( \38258 , \38256 , \38257 );
and \U$37916 ( \38259 , \38258 , \421 );
not \U$37917 ( \38260 , \38258 );
and \U$37918 ( \38261 , \38260 , \422 );
nor \U$37919 ( \38262 , \38259 , \38261 );
nand \U$37920 ( \38263 , RI98712a8_116, RI9871fc8_144);
or \U$37921 ( \38264 , \38262 , \38263 );
not \U$37922 ( \38265 , \38263 );
not \U$37923 ( \38266 , \38262 );
or \U$37924 ( \38267 , \38265 , \38266 );
not \U$37925 ( \38268 , \361 );
and \U$37926 ( \38269 , \354 , RI9871488_120);
and \U$37927 ( \38270 , RI9871758_126, \352 );
nor \U$37928 ( \38271 , \38269 , \38270 );
not \U$37929 ( \38272 , \38271 );
or \U$37930 ( \38273 , \38268 , \38272 );
or \U$37931 ( \38274 , \38271 , \345 );
nand \U$37932 ( \38275 , \38273 , \38274 );
nand \U$37933 ( \38276 , \38267 , \38275 );
nand \U$37934 ( \38277 , \38264 , \38276 );
xor \U$37935 ( \38278 , \38255 , \38277 );
xor \U$37936 ( \38279 , \37309 , \37317 );
xor \U$37937 ( \38280 , \38279 , \37326 );
and \U$37938 ( \38281 , \38278 , \38280 );
and \U$37939 ( \38282 , \38255 , \38277 );
or \U$37940 ( \38283 , \38281 , \38282 );
and \U$37941 ( \38284 , \38253 , \38283 );
and \U$37942 ( \38285 , \38168 , \38252 );
or \U$37943 ( \38286 , \38284 , \38285 );
xor \U$37944 ( \38287 , \38088 , \38286 );
xor \U$37945 ( \38288 , \37282 , \37289 );
xor \U$37946 ( \38289 , \38288 , \37298 );
xor \U$37947 ( \38290 , \37412 , \37419 );
xor \U$37948 ( \38291 , \38290 , \37428 );
and \U$37949 ( \38292 , \38289 , \38291 );
xor \U$37950 ( \38293 , \37337 , \37344 );
xor \U$37951 ( \38294 , \38293 , \37353 );
xor \U$37952 ( \38295 , \37412 , \37419 );
xor \U$37953 ( \38296 , \38295 , \37428 );
and \U$37954 ( \38297 , \38294 , \38296 );
and \U$37955 ( \38298 , \38289 , \38294 );
or \U$37956 ( \38299 , \38292 , \38297 , \38298 );
xor \U$37957 ( \38300 , \37527 , \37549 );
xor \U$37958 ( \38301 , \38299 , \38300 );
xor \U$37959 ( \38302 , \37119 , \37126 );
xor \U$37960 ( \38303 , \38302 , \37134 );
xor \U$37961 ( \38304 , \37470 , \37497 );
xor \U$37962 ( \38305 , \38303 , \38304 );
and \U$37963 ( \38306 , \38301 , \38305 );
and \U$37964 ( \38307 , \38299 , \38300 );
or \U$37965 ( \38308 , \38306 , \38307 );
and \U$37966 ( \38309 , \38287 , \38308 );
and \U$37967 ( \38310 , \38088 , \38286 );
or \U$37968 ( \38311 , \38309 , \38310 );
xor \U$37969 ( \38312 , \37917 , \37919 );
xor \U$37970 ( \38313 , \38312 , \37928 );
xor \U$37971 ( \38314 , \38311 , \38313 );
xor \U$37972 ( \38315 , \37935 , \37939 );
xor \U$37973 ( \38316 , \38315 , \37944 );
xor \U$37974 ( \38317 , \37502 , \37550 );
xor \U$37975 ( \38318 , \38317 , \37619 );
and \U$37976 ( \38319 , \38316 , \38318 );
xor \U$37977 ( \38320 , \37137 , \37165 );
xor \U$37978 ( \38321 , \38320 , \37192 );
xor \U$37979 ( \38322 , \37111 , \37270 );
xor \U$37980 ( \38323 , \38321 , \38322 );
xor \U$37981 ( \38324 , \37502 , \37550 );
xor \U$37982 ( \38325 , \38324 , \37619 );
and \U$37983 ( \38326 , \38323 , \38325 );
and \U$37984 ( \38327 , \38316 , \38323 );
or \U$37985 ( \38328 , \38319 , \38326 , \38327 );
and \U$37986 ( \38329 , \38314 , \38328 );
and \U$37987 ( \38330 , \38311 , \38313 );
or \U$37988 ( \38331 , \38329 , \38330 );
and \U$37989 ( \38332 , \38078 , \38331 );
and \U$37990 ( \38333 , \38065 , \38077 );
nor \U$37991 ( \38334 , \38332 , \38333 );
not \U$37992 ( \38335 , \38334 );
xor \U$37993 ( \38336 , \37882 , \37900 );
xor \U$37994 ( \38337 , \38336 , \38013 );
nand \U$37995 ( \38338 , \38335 , \38337 );
or \U$37996 ( \38339 , \38063 , \38338 );
not \U$37997 ( \38340 , \38062 );
not \U$37998 ( \38341 , \38338 );
and \U$37999 ( \38342 , \38340 , \38341 );
and \U$38000 ( \38343 , \38062 , \38338 );
nor \U$38001 ( \38344 , \38342 , \38343 );
xor \U$38002 ( \38345 , \38202 , \38210 );
xor \U$38003 ( \38346 , \38345 , \38219 );
xor \U$38004 ( \38347 , \38230 , \38237 );
xor \U$38005 ( \38348 , \38347 , \38246 );
and \U$38006 ( \38349 , \38346 , \38348 );
xor \U$38007 ( \38350 , \38175 , \38182 );
xor \U$38008 ( \38351 , \38350 , \38191 );
xor \U$38009 ( \38352 , \38230 , \38237 );
xor \U$38010 ( \38353 , \38352 , \38246 );
and \U$38011 ( \38354 , \38351 , \38353 );
and \U$38012 ( \38355 , \38346 , \38351 );
or \U$38013 ( \38356 , \38349 , \38354 , \38355 );
xor \U$38014 ( \38357 , \37367 , \37374 );
xor \U$38015 ( \38358 , \38357 , \37383 );
xor \U$38016 ( \38359 , \38356 , \38358 );
xor \U$38017 ( \38360 , \38122 , \38127 );
xor \U$38018 ( \38361 , \38360 , \38135 );
xor \U$38019 ( \38362 , \38096 , \38103 );
xor \U$38020 ( \38363 , \38362 , \38112 );
and \U$38021 ( \38364 , \38361 , \38363 );
xor \U$38022 ( \38365 , \38147 , \38154 );
xor \U$38023 ( \38366 , \38365 , \38162 );
xor \U$38024 ( \38367 , \38096 , \38103 );
xor \U$38025 ( \38368 , \38367 , \38112 );
and \U$38026 ( \38369 , \38366 , \38368 );
and \U$38027 ( \38370 , \38361 , \38366 );
or \U$38028 ( \38371 , \38364 , \38369 , \38370 );
and \U$38029 ( \38372 , \38359 , \38371 );
and \U$38030 ( \38373 , \38356 , \38358 );
or \U$38031 ( \38374 , \38372 , \38373 );
not \U$38032 ( \38375 , \3406 );
and \U$38033 ( \38376 , \3254 , RI986fa48_64);
and \U$38034 ( \38377 , RI986f958_62, \3252 );
nor \U$38035 ( \38378 , \38376 , \38377 );
not \U$38036 ( \38379 , \38378 );
or \U$38037 ( \38380 , \38375 , \38379 );
or \U$38038 ( \38381 , \38378 , \3406 );
nand \U$38039 ( \38382 , \38380 , \38381 );
and \U$38040 ( \38383 , \2464 , RI986f868_60);
and \U$38041 ( \38384 , RI986f778_58, \2462 );
nor \U$38042 ( \38385 , \38383 , \38384 );
and \U$38043 ( \38386 , \38385 , \2468 );
not \U$38044 ( \38387 , \38385 );
and \U$38045 ( \38388 , \38387 , \2263 );
nor \U$38046 ( \38389 , \38386 , \38388 );
xor \U$38047 ( \38390 , \38382 , \38389 );
not \U$38048 ( \38391 , \3412 );
and \U$38049 ( \38392 , \3683 , RI986f4a8_52);
and \U$38050 ( \38393 , RI986f3b8_50, \3681 );
nor \U$38051 ( \38394 , \38392 , \38393 );
not \U$38052 ( \38395 , \38394 );
or \U$38053 ( \38396 , \38391 , \38395 );
or \U$38054 ( \38397 , \38394 , \3412 );
nand \U$38055 ( \38398 , \38396 , \38397 );
and \U$38056 ( \38399 , \38390 , \38398 );
and \U$38057 ( \38400 , \38382 , \38389 );
or \U$38058 ( \38401 , \38399 , \38400 );
and \U$38059 ( \38402 , \5881 , RI986e1e8_12);
and \U$38060 ( \38403 , RI986e0f8_10, \5879 );
nor \U$38061 ( \38404 , \38402 , \38403 );
and \U$38062 ( \38405 , \38404 , \5594 );
not \U$38063 ( \38406 , \38404 );
and \U$38064 ( \38407 , \38406 , \5885 );
nor \U$38065 ( \38408 , \38405 , \38407 );
xor \U$38066 ( \38409 , \38408 , \6710 );
and \U$38067 ( \38410 , \6453 , RI986e2d8_14);
and \U$38068 ( \38411 , RI986e3c8_16, \6451 );
nor \U$38069 ( \38412 , \38410 , \38411 );
and \U$38070 ( \38413 , \38412 , \6190 );
not \U$38071 ( \38414 , \38412 );
and \U$38072 ( \38415 , \38414 , \6705 );
nor \U$38073 ( \38416 , \38413 , \38415 );
and \U$38074 ( \38417 , \38409 , \38416 );
and \U$38075 ( \38418 , \38408 , \6710 );
or \U$38076 ( \38419 , \38417 , \38418 );
xor \U$38077 ( \38420 , \38401 , \38419 );
and \U$38078 ( \38421 , \4203 , RI986f598_54);
and \U$38079 ( \38422 , RI986f688_56, \4201 );
nor \U$38080 ( \38423 , \38421 , \38422 );
and \U$38081 ( \38424 , \38423 , \4207 );
not \U$38082 ( \38425 , \38423 );
and \U$38083 ( \38426 , \38425 , \3923 );
nor \U$38084 ( \38427 , \38424 , \38426 );
not \U$38085 ( \38428 , \4521 );
and \U$38086 ( \38429 , \4710 , RI986e008_8);
and \U$38087 ( \38430 , RI986df18_6, \4708 );
nor \U$38088 ( \38431 , \38429 , \38430 );
not \U$38089 ( \38432 , \38431 );
or \U$38090 ( \38433 , \38428 , \38432 );
or \U$38091 ( \38434 , \38431 , \4519 );
nand \U$38092 ( \38435 , \38433 , \38434 );
xor \U$38093 ( \38436 , \38427 , \38435 );
and \U$38094 ( \38437 , \5318 , RI986de28_4);
and \U$38095 ( \38438 , RI986dd38_2, \5316 );
nor \U$38096 ( \38439 , \38437 , \38438 );
and \U$38097 ( \38440 , \38439 , \5052 );
not \U$38098 ( \38441 , \38439 );
and \U$38099 ( \38442 , \38441 , \5322 );
nor \U$38100 ( \38443 , \38440 , \38442 );
and \U$38101 ( \38444 , \38436 , \38443 );
and \U$38102 ( \38445 , \38427 , \38435 );
or \U$38103 ( \38446 , \38444 , \38445 );
and \U$38104 ( \38447 , \38420 , \38446 );
and \U$38105 ( \38448 , \38401 , \38419 );
or \U$38106 ( \38449 , \38447 , \38448 );
not \U$38107 ( \38450 , \386 );
and \U$38108 ( \38451 , \395 , RI9871758_126);
and \U$38109 ( \38452 , RI9871848_128, \393 );
nor \U$38110 ( \38453 , \38451 , \38452 );
not \U$38111 ( \38454 , \38453 );
or \U$38112 ( \38455 , \38450 , \38454 );
or \U$38113 ( \38456 , \38453 , \487 );
nand \U$38114 ( \38457 , \38455 , \38456 );
not \U$38115 ( \38458 , \361 );
and \U$38116 ( \38459 , \354 , RI9871398_118);
and \U$38117 ( \38460 , RI9871488_120, \352 );
nor \U$38118 ( \38461 , \38459 , \38460 );
not \U$38119 ( \38462 , \38461 );
or \U$38120 ( \38463 , \38458 , \38462 );
or \U$38121 ( \38464 , \38461 , \345 );
nand \U$38122 ( \38465 , \38463 , \38464 );
xor \U$38123 ( \38466 , \38457 , \38465 );
and \U$38124 ( \38467 , \416 , RI98712a8_116);
and \U$38125 ( \38468 , RI98711b8_114, \414 );
nor \U$38126 ( \38469 , \38467 , \38468 );
and \U$38127 ( \38470 , \38469 , \422 );
not \U$38128 ( \38471 , \38469 );
and \U$38129 ( \38472 , \38471 , \421 );
nor \U$38130 ( \38473 , \38470 , \38472 );
and \U$38131 ( \38474 , \38466 , \38473 );
and \U$38132 ( \38475 , \38457 , \38465 );
nor \U$38133 ( \38476 , \38474 , \38475 );
not \U$38134 ( \38477 , \38262 );
not \U$38135 ( \38478 , \38275 );
or \U$38136 ( \38479 , \38477 , \38478 );
or \U$38137 ( \38480 , \38262 , \38275 );
nand \U$38138 ( \38481 , \38479 , \38480 );
not \U$38139 ( \38482 , \38481 );
not \U$38140 ( \38483 , \38263 );
and \U$38141 ( \38484 , \38482 , \38483 );
and \U$38142 ( \38485 , \38481 , \38263 );
nor \U$38143 ( \38486 , \38484 , \38485 );
nand \U$38144 ( \38487 , \38476 , \38486 );
xor \U$38145 ( \38488 , \38449 , \38487 );
and \U$38146 ( \38489 , \2274 , RI986e788_24);
and \U$38147 ( \38490 , RI986e698_22, \2272 );
nor \U$38148 ( \38491 , \38489 , \38490 );
and \U$38149 ( \38492 , \38491 , \2030 );
not \U$38150 ( \38493 , \38491 );
and \U$38151 ( \38494 , \38493 , \2031 );
nor \U$38152 ( \38495 , \38492 , \38494 );
and \U$38153 ( \38496 , \1311 , RI986f2c8_48);
and \U$38154 ( \38497 , RI986f1d8_46, \1309 );
nor \U$38155 ( \38498 , \38496 , \38497 );
and \U$38156 ( \38499 , \38498 , \1319 );
not \U$38157 ( \38500 , \38498 );
and \U$38158 ( \38501 , \38500 , \1318 );
nor \U$38159 ( \38502 , \38499 , \38501 );
xor \U$38160 ( \38503 , \38495 , \38502 );
not \U$38161 ( \38504 , \1462 );
and \U$38162 ( \38505 , \2042 , RI986e5a8_20);
and \U$38163 ( \38506 , RI986e4b8_18, \2040 );
nor \U$38164 ( \38507 , \38505 , \38506 );
not \U$38165 ( \38508 , \38507 );
or \U$38166 ( \38509 , \38504 , \38508 );
or \U$38167 ( \38510 , \38507 , \2034 );
nand \U$38168 ( \38511 , \38509 , \38510 );
and \U$38169 ( \38512 , \38503 , \38511 );
and \U$38170 ( \38513 , \38495 , \38502 );
or \U$38171 ( \38514 , \38512 , \38513 );
not \U$38172 ( \38515 , \456 );
and \U$38173 ( \38516 , \465 , RI986eb48_32);
and \U$38174 ( \38517 , RI986ea58_30, \463 );
nor \U$38175 ( \38518 , \38516 , \38517 );
not \U$38176 ( \38519 , \38518 );
or \U$38177 ( \38520 , \38515 , \38519 );
or \U$38178 ( \38521 , \38518 , \456 );
nand \U$38179 ( \38522 , \38520 , \38521 );
and \U$38180 ( \38523 , \438 , RI986e968_28);
and \U$38181 ( \38524 , RI986e878_26, \436 );
nor \U$38182 ( \38525 , \38523 , \38524 );
and \U$38183 ( \38526 , \38525 , \444 );
not \U$38184 ( \38527 , \38525 );
and \U$38185 ( \38528 , \38527 , \443 );
nor \U$38186 ( \38529 , \38526 , \38528 );
xor \U$38187 ( \38530 , \38522 , \38529 );
not \U$38188 ( \38531 , \367 );
and \U$38189 ( \38532 , \376 , RI9871578_122);
and \U$38190 ( \38533 , RI9871668_124, \374 );
nor \U$38191 ( \38534 , \38532 , \38533 );
not \U$38192 ( \38535 , \38534 );
or \U$38193 ( \38536 , \38531 , \38535 );
or \U$38194 ( \38537 , \38534 , \367 );
nand \U$38195 ( \38538 , \38536 , \38537 );
and \U$38196 ( \38539 , \38530 , \38538 );
and \U$38197 ( \38540 , \38522 , \38529 );
or \U$38198 ( \38541 , \38539 , \38540 );
xor \U$38199 ( \38542 , \38514 , \38541 );
and \U$38200 ( \38543 , \1329 , RI986f0e8_44);
and \U$38201 ( \38544 , RI986eff8_42, \1327 );
nor \U$38202 ( \38545 , \38543 , \38544 );
and \U$38203 ( \38546 , \38545 , \1336 );
not \U$38204 ( \38547 , \38545 );
and \U$38205 ( \38548 , \38547 , \1337 );
nor \U$38206 ( \38549 , \38546 , \38548 );
and \U$38207 ( \38550 , \776 , RI986ef08_40);
and \U$38208 ( \38551 , RI986ee18_38, \774 );
nor \U$38209 ( \38552 , \38550 , \38551 );
and \U$38210 ( \38553 , \38552 , \474 );
not \U$38211 ( \38554 , \38552 );
and \U$38212 ( \38555 , \38554 , \451 );
nor \U$38213 ( \38556 , \38553 , \38555 );
xor \U$38214 ( \38557 , \38549 , \38556 );
not \U$38215 ( \38558 , \1301 );
and \U$38216 ( \38559 , \1293 , RI986ec38_34);
and \U$38217 ( \38560 , RI986ed28_36, \1291 );
nor \U$38218 ( \38561 , \38559 , \38560 );
not \U$38219 ( \38562 , \38561 );
or \U$38220 ( \38563 , \38558 , \38562 );
or \U$38221 ( \38564 , \38561 , \1301 );
nand \U$38222 ( \38565 , \38563 , \38564 );
and \U$38223 ( \38566 , \38557 , \38565 );
and \U$38224 ( \38567 , \38549 , \38556 );
or \U$38225 ( \38568 , \38566 , \38567 );
and \U$38226 ( \38569 , \38542 , \38568 );
and \U$38227 ( \38570 , \38514 , \38541 );
or \U$38228 ( \38571 , \38569 , \38570 );
and \U$38229 ( \38572 , \38488 , \38571 );
and \U$38230 ( \38573 , \38449 , \38487 );
or \U$38231 ( \38574 , \38572 , \38573 );
xor \U$38232 ( \38575 , \38374 , \38574 );
xor \U$38233 ( \38576 , \37393 , \6190 );
xor \U$38234 ( \38577 , \38576 , \37401 );
xor \U$38235 ( \38578 , \38255 , \38277 );
xor \U$38236 ( \38579 , \38578 , \38280 );
and \U$38237 ( \38580 , \38577 , \38579 );
xor \U$38238 ( \38581 , \37412 , \37419 );
xor \U$38239 ( \38582 , \38581 , \37428 );
xor \U$38240 ( \38583 , \38289 , \38294 );
xor \U$38241 ( \38584 , \38582 , \38583 );
xor \U$38242 ( \38585 , \38255 , \38277 );
xor \U$38243 ( \38586 , \38585 , \38280 );
and \U$38244 ( \38587 , \38584 , \38586 );
and \U$38245 ( \38588 , \38577 , \38584 );
or \U$38246 ( \38589 , \38580 , \38587 , \38588 );
and \U$38247 ( \38590 , \38575 , \38589 );
and \U$38248 ( \38591 , \38374 , \38574 );
or \U$38249 ( \38592 , \38590 , \38591 );
xor \U$38250 ( \38593 , \37359 , \37434 );
xor \U$38251 ( \38594 , \38593 , \37464 );
xor \U$38252 ( \38595 , \38592 , \38594 );
xor \U$38253 ( \38596 , \38168 , \38252 );
xor \U$38254 ( \38597 , \38596 , \38283 );
xor \U$38255 ( \38598 , \38080 , \38082 );
xor \U$38256 ( \38599 , \38598 , \38085 );
and \U$38257 ( \38600 , \38597 , \38599 );
xor \U$38258 ( \38601 , \38299 , \38300 );
xor \U$38259 ( \38602 , \38601 , \38305 );
xor \U$38260 ( \38603 , \38080 , \38082 );
xor \U$38261 ( \38604 , \38603 , \38085 );
and \U$38262 ( \38605 , \38602 , \38604 );
and \U$38263 ( \38606 , \38597 , \38602 );
or \U$38264 ( \38607 , \38600 , \38605 , \38606 );
and \U$38265 ( \38608 , \38595 , \38607 );
and \U$38266 ( \38609 , \38592 , \38594 );
or \U$38267 ( \38610 , \38608 , \38609 );
xor \U$38268 ( \38611 , \38088 , \38286 );
xor \U$38269 ( \38612 , \38611 , \38308 );
xor \U$38270 ( \38613 , \37502 , \37550 );
xor \U$38271 ( \38614 , \38613 , \37619 );
xor \U$38272 ( \38615 , \38316 , \38323 );
xor \U$38273 ( \38616 , \38614 , \38615 );
and \U$38274 ( \38617 , \38612 , \38616 );
xor \U$38275 ( \38618 , \38610 , \38617 );
xor \U$38276 ( \38619 , \37639 , \37653 );
xor \U$38277 ( \38620 , \38619 , \37782 );
xor \U$38278 ( \38621 , \38067 , \38072 );
xor \U$38279 ( \38622 , \38620 , \38621 );
and \U$38280 ( \38623 , \38618 , \38622 );
and \U$38281 ( \38624 , \38610 , \38617 );
or \U$38282 ( \38625 , \38623 , \38624 );
xor \U$38283 ( \38626 , \37625 , \37785 );
xor \U$38284 ( \38627 , \38626 , \37879 );
xor \U$38285 ( \38628 , \38625 , \38627 );
xor \U$38286 ( \38629 , \38065 , \38077 );
xor \U$38287 ( \38630 , \38629 , \38331 );
and \U$38288 ( \38631 , \38628 , \38630 );
and \U$38289 ( \38632 , \38625 , \38627 );
or \U$38290 ( \38633 , \38631 , \38632 );
not \U$38291 ( \38634 , \38334 );
not \U$38292 ( \38635 , \38337 );
or \U$38293 ( \38636 , \38634 , \38635 );
or \U$38294 ( \38637 , \38337 , \38334 );
nand \U$38295 ( \38638 , \38636 , \38637 );
and \U$38296 ( \38639 , \38633 , \38638 );
xor \U$38297 ( \38640 , \38638 , \38633 );
xor \U$38298 ( \38641 , \38449 , \38487 );
xor \U$38299 ( \38642 , \38641 , \38571 );
xor \U$38300 ( \38643 , \38194 , \38222 );
xor \U$38301 ( \38644 , \38643 , \38249 );
xor \U$38302 ( \38645 , \38115 , \38138 );
xor \U$38303 ( \38646 , \38645 , \38165 );
xor \U$38304 ( \38647 , \38644 , \38646 );
xor \U$38305 ( \38648 , \38255 , \38277 );
xor \U$38306 ( \38649 , \38648 , \38280 );
xor \U$38307 ( \38650 , \38577 , \38584 );
xor \U$38308 ( \38651 , \38649 , \38650 );
xor \U$38309 ( \38652 , \38647 , \38651 );
and \U$38310 ( \38653 , \38642 , \38652 );
or \U$38311 ( \38654 , \38486 , \38476 );
nand \U$38312 ( \38655 , \38654 , \38487 );
xor \U$38313 ( \38656 , \38514 , \38541 );
xor \U$38314 ( \38657 , \38656 , \38568 );
and \U$38315 ( \38658 , \38655 , \38657 );
xor \U$38316 ( \38659 , \38230 , \38237 );
xor \U$38317 ( \38660 , \38659 , \38246 );
xor \U$38318 ( \38661 , \38346 , \38351 );
xor \U$38319 ( \38662 , \38660 , \38661 );
xor \U$38320 ( \38663 , \38514 , \38541 );
xor \U$38321 ( \38664 , \38663 , \38568 );
and \U$38322 ( \38665 , \38662 , \38664 );
and \U$38323 ( \38666 , \38655 , \38662 );
or \U$38324 ( \38667 , \38658 , \38665 , \38666 );
not \U$38325 ( \38668 , \3406 );
and \U$38326 ( \38669 , \3254 , RI986f778_58);
and \U$38327 ( \38670 , RI986fa48_64, \3252 );
nor \U$38328 ( \38671 , \38669 , \38670 );
not \U$38329 ( \38672 , \38671 );
or \U$38330 ( \38673 , \38668 , \38672 );
or \U$38331 ( \38674 , \38671 , \3406 );
nand \U$38332 ( \38675 , \38673 , \38674 );
and \U$38333 ( \38676 , \2464 , RI986e698_22);
and \U$38334 ( \38677 , RI986f868_60, \2462 );
nor \U$38335 ( \38678 , \38676 , \38677 );
and \U$38336 ( \38679 , \38678 , \2468 );
not \U$38337 ( \38680 , \38678 );
and \U$38338 ( \38681 , \38680 , \2263 );
nor \U$38339 ( \38682 , \38679 , \38681 );
xor \U$38340 ( \38683 , \38675 , \38682 );
not \U$38341 ( \38684 , \3412 );
and \U$38342 ( \38685 , \3683 , RI986f958_62);
and \U$38343 ( \38686 , RI986f4a8_52, \3681 );
nor \U$38344 ( \38687 , \38685 , \38686 );
not \U$38345 ( \38688 , \38687 );
or \U$38346 ( \38689 , \38684 , \38688 );
or \U$38347 ( \38690 , \38687 , \3412 );
nand \U$38348 ( \38691 , \38689 , \38690 );
and \U$38349 ( \38692 , \38683 , \38691 );
and \U$38350 ( \38693 , \38675 , \38682 );
or \U$38351 ( \38694 , \38692 , \38693 );
and \U$38352 ( \38695 , \5881 , RI986dd38_2);
and \U$38353 ( \38696 , RI986e1e8_12, \5879 );
nor \U$38354 ( \38697 , \38695 , \38696 );
and \U$38355 ( \38698 , \38697 , \5594 );
not \U$38356 ( \38699 , \38697 );
and \U$38357 ( \38700 , \38699 , \5885 );
nor \U$38358 ( \38701 , \38698 , \38700 );
nand \U$38359 ( \38702 , RI986e3c8_16, \7079 );
and \U$38360 ( \38703 , \38702 , \6710 );
not \U$38361 ( \38704 , \38702 );
and \U$38362 ( \38705 , \38704 , \6709 );
nor \U$38363 ( \38706 , \38703 , \38705 );
xor \U$38364 ( \38707 , \38701 , \38706 );
and \U$38365 ( \38708 , \6453 , RI986e0f8_10);
and \U$38366 ( \38709 , RI986e2d8_14, \6451 );
nor \U$38367 ( \38710 , \38708 , \38709 );
and \U$38368 ( \38711 , \38710 , \6190 );
not \U$38369 ( \38712 , \38710 );
and \U$38370 ( \38713 , \38712 , \6705 );
nor \U$38371 ( \38714 , \38711 , \38713 );
and \U$38372 ( \38715 , \38707 , \38714 );
and \U$38373 ( \38716 , \38701 , \38706 );
or \U$38374 ( \38717 , \38715 , \38716 );
xor \U$38375 ( \38718 , \38694 , \38717 );
and \U$38376 ( \38719 , \5318 , RI986df18_6);
and \U$38377 ( \38720 , RI986de28_4, \5316 );
nor \U$38378 ( \38721 , \38719 , \38720 );
and \U$38379 ( \38722 , \38721 , \5052 );
not \U$38380 ( \38723 , \38721 );
and \U$38381 ( \38724 , \38723 , \5322 );
nor \U$38382 ( \38725 , \38722 , \38724 );
and \U$38383 ( \38726 , \4203 , RI986f3b8_50);
and \U$38384 ( \38727 , RI986f598_54, \4201 );
nor \U$38385 ( \38728 , \38726 , \38727 );
and \U$38386 ( \38729 , \38728 , \4207 );
not \U$38387 ( \38730 , \38728 );
and \U$38388 ( \38731 , \38730 , \3923 );
nor \U$38389 ( \38732 , \38729 , \38731 );
xor \U$38390 ( \38733 , \38725 , \38732 );
not \U$38391 ( \38734 , \4519 );
and \U$38392 ( \38735 , \4710 , RI986f688_56);
and \U$38393 ( \38736 , RI986e008_8, \4708 );
nor \U$38394 ( \38737 , \38735 , \38736 );
not \U$38395 ( \38738 , \38737 );
or \U$38396 ( \38739 , \38734 , \38738 );
or \U$38397 ( \38740 , \38737 , \4519 );
nand \U$38398 ( \38741 , \38739 , \38740 );
and \U$38399 ( \38742 , \38733 , \38741 );
and \U$38400 ( \38743 , \38725 , \38732 );
or \U$38401 ( \38744 , \38742 , \38743 );
and \U$38402 ( \38745 , \38718 , \38744 );
and \U$38403 ( \38746 , \38694 , \38717 );
or \U$38404 ( \38747 , \38745 , \38746 );
nand \U$38405 ( \38748 , RI98710c8_112, RI9871fc8_144);
not \U$38406 ( \38749 , \38748 );
not \U$38407 ( \38750 , RI9870d08_104);
nor \U$38408 ( \38751 , \38750 , \407 );
xor \U$38409 ( \38752 , \38749 , \38751 );
and \U$38410 ( \38753 , \416 , RI9870d08_104);
and \U$38411 ( \38754 , RI98712a8_116, \414 );
nor \U$38412 ( \38755 , \38753 , \38754 );
and \U$38413 ( \38756 , \38755 , \422 );
not \U$38414 ( \38757 , \38755 );
and \U$38415 ( \38758 , \38757 , \421 );
nor \U$38416 ( \38759 , \38756 , \38758 );
not \U$38417 ( \38760 , \487 );
and \U$38418 ( \38761 , \395 , RI9871488_120);
and \U$38419 ( \38762 , RI9871758_126, \393 );
nor \U$38420 ( \38763 , \38761 , \38762 );
not \U$38421 ( \38764 , \38763 );
or \U$38422 ( \38765 , \38760 , \38764 );
or \U$38423 ( \38766 , \38763 , \386 );
nand \U$38424 ( \38767 , \38765 , \38766 );
xor \U$38425 ( \38768 , \38759 , \38767 );
not \U$38426 ( \38769 , \345 );
and \U$38427 ( \38770 , \354 , RI98711b8_114);
and \U$38428 ( \38771 , RI9871398_118, \352 );
nor \U$38429 ( \38772 , \38770 , \38771 );
not \U$38430 ( \38773 , \38772 );
or \U$38431 ( \38774 , \38769 , \38773 );
or \U$38432 ( \38775 , \38772 , \361 );
nand \U$38433 ( \38776 , \38774 , \38775 );
and \U$38434 ( \38777 , \38768 , \38776 );
and \U$38435 ( \38778 , \38759 , \38767 );
or \U$38436 ( \38779 , \38777 , \38778 );
and \U$38437 ( \38780 , \38752 , \38779 );
and \U$38438 ( \38781 , \38749 , \38751 );
or \U$38439 ( \38782 , \38780 , \38781 );
xor \U$38440 ( \38783 , \38747 , \38782 );
and \U$38441 ( \38784 , \1311 , RI986eff8_42);
and \U$38442 ( \38785 , RI986f2c8_48, \1309 );
nor \U$38443 ( \38786 , \38784 , \38785 );
and \U$38444 ( \38787 , \38786 , \1458 );
not \U$38445 ( \38788 , \38786 );
and \U$38446 ( \38789 , \38788 , \1318 );
nor \U$38447 ( \38790 , \38787 , \38789 );
not \U$38448 ( \38791 , \1462 );
and \U$38449 ( \38792 , \2042 , RI986f1d8_46);
and \U$38450 ( \38793 , RI986e5a8_20, \2040 );
nor \U$38451 ( \38794 , \38792 , \38793 );
not \U$38452 ( \38795 , \38794 );
or \U$38453 ( \38796 , \38791 , \38795 );
or \U$38454 ( \38797 , \38794 , \1462 );
nand \U$38455 ( \38798 , \38796 , \38797 );
xor \U$38456 ( \38799 , \38790 , \38798 );
and \U$38457 ( \38800 , \2274 , RI986e4b8_18);
and \U$38458 ( \38801 , RI986e788_24, \2272 );
nor \U$38459 ( \38802 , \38800 , \38801 );
and \U$38460 ( \38803 , \38802 , \2030 );
not \U$38461 ( \38804 , \38802 );
and \U$38462 ( \38805 , \38804 , \2031 );
nor \U$38463 ( \38806 , \38803 , \38805 );
and \U$38464 ( \38807 , \38799 , \38806 );
and \U$38465 ( \38808 , \38790 , \38798 );
or \U$38466 ( \38809 , \38807 , \38808 );
not \U$38467 ( \38810 , \365 );
and \U$38468 ( \38811 , \376 , RI9871848_128);
and \U$38469 ( \38812 , RI9871578_122, \374 );
nor \U$38470 ( \38813 , \38811 , \38812 );
not \U$38471 ( \38814 , \38813 );
or \U$38472 ( \38815 , \38810 , \38814 );
or \U$38473 ( \38816 , \38813 , \367 );
nand \U$38474 ( \38817 , \38815 , \38816 );
and \U$38475 ( \38818 , \438 , RI986ea58_30);
and \U$38476 ( \38819 , RI986e968_28, \436 );
nor \U$38477 ( \38820 , \38818 , \38819 );
and \U$38478 ( \38821 , \38820 , \444 );
not \U$38479 ( \38822 , \38820 );
and \U$38480 ( \38823 , \38822 , \443 );
nor \U$38481 ( \38824 , \38821 , \38823 );
xor \U$38482 ( \38825 , \38817 , \38824 );
not \U$38483 ( \38826 , \456 );
and \U$38484 ( \38827 , \465 , RI9871668_124);
and \U$38485 ( \38828 , RI986eb48_32, \463 );
nor \U$38486 ( \38829 , \38827 , \38828 );
not \U$38487 ( \38830 , \38829 );
or \U$38488 ( \38831 , \38826 , \38830 );
or \U$38489 ( \38832 , \38829 , \456 );
nand \U$38490 ( \38833 , \38831 , \38832 );
and \U$38491 ( \38834 , \38825 , \38833 );
and \U$38492 ( \38835 , \38817 , \38824 );
or \U$38493 ( \38836 , \38834 , \38835 );
xor \U$38494 ( \38837 , \38809 , \38836 );
and \U$38495 ( \38838 , \1329 , RI986ed28_36);
and \U$38496 ( \38839 , RI986f0e8_44, \1327 );
nor \U$38497 ( \38840 , \38838 , \38839 );
and \U$38498 ( \38841 , \38840 , \1336 );
not \U$38499 ( \38842 , \38840 );
and \U$38500 ( \38843 , \38842 , \1337 );
nor \U$38501 ( \38844 , \38841 , \38843 );
and \U$38502 ( \38845 , \776 , RI986e878_26);
and \U$38503 ( \38846 , RI986ef08_40, \774 );
nor \U$38504 ( \38847 , \38845 , \38846 );
and \U$38505 ( \38848 , \38847 , \474 );
not \U$38506 ( \38849 , \38847 );
and \U$38507 ( \38850 , \38849 , \451 );
nor \U$38508 ( \38851 , \38848 , \38850 );
xor \U$38509 ( \38852 , \38844 , \38851 );
not \U$38510 ( \38853 , \1128 );
and \U$38511 ( \38854 , \1293 , RI986ee18_38);
and \U$38512 ( \38855 , RI986ec38_34, \1291 );
nor \U$38513 ( \38856 , \38854 , \38855 );
not \U$38514 ( \38857 , \38856 );
or \U$38515 ( \38858 , \38853 , \38857 );
or \U$38516 ( \38859 , \38856 , \1301 );
nand \U$38517 ( \38860 , \38858 , \38859 );
and \U$38518 ( \38861 , \38852 , \38860 );
and \U$38519 ( \38862 , \38844 , \38851 );
or \U$38520 ( \38863 , \38861 , \38862 );
and \U$38521 ( \38864 , \38837 , \38863 );
and \U$38522 ( \38865 , \38809 , \38836 );
or \U$38523 ( \38866 , \38864 , \38865 );
and \U$38524 ( \38867 , \38783 , \38866 );
and \U$38525 ( \38868 , \38747 , \38782 );
or \U$38526 ( \38869 , \38867 , \38868 );
xor \U$38527 ( \38870 , \38667 , \38869 );
xor \U$38528 ( \38871 , \38457 , \38465 );
xor \U$38529 ( \38872 , \38871 , \38473 );
xor \U$38530 ( \38873 , \38522 , \38529 );
xor \U$38531 ( \38874 , \38873 , \38538 );
and \U$38532 ( \38875 , \38872 , \38874 );
xor \U$38533 ( \38876 , \38549 , \38556 );
xor \U$38534 ( \38877 , \38876 , \38565 );
xor \U$38535 ( \38878 , \38522 , \38529 );
xor \U$38536 ( \38879 , \38878 , \38538 );
and \U$38537 ( \38880 , \38877 , \38879 );
and \U$38538 ( \38881 , \38872 , \38877 );
or \U$38539 ( \38882 , \38875 , \38880 , \38881 );
xor \U$38540 ( \38883 , \38427 , \38435 );
xor \U$38541 ( \38884 , \38883 , \38443 );
xor \U$38542 ( \38885 , \38495 , \38502 );
xor \U$38543 ( \38886 , \38885 , \38511 );
xor \U$38544 ( \38887 , \38884 , \38886 );
xor \U$38545 ( \38888 , \38382 , \38389 );
xor \U$38546 ( \38889 , \38888 , \38398 );
and \U$38547 ( \38890 , \38887 , \38889 );
and \U$38548 ( \38891 , \38884 , \38886 );
or \U$38549 ( \38892 , \38890 , \38891 );
xor \U$38550 ( \38893 , \38882 , \38892 );
xor \U$38551 ( \38894 , \38096 , \38103 );
xor \U$38552 ( \38895 , \38894 , \38112 );
xor \U$38553 ( \38896 , \38361 , \38366 );
xor \U$38554 ( \38897 , \38895 , \38896 );
and \U$38555 ( \38898 , \38893 , \38897 );
and \U$38556 ( \38899 , \38882 , \38892 );
or \U$38557 ( \38900 , \38898 , \38899 );
xor \U$38558 ( \38901 , \38870 , \38900 );
xor \U$38559 ( \38902 , \38644 , \38646 );
xor \U$38560 ( \38903 , \38902 , \38651 );
and \U$38561 ( \38904 , \38901 , \38903 );
and \U$38562 ( \38905 , \38642 , \38901 );
or \U$38563 ( \38906 , \38653 , \38904 , \38905 );
xor \U$38564 ( \38907 , \38374 , \38574 );
xor \U$38565 ( \38908 , \38907 , \38589 );
xor \U$38566 ( \38909 , \38906 , \38908 );
xor \U$38567 ( \38910 , \38701 , \38706 );
xor \U$38568 ( \38911 , \38910 , \38714 );
xor \U$38569 ( \38912 , \38675 , \38682 );
xor \U$38570 ( \38913 , \38912 , \38691 );
and \U$38571 ( \38914 , \38911 , \38913 );
xor \U$38572 ( \38915 , \38725 , \38732 );
xor \U$38573 ( \38916 , \38915 , \38741 );
xor \U$38574 ( \38917 , \38675 , \38682 );
xor \U$38575 ( \38918 , \38917 , \38691 );
and \U$38576 ( \38919 , \38916 , \38918 );
and \U$38577 ( \38920 , \38911 , \38916 );
or \U$38578 ( \38921 , \38914 , \38919 , \38920 );
xor \U$38579 ( \38922 , \38408 , \6710 );
xor \U$38580 ( \38923 , \38922 , \38416 );
xor \U$38581 ( \38924 , \38921 , \38923 );
xor \U$38582 ( \38925 , \38817 , \38824 );
xor \U$38583 ( \38926 , \38925 , \38833 );
xor \U$38584 ( \38927 , \38844 , \38851 );
xor \U$38585 ( \38928 , \38927 , \38860 );
and \U$38586 ( \38929 , \38926 , \38928 );
xor \U$38587 ( \38930 , \38790 , \38798 );
xor \U$38588 ( \38931 , \38930 , \38806 );
xor \U$38589 ( \38932 , \38844 , \38851 );
xor \U$38590 ( \38933 , \38932 , \38860 );
and \U$38591 ( \38934 , \38931 , \38933 );
and \U$38592 ( \38935 , \38926 , \38931 );
or \U$38593 ( \38936 , \38929 , \38934 , \38935 );
and \U$38594 ( \38937 , \38924 , \38936 );
and \U$38595 ( \38938 , \38921 , \38923 );
or \U$38596 ( \38939 , \38937 , \38938 );
and \U$38597 ( \38940 , \2274 , RI986e5a8_20);
and \U$38598 ( \38941 , RI986e4b8_18, \2272 );
nor \U$38599 ( \38942 , \38940 , \38941 );
and \U$38600 ( \38943 , \38942 , \2030 );
not \U$38601 ( \38944 , \38942 );
and \U$38602 ( \38945 , \38944 , \2031 );
nor \U$38603 ( \38946 , \38943 , \38945 );
not \U$38604 ( \38947 , \1462 );
and \U$38605 ( \38948 , \2042 , RI986f2c8_48);
and \U$38606 ( \38949 , RI986f1d8_46, \2040 );
nor \U$38607 ( \38950 , \38948 , \38949 );
not \U$38608 ( \38951 , \38950 );
or \U$38609 ( \38952 , \38947 , \38951 );
or \U$38610 ( \38953 , \38950 , \1462 );
nand \U$38611 ( \38954 , \38952 , \38953 );
xor \U$38612 ( \38955 , \38946 , \38954 );
and \U$38613 ( \38956 , \2464 , RI986e788_24);
and \U$38614 ( \38957 , RI986e698_22, \2462 );
nor \U$38615 ( \38958 , \38956 , \38957 );
and \U$38616 ( \38959 , \38958 , \2468 );
not \U$38617 ( \38960 , \38958 );
and \U$38618 ( \38961 , \38960 , \2263 );
nor \U$38619 ( \38962 , \38959 , \38961 );
and \U$38620 ( \38963 , \38955 , \38962 );
and \U$38621 ( \38964 , \38946 , \38954 );
or \U$38622 ( \38965 , \38963 , \38964 );
not \U$38623 ( \38966 , \456 );
and \U$38624 ( \38967 , \465 , RI9871578_122);
and \U$38625 ( \38968 , RI9871668_124, \463 );
nor \U$38626 ( \38969 , \38967 , \38968 );
not \U$38627 ( \38970 , \38969 );
or \U$38628 ( \38971 , \38966 , \38970 );
or \U$38629 ( \38972 , \38969 , \456 );
nand \U$38630 ( \38973 , \38971 , \38972 );
and \U$38631 ( \38974 , \776 , RI986e968_28);
and \U$38632 ( \38975 , RI986e878_26, \774 );
nor \U$38633 ( \38976 , \38974 , \38975 );
and \U$38634 ( \38977 , \38976 , \474 );
not \U$38635 ( \38978 , \38976 );
and \U$38636 ( \38979 , \38978 , \451 );
nor \U$38637 ( \38980 , \38977 , \38979 );
xor \U$38638 ( \38981 , \38973 , \38980 );
and \U$38639 ( \38982 , \438 , RI986eb48_32);
and \U$38640 ( \38983 , RI986ea58_30, \436 );
nor \U$38641 ( \38984 , \38982 , \38983 );
and \U$38642 ( \38985 , \38984 , \444 );
not \U$38643 ( \38986 , \38984 );
and \U$38644 ( \38987 , \38986 , \443 );
nor \U$38645 ( \38988 , \38985 , \38987 );
and \U$38646 ( \38989 , \38981 , \38988 );
and \U$38647 ( \38990 , \38973 , \38980 );
or \U$38648 ( \38991 , \38989 , \38990 );
xor \U$38649 ( \38992 , \38965 , \38991 );
not \U$38650 ( \38993 , \1128 );
and \U$38651 ( \38994 , \1293 , RI986ef08_40);
and \U$38652 ( \38995 , RI986ee18_38, \1291 );
nor \U$38653 ( \38996 , \38994 , \38995 );
not \U$38654 ( \38997 , \38996 );
or \U$38655 ( \38998 , \38993 , \38997 );
or \U$38656 ( \38999 , \38996 , \1128 );
nand \U$38657 ( \39000 , \38998 , \38999 );
and \U$38658 ( \39001 , \1329 , RI986ec38_34);
and \U$38659 ( \39002 , RI986ed28_36, \1327 );
nor \U$38660 ( \39003 , \39001 , \39002 );
and \U$38661 ( \39004 , \39003 , \1336 );
not \U$38662 ( \39005 , \39003 );
and \U$38663 ( \39006 , \39005 , \1337 );
nor \U$38664 ( \39007 , \39004 , \39006 );
xor \U$38665 ( \39008 , \39000 , \39007 );
and \U$38666 ( \39009 , \1311 , RI986f0e8_44);
and \U$38667 ( \39010 , RI986eff8_42, \1309 );
nor \U$38668 ( \39011 , \39009 , \39010 );
and \U$38669 ( \39012 , \39011 , \1319 );
not \U$38670 ( \39013 , \39011 );
and \U$38671 ( \39014 , \39013 , \1318 );
nor \U$38672 ( \39015 , \39012 , \39014 );
and \U$38673 ( \39016 , \39008 , \39015 );
and \U$38674 ( \39017 , \39000 , \39007 );
or \U$38675 ( \39018 , \39016 , \39017 );
and \U$38676 ( \39019 , \38992 , \39018 );
and \U$38677 ( \39020 , \38965 , \38991 );
or \U$38678 ( \39021 , \39019 , \39020 );
and \U$38679 ( \39022 , \4203 , RI986f4a8_52);
and \U$38680 ( \39023 , RI986f3b8_50, \4201 );
nor \U$38681 ( \39024 , \39022 , \39023 );
and \U$38682 ( \39025 , \39024 , \4207 );
not \U$38683 ( \39026 , \39024 );
and \U$38684 ( \39027 , \39026 , \3923 );
nor \U$38685 ( \39028 , \39025 , \39027 );
not \U$38686 ( \39029 , \3406 );
and \U$38687 ( \39030 , \3254 , RI986f868_60);
and \U$38688 ( \39031 , RI986f778_58, \3252 );
nor \U$38689 ( \39032 , \39030 , \39031 );
not \U$38690 ( \39033 , \39032 );
or \U$38691 ( \39034 , \39029 , \39033 );
or \U$38692 ( \39035 , \39032 , \2935 );
nand \U$38693 ( \39036 , \39034 , \39035 );
xor \U$38694 ( \39037 , \39028 , \39036 );
not \U$38695 ( \39038 , \3412 );
and \U$38696 ( \39039 , \3683 , RI986fa48_64);
and \U$38697 ( \39040 , RI986f958_62, \3681 );
nor \U$38698 ( \39041 , \39039 , \39040 );
not \U$38699 ( \39042 , \39041 );
or \U$38700 ( \39043 , \39038 , \39042 );
or \U$38701 ( \39044 , \39041 , \3918 );
nand \U$38702 ( \39045 , \39043 , \39044 );
and \U$38703 ( \39046 , \39037 , \39045 );
and \U$38704 ( \39047 , \39028 , \39036 );
or \U$38705 ( \39048 , \39046 , \39047 );
and \U$38706 ( \39049 , \6453 , RI986e1e8_12);
and \U$38707 ( \39050 , RI986e0f8_10, \6451 );
nor \U$38708 ( \39051 , \39049 , \39050 );
and \U$38709 ( \39052 , \39051 , \6190 );
not \U$38710 ( \39053 , \39051 );
and \U$38711 ( \39054 , \39053 , \6180 );
nor \U$38712 ( \39055 , \39052 , \39054 );
xor \U$38713 ( \39056 , \39055 , \7480 );
and \U$38714 ( \39057 , \7079 , RI986e2d8_14);
and \U$38715 ( \39058 , RI986e3c8_16, \7077 );
nor \U$38716 ( \39059 , \39057 , \39058 );
and \U$38717 ( \39060 , \39059 , \6710 );
not \U$38718 ( \39061 , \39059 );
and \U$38719 ( \39062 , \39061 , \6709 );
nor \U$38720 ( \39063 , \39060 , \39062 );
and \U$38721 ( \39064 , \39056 , \39063 );
and \U$38722 ( \39065 , \39055 , \7480 );
or \U$38723 ( \39066 , \39064 , \39065 );
xor \U$38724 ( \39067 , \39048 , \39066 );
and \U$38725 ( \39068 , \5881 , RI986de28_4);
and \U$38726 ( \39069 , RI986dd38_2, \5879 );
nor \U$38727 ( \39070 , \39068 , \39069 );
and \U$38728 ( \39071 , \39070 , \5594 );
not \U$38729 ( \39072 , \39070 );
and \U$38730 ( \39073 , \39072 , \5885 );
nor \U$38731 ( \39074 , \39071 , \39073 );
not \U$38732 ( \39075 , \4521 );
and \U$38733 ( \39076 , \4710 , RI986f598_54);
and \U$38734 ( \39077 , RI986f688_56, \4708 );
nor \U$38735 ( \39078 , \39076 , \39077 );
not \U$38736 ( \39079 , \39078 );
or \U$38737 ( \39080 , \39075 , \39079 );
or \U$38738 ( \39081 , \39078 , \4519 );
nand \U$38739 ( \39082 , \39080 , \39081 );
xor \U$38740 ( \39083 , \39074 , \39082 );
and \U$38741 ( \39084 , \5318 , RI986e008_8);
and \U$38742 ( \39085 , RI986df18_6, \5316 );
nor \U$38743 ( \39086 , \39084 , \39085 );
and \U$38744 ( \39087 , \39086 , \5052 );
not \U$38745 ( \39088 , \39086 );
and \U$38746 ( \39089 , \39088 , \5322 );
nor \U$38747 ( \39090 , \39087 , \39089 );
and \U$38748 ( \39091 , \39083 , \39090 );
and \U$38749 ( \39092 , \39074 , \39082 );
or \U$38750 ( \39093 , \39091 , \39092 );
and \U$38751 ( \39094 , \39067 , \39093 );
and \U$38752 ( \39095 , \39048 , \39066 );
or \U$38753 ( \39096 , \39094 , \39095 );
xor \U$38754 ( \39097 , \39021 , \39096 );
not \U$38755 ( \39098 , \361 );
and \U$38756 ( \39099 , \354 , RI98712a8_116);
and \U$38757 ( \39100 , RI98711b8_114, \352 );
nor \U$38758 ( \39101 , \39099 , \39100 );
not \U$38759 ( \39102 , \39101 );
or \U$38760 ( \39103 , \39098 , \39102 );
or \U$38761 ( \39104 , \39101 , \345 );
nand \U$38762 ( \39105 , \39103 , \39104 );
not \U$38763 ( \39106 , \367 );
and \U$38764 ( \39107 , \376 , RI9871758_126);
and \U$38765 ( \39108 , RI9871848_128, \374 );
nor \U$38766 ( \39109 , \39107 , \39108 );
not \U$38767 ( \39110 , \39109 );
or \U$38768 ( \39111 , \39106 , \39110 );
or \U$38769 ( \39112 , \39109 , \367 );
nand \U$38770 ( \39113 , \39111 , \39112 );
xor \U$38771 ( \39114 , \39105 , \39113 );
not \U$38772 ( \39115 , \487 );
and \U$38773 ( \39116 , \395 , RI9871398_118);
and \U$38774 ( \39117 , RI9871488_120, \393 );
nor \U$38775 ( \39118 , \39116 , \39117 );
not \U$38776 ( \39119 , \39118 );
or \U$38777 ( \39120 , \39115 , \39119 );
or \U$38778 ( \39121 , \39118 , \386 );
nand \U$38779 ( \39122 , \39120 , \39121 );
and \U$38780 ( \39123 , \39114 , \39122 );
and \U$38781 ( \39124 , \39105 , \39113 );
or \U$38782 ( \39125 , \39123 , \39124 );
xor \U$38783 ( \39126 , \39125 , \38748 );
xor \U$38784 ( \39127 , \38759 , \38767 );
xor \U$38785 ( \39128 , \39127 , \38776 );
and \U$38786 ( \39129 , \39126 , \39128 );
and \U$38787 ( \39130 , \39125 , \38748 );
or \U$38788 ( \39131 , \39129 , \39130 );
and \U$38789 ( \39132 , \39097 , \39131 );
and \U$38790 ( \39133 , \39021 , \39096 );
or \U$38791 ( \39134 , \39132 , \39133 );
xor \U$38792 ( \39135 , \38939 , \39134 );
xor \U$38793 ( \39136 , \38749 , \38751 );
xor \U$38794 ( \39137 , \39136 , \38779 );
xor \U$38795 ( \39138 , \38884 , \38886 );
xor \U$38796 ( \39139 , \39138 , \38889 );
and \U$38797 ( \39140 , \39137 , \39139 );
xor \U$38798 ( \39141 , \38522 , \38529 );
xor \U$38799 ( \39142 , \39141 , \38538 );
xor \U$38800 ( \39143 , \38872 , \38877 );
xor \U$38801 ( \39144 , \39142 , \39143 );
xor \U$38802 ( \39145 , \38884 , \38886 );
xor \U$38803 ( \39146 , \39145 , \38889 );
and \U$38804 ( \39147 , \39144 , \39146 );
and \U$38805 ( \39148 , \39137 , \39144 );
or \U$38806 ( \39149 , \39140 , \39147 , \39148 );
and \U$38807 ( \39150 , \39135 , \39149 );
and \U$38808 ( \39151 , \38939 , \39134 );
or \U$38809 ( \39152 , \39150 , \39151 );
xor \U$38810 ( \39153 , \38356 , \38358 );
xor \U$38811 ( \39154 , \39153 , \38371 );
xor \U$38812 ( \39155 , \39152 , \39154 );
xor \U$38813 ( \39156 , \38401 , \38419 );
xor \U$38814 ( \39157 , \39156 , \38446 );
xor \U$38815 ( \39158 , \38882 , \38892 );
xor \U$38816 ( \39159 , \39158 , \38897 );
and \U$38817 ( \39160 , \39157 , \39159 );
xor \U$38818 ( \39161 , \38514 , \38541 );
xor \U$38819 ( \39162 , \39161 , \38568 );
xor \U$38820 ( \39163 , \38655 , \38662 );
xor \U$38821 ( \39164 , \39162 , \39163 );
xor \U$38822 ( \39165 , \38882 , \38892 );
xor \U$38823 ( \39166 , \39165 , \38897 );
and \U$38824 ( \39167 , \39164 , \39166 );
and \U$38825 ( \39168 , \39157 , \39164 );
or \U$38826 ( \39169 , \39160 , \39167 , \39168 );
and \U$38827 ( \39170 , \39155 , \39169 );
and \U$38828 ( \39171 , \39152 , \39154 );
or \U$38829 ( \39172 , \39170 , \39171 );
and \U$38830 ( \39173 , \38909 , \39172 );
and \U$38831 ( \39174 , \38906 , \38908 );
or \U$38832 ( \39175 , \39173 , \39174 );
xor \U$38833 ( \39176 , \38667 , \38869 );
and \U$38834 ( \39177 , \39176 , \38900 );
and \U$38835 ( \39178 , \38667 , \38869 );
or \U$38836 ( \39179 , \39177 , \39178 );
xor \U$38837 ( \39180 , \38644 , \38646 );
and \U$38838 ( \39181 , \39180 , \38651 );
and \U$38839 ( \39182 , \38644 , \38646 );
or \U$38840 ( \39183 , \39181 , \39182 );
xor \U$38841 ( \39184 , \39179 , \39183 );
xor \U$38842 ( \39185 , \38080 , \38082 );
xor \U$38843 ( \39186 , \39185 , \38085 );
xor \U$38844 ( \39187 , \38597 , \38602 );
xor \U$38845 ( \39188 , \39186 , \39187 );
and \U$38846 ( \39189 , \39184 , \39188 );
and \U$38847 ( \39190 , \39179 , \39183 );
or \U$38848 ( \39191 , \39189 , \39190 );
xor \U$38849 ( \39192 , \38612 , \38616 );
xor \U$38850 ( \39193 , \39191 , \39192 );
xor \U$38851 ( \39194 , \38592 , \38594 );
xor \U$38852 ( \39195 , \39194 , \38607 );
xor \U$38853 ( \39196 , \39193 , \39195 );
and \U$38854 ( \39197 , \39175 , \39196 );
xor \U$38855 ( \39198 , \38946 , \38954 );
xor \U$38856 ( \39199 , \39198 , \38962 );
xor \U$38857 ( \39200 , \39000 , \39007 );
xor \U$38858 ( \39201 , \39200 , \39015 );
and \U$38859 ( \39202 , \39199 , \39201 );
xor \U$38860 ( \39203 , \39028 , \39036 );
xor \U$38861 ( \39204 , \39203 , \39045 );
xor \U$38862 ( \39205 , \39000 , \39007 );
xor \U$38863 ( \39206 , \39205 , \39015 );
and \U$38864 ( \39207 , \39204 , \39206 );
and \U$38865 ( \39208 , \39199 , \39204 );
or \U$38866 ( \39209 , \39202 , \39207 , \39208 );
xor \U$38867 ( \39210 , \38973 , \38980 );
xor \U$38868 ( \39211 , \39210 , \38988 );
not \U$38869 ( \39212 , RI9870c18_102);
nor \U$38870 ( \39213 , \39212 , \407 );
xor \U$38871 ( \39214 , \39211 , \39213 );
xor \U$38872 ( \39215 , \39105 , \39113 );
xor \U$38873 ( \39216 , \39215 , \39122 );
and \U$38874 ( \39217 , \39214 , \39216 );
and \U$38875 ( \39218 , \39211 , \39213 );
or \U$38876 ( \39219 , \39217 , \39218 );
xor \U$38877 ( \39220 , \39209 , \39219 );
xor \U$38878 ( \39221 , \38675 , \38682 );
xor \U$38879 ( \39222 , \39221 , \38691 );
xor \U$38880 ( \39223 , \38911 , \38916 );
xor \U$38881 ( \39224 , \39222 , \39223 );
and \U$38882 ( \39225 , \39220 , \39224 );
and \U$38883 ( \39226 , \39209 , \39219 );
or \U$38884 ( \39227 , \39225 , \39226 );
and \U$38885 ( \39228 , \4203 , RI986f958_62);
and \U$38886 ( \39229 , RI986f4a8_52, \4201 );
nor \U$38887 ( \39230 , \39228 , \39229 );
and \U$38888 ( \39231 , \39230 , \4207 );
not \U$38889 ( \39232 , \39230 );
and \U$38890 ( \39233 , \39232 , \3923 );
nor \U$38891 ( \39234 , \39231 , \39233 );
not \U$38892 ( \39235 , \2935 );
and \U$38893 ( \39236 , \3254 , RI986e698_22);
and \U$38894 ( \39237 , RI986f868_60, \3252 );
nor \U$38895 ( \39238 , \39236 , \39237 );
not \U$38896 ( \39239 , \39238 );
or \U$38897 ( \39240 , \39235 , \39239 );
or \U$38898 ( \39241 , \39238 , \3406 );
nand \U$38899 ( \39242 , \39240 , \39241 );
xor \U$38900 ( \39243 , \39234 , \39242 );
not \U$38901 ( \39244 , \3918 );
and \U$38902 ( \39245 , \3683 , RI986f778_58);
and \U$38903 ( \39246 , RI986fa48_64, \3681 );
nor \U$38904 ( \39247 , \39245 , \39246 );
not \U$38905 ( \39248 , \39247 );
or \U$38906 ( \39249 , \39244 , \39248 );
or \U$38907 ( \39250 , \39247 , \3918 );
nand \U$38908 ( \39251 , \39249 , \39250 );
and \U$38909 ( \39252 , \39243 , \39251 );
and \U$38910 ( \39253 , \39234 , \39242 );
or \U$38911 ( \39254 , \39252 , \39253 );
and \U$38912 ( \39255 , \6453 , RI986dd38_2);
and \U$38913 ( \39256 , RI986e1e8_12, \6451 );
nor \U$38914 ( \39257 , \39255 , \39256 );
and \U$38915 ( \39258 , \39257 , \6190 );
not \U$38916 ( \39259 , \39257 );
and \U$38917 ( \39260 , \39259 , \6705 );
nor \U$38918 ( \39261 , \39258 , \39260 );
nand \U$38919 ( \39262 , RI986e3c8_16, \7729 );
and \U$38920 ( \39263 , \39262 , \7480 );
not \U$38921 ( \39264 , \39262 );
and \U$38922 ( \39265 , \39264 , \7733 );
nor \U$38923 ( \39266 , \39263 , \39265 );
xor \U$38924 ( \39267 , \39261 , \39266 );
and \U$38925 ( \39268 , \7079 , RI986e0f8_10);
and \U$38926 ( \39269 , RI986e2d8_14, \7077 );
nor \U$38927 ( \39270 , \39268 , \39269 );
and \U$38928 ( \39271 , \39270 , \6710 );
not \U$38929 ( \39272 , \39270 );
and \U$38930 ( \39273 , \39272 , \6709 );
nor \U$38931 ( \39274 , \39271 , \39273 );
and \U$38932 ( \39275 , \39267 , \39274 );
and \U$38933 ( \39276 , \39261 , \39266 );
or \U$38934 ( \39277 , \39275 , \39276 );
xor \U$38935 ( \39278 , \39254 , \39277 );
and \U$38936 ( \39279 , \5881 , RI986df18_6);
and \U$38937 ( \39280 , RI986de28_4, \5879 );
nor \U$38938 ( \39281 , \39279 , \39280 );
and \U$38939 ( \39282 , \39281 , \5594 );
not \U$38940 ( \39283 , \39281 );
and \U$38941 ( \39284 , \39283 , \5885 );
nor \U$38942 ( \39285 , \39282 , \39284 );
not \U$38943 ( \39286 , \4521 );
and \U$38944 ( \39287 , \4710 , RI986f3b8_50);
and \U$38945 ( \39288 , RI986f598_54, \4708 );
nor \U$38946 ( \39289 , \39287 , \39288 );
not \U$38947 ( \39290 , \39289 );
or \U$38948 ( \39291 , \39286 , \39290 );
or \U$38949 ( \39292 , \39289 , \4519 );
nand \U$38950 ( \39293 , \39291 , \39292 );
xor \U$38951 ( \39294 , \39285 , \39293 );
and \U$38952 ( \39295 , \5318 , RI986f688_56);
and \U$38953 ( \39296 , RI986e008_8, \5316 );
nor \U$38954 ( \39297 , \39295 , \39296 );
and \U$38955 ( \39298 , \39297 , \5052 );
not \U$38956 ( \39299 , \39297 );
and \U$38957 ( \39300 , \39299 , \5322 );
nor \U$38958 ( \39301 , \39298 , \39300 );
and \U$38959 ( \39302 , \39294 , \39301 );
and \U$38960 ( \39303 , \39285 , \39293 );
or \U$38961 ( \39304 , \39302 , \39303 );
and \U$38962 ( \39305 , \39278 , \39304 );
and \U$38963 ( \39306 , \39254 , \39277 );
or \U$38964 ( \39307 , \39305 , \39306 );
nand \U$38965 ( \39308 , RI9870ee8_108, RI9871fc8_144);
and \U$38966 ( \39309 , \416 , RI9870c18_102);
and \U$38967 ( \39310 , RI98710c8_112, \414 );
nor \U$38968 ( \39311 , \39309 , \39310 );
and \U$38969 ( \39312 , \39311 , \421 );
not \U$38970 ( \39313 , \39311 );
and \U$38971 ( \39314 , \39313 , \422 );
nor \U$38972 ( \39315 , \39312 , \39314 );
nand \U$38973 ( \39316 , \39308 , \39315 );
and \U$38974 ( \39317 , \416 , RI98710c8_112);
and \U$38975 ( \39318 , RI9870d08_104, \414 );
nor \U$38976 ( \39319 , \39317 , \39318 );
and \U$38977 ( \39320 , \39319 , \422 );
not \U$38978 ( \39321 , \39319 );
and \U$38979 ( \39322 , \39321 , \421 );
nor \U$38980 ( \39323 , \39320 , \39322 );
xor \U$38981 ( \39324 , \39316 , \39323 );
not \U$38982 ( \39325 , \361 );
and \U$38983 ( \39326 , \354 , RI9870d08_104);
and \U$38984 ( \39327 , RI98712a8_116, \352 );
nor \U$38985 ( \39328 , \39326 , \39327 );
not \U$38986 ( \39329 , \39328 );
or \U$38987 ( \39330 , \39325 , \39329 );
or \U$38988 ( \39331 , \39328 , \361 );
nand \U$38989 ( \39332 , \39330 , \39331 );
not \U$38990 ( \39333 , \367 );
and \U$38991 ( \39334 , \376 , RI9871488_120);
and \U$38992 ( \39335 , RI9871758_126, \374 );
nor \U$38993 ( \39336 , \39334 , \39335 );
not \U$38994 ( \39337 , \39336 );
or \U$38995 ( \39338 , \39333 , \39337 );
or \U$38996 ( \39339 , \39336 , \367 );
nand \U$38997 ( \39340 , \39338 , \39339 );
xor \U$38998 ( \39341 , \39332 , \39340 );
not \U$38999 ( \39342 , \386 );
and \U$39000 ( \39343 , \395 , RI98711b8_114);
and \U$39001 ( \39344 , RI9871398_118, \393 );
nor \U$39002 ( \39345 , \39343 , \39344 );
not \U$39003 ( \39346 , \39345 );
or \U$39004 ( \39347 , \39342 , \39346 );
or \U$39005 ( \39348 , \39345 , \487 );
nand \U$39006 ( \39349 , \39347 , \39348 );
and \U$39007 ( \39350 , \39341 , \39349 );
and \U$39008 ( \39351 , \39332 , \39340 );
or \U$39009 ( \39352 , \39350 , \39351 );
and \U$39010 ( \39353 , \39324 , \39352 );
and \U$39011 ( \39354 , \39316 , \39323 );
or \U$39012 ( \39355 , \39353 , \39354 );
xor \U$39013 ( \39356 , \39307 , \39355 );
and \U$39014 ( \39357 , \2464 , RI986e4b8_18);
and \U$39015 ( \39358 , RI986e788_24, \2462 );
nor \U$39016 ( \39359 , \39357 , \39358 );
and \U$39017 ( \39360 , \39359 , \2468 );
not \U$39018 ( \39361 , \39359 );
and \U$39019 ( \39362 , \39361 , \2263 );
nor \U$39020 ( \39363 , \39360 , \39362 );
not \U$39021 ( \39364 , \2034 );
and \U$39022 ( \39365 , \2042 , RI986eff8_42);
and \U$39023 ( \39366 , RI986f2c8_48, \2040 );
nor \U$39024 ( \39367 , \39365 , \39366 );
not \U$39025 ( \39368 , \39367 );
or \U$39026 ( \39369 , \39364 , \39368 );
or \U$39027 ( \39370 , \39367 , \2034 );
nand \U$39028 ( \39371 , \39369 , \39370 );
xor \U$39029 ( \39372 , \39363 , \39371 );
and \U$39030 ( \39373 , \2274 , RI986f1d8_46);
and \U$39031 ( \39374 , RI986e5a8_20, \2272 );
nor \U$39032 ( \39375 , \39373 , \39374 );
and \U$39033 ( \39376 , \39375 , \2030 );
not \U$39034 ( \39377 , \39375 );
and \U$39035 ( \39378 , \39377 , \2031 );
nor \U$39036 ( \39379 , \39376 , \39378 );
and \U$39037 ( \39380 , \39372 , \39379 );
and \U$39038 ( \39381 , \39363 , \39371 );
or \U$39039 ( \39382 , \39380 , \39381 );
and \U$39040 ( \39383 , \1311 , RI986ed28_36);
and \U$39041 ( \39384 , RI986f0e8_44, \1309 );
nor \U$39042 ( \39385 , \39383 , \39384 );
and \U$39043 ( \39386 , \39385 , \1458 );
not \U$39044 ( \39387 , \39385 );
and \U$39045 ( \39388 , \39387 , \1315 );
nor \U$39046 ( \39389 , \39386 , \39388 );
not \U$39047 ( \39390 , \1301 );
and \U$39048 ( \39391 , \1293 , RI986e878_26);
and \U$39049 ( \39392 , RI986ef08_40, \1291 );
nor \U$39050 ( \39393 , \39391 , \39392 );
not \U$39051 ( \39394 , \39393 );
or \U$39052 ( \39395 , \39390 , \39394 );
or \U$39053 ( \39396 , \39393 , \1301 );
nand \U$39054 ( \39397 , \39395 , \39396 );
xor \U$39055 ( \39398 , \39389 , \39397 );
and \U$39056 ( \39399 , \1329 , RI986ee18_38);
and \U$39057 ( \39400 , RI986ec38_34, \1327 );
nor \U$39058 ( \39401 , \39399 , \39400 );
and \U$39059 ( \39402 , \39401 , \1336 );
not \U$39060 ( \39403 , \39401 );
and \U$39061 ( \39404 , \39403 , \1337 );
nor \U$39062 ( \39405 , \39402 , \39404 );
and \U$39063 ( \39406 , \39398 , \39405 );
and \U$39064 ( \39407 , \39389 , \39397 );
or \U$39065 ( \39408 , \39406 , \39407 );
xor \U$39066 ( \39409 , \39382 , \39408 );
and \U$39067 ( \39410 , \776 , RI986ea58_30);
and \U$39068 ( \39411 , RI986e968_28, \774 );
nor \U$39069 ( \39412 , \39410 , \39411 );
and \U$39070 ( \39413 , \39412 , \474 );
not \U$39071 ( \39414 , \39412 );
and \U$39072 ( \39415 , \39414 , \451 );
nor \U$39073 ( \39416 , \39413 , \39415 );
and \U$39074 ( \39417 , \438 , RI9871668_124);
and \U$39075 ( \39418 , RI986eb48_32, \436 );
nor \U$39076 ( \39419 , \39417 , \39418 );
and \U$39077 ( \39420 , \39419 , \444 );
not \U$39078 ( \39421 , \39419 );
and \U$39079 ( \39422 , \39421 , \443 );
nor \U$39080 ( \39423 , \39420 , \39422 );
xor \U$39081 ( \39424 , \39416 , \39423 );
not \U$39082 ( \39425 , \456 );
and \U$39083 ( \39426 , \465 , RI9871848_128);
and \U$39084 ( \39427 , RI9871578_122, \463 );
nor \U$39085 ( \39428 , \39426 , \39427 );
not \U$39086 ( \39429 , \39428 );
or \U$39087 ( \39430 , \39425 , \39429 );
or \U$39088 ( \39431 , \39428 , \454 );
nand \U$39089 ( \39432 , \39430 , \39431 );
and \U$39090 ( \39433 , \39424 , \39432 );
and \U$39091 ( \39434 , \39416 , \39423 );
or \U$39092 ( \39435 , \39433 , \39434 );
and \U$39093 ( \39436 , \39409 , \39435 );
and \U$39094 ( \39437 , \39382 , \39408 );
or \U$39095 ( \39438 , \39436 , \39437 );
and \U$39096 ( \39439 , \39356 , \39438 );
and \U$39097 ( \39440 , \39307 , \39355 );
or \U$39098 ( \39441 , \39439 , \39440 );
xor \U$39099 ( \39442 , \39227 , \39441 );
xor \U$39100 ( \39443 , \38965 , \38991 );
xor \U$39101 ( \39444 , \39443 , \39018 );
xor \U$39102 ( \39445 , \39125 , \38748 );
xor \U$39103 ( \39446 , \39445 , \39128 );
and \U$39104 ( \39447 , \39444 , \39446 );
xor \U$39105 ( \39448 , \38844 , \38851 );
xor \U$39106 ( \39449 , \39448 , \38860 );
xor \U$39107 ( \39450 , \38926 , \38931 );
xor \U$39108 ( \39451 , \39449 , \39450 );
xor \U$39109 ( \39452 , \39125 , \38748 );
xor \U$39110 ( \39453 , \39452 , \39128 );
and \U$39111 ( \39454 , \39451 , \39453 );
and \U$39112 ( \39455 , \39444 , \39451 );
or \U$39113 ( \39456 , \39447 , \39454 , \39455 );
and \U$39114 ( \39457 , \39442 , \39456 );
and \U$39115 ( \39458 , \39227 , \39441 );
or \U$39116 ( \39459 , \39457 , \39458 );
xor \U$39117 ( \39460 , \38747 , \38782 );
xor \U$39118 ( \39461 , \39460 , \38866 );
xor \U$39119 ( \39462 , \39459 , \39461 );
xor \U$39120 ( \39463 , \38809 , \38836 );
xor \U$39121 ( \39464 , \39463 , \38863 );
xor \U$39122 ( \39465 , \38694 , \38717 );
xor \U$39123 ( \39466 , \39465 , \38744 );
xor \U$39124 ( \39467 , \39464 , \39466 );
xor \U$39125 ( \39468 , \38884 , \38886 );
xor \U$39126 ( \39469 , \39468 , \38889 );
xor \U$39127 ( \39470 , \39137 , \39144 );
xor \U$39128 ( \39471 , \39469 , \39470 );
and \U$39129 ( \39472 , \39467 , \39471 );
and \U$39130 ( \39473 , \39464 , \39466 );
or \U$39131 ( \39474 , \39472 , \39473 );
and \U$39132 ( \39475 , \39462 , \39474 );
and \U$39133 ( \39476 , \39459 , \39461 );
or \U$39134 ( \39477 , \39475 , \39476 );
xor \U$39135 ( \39478 , \39152 , \39154 );
xor \U$39136 ( \39479 , \39478 , \39169 );
and \U$39137 ( \39480 , \39477 , \39479 );
xor \U$39138 ( \39481 , \38644 , \38646 );
xor \U$39139 ( \39482 , \39481 , \38651 );
xor \U$39140 ( \39483 , \38642 , \38901 );
xor \U$39141 ( \39484 , \39482 , \39483 );
xor \U$39142 ( \39485 , \39152 , \39154 );
xor \U$39143 ( \39486 , \39485 , \39169 );
and \U$39144 ( \39487 , \39484 , \39486 );
and \U$39145 ( \39488 , \39477 , \39484 );
or \U$39146 ( \39489 , \39480 , \39487 , \39488 );
xor \U$39147 ( \39490 , \39179 , \39183 );
xor \U$39148 ( \39491 , \39490 , \39188 );
xor \U$39149 ( \39492 , \39489 , \39491 );
xor \U$39150 ( \39493 , \38906 , \38908 );
xor \U$39151 ( \39494 , \39493 , \39172 );
and \U$39152 ( \39495 , \39492 , \39494 );
and \U$39153 ( \39496 , \39489 , \39491 );
or \U$39154 ( \39497 , \39495 , \39496 );
xor \U$39155 ( \39498 , \39191 , \39192 );
xor \U$39156 ( \39499 , \39498 , \39195 );
and \U$39157 ( \39500 , \39497 , \39499 );
and \U$39158 ( \39501 , \39175 , \39497 );
or \U$39159 ( \39502 , \39197 , \39500 , \39501 );
xor \U$39160 ( \39503 , \39191 , \39192 );
and \U$39161 ( \39504 , \39503 , \39195 );
and \U$39162 ( \39505 , \39191 , \39192 );
or \U$39163 ( \39506 , \39504 , \39505 );
xor \U$39164 ( \39507 , \38311 , \38313 );
xor \U$39165 ( \39508 , \39507 , \38328 );
xor \U$39166 ( \39509 , \39506 , \39508 );
xor \U$39167 ( \39510 , \38610 , \38617 );
xor \U$39168 ( \39511 , \39510 , \38622 );
xor \U$39169 ( \39512 , \39509 , \39511 );
and \U$39170 ( \39513 , \39502 , \39512 );
xor \U$39171 ( \39514 , \39512 , \39502 );
xor \U$39172 ( \39515 , \39332 , \39340 );
xor \U$39173 ( \39516 , \39515 , \39349 );
xor \U$39174 ( \39517 , \39416 , \39423 );
xor \U$39175 ( \39518 , \39517 , \39432 );
and \U$39176 ( \39519 , \39516 , \39518 );
xor \U$39177 ( \39520 , \39389 , \39397 );
xor \U$39178 ( \39521 , \39520 , \39405 );
xor \U$39179 ( \39522 , \39416 , \39423 );
xor \U$39180 ( \39523 , \39522 , \39432 );
and \U$39181 ( \39524 , \39521 , \39523 );
and \U$39182 ( \39525 , \39516 , \39521 );
or \U$39183 ( \39526 , \39519 , \39524 , \39525 );
xor \U$39184 ( \39527 , \39074 , \39082 );
xor \U$39185 ( \39528 , \39527 , \39090 );
xor \U$39186 ( \39529 , \39526 , \39528 );
xor \U$39187 ( \39530 , \39363 , \39371 );
xor \U$39188 ( \39531 , \39530 , \39379 );
xor \U$39189 ( \39532 , \39234 , \39242 );
xor \U$39190 ( \39533 , \39532 , \39251 );
xor \U$39191 ( \39534 , \39531 , \39533 );
xor \U$39192 ( \39535 , \39285 , \39293 );
xor \U$39193 ( \39536 , \39535 , \39301 );
and \U$39194 ( \39537 , \39534 , \39536 );
and \U$39195 ( \39538 , \39531 , \39533 );
or \U$39196 ( \39539 , \39537 , \39538 );
and \U$39197 ( \39540 , \39529 , \39539 );
and \U$39198 ( \39541 , \39526 , \39528 );
or \U$39199 ( \39542 , \39540 , \39541 );
and \U$39200 ( \39543 , \5318 , RI986f598_54);
and \U$39201 ( \39544 , RI986f688_56, \5316 );
nor \U$39202 ( \39545 , \39543 , \39544 );
and \U$39203 ( \39546 , \39545 , \5052 );
not \U$39204 ( \39547 , \39545 );
and \U$39205 ( \39548 , \39547 , \5322 );
nor \U$39206 ( \39549 , \39546 , \39548 );
and \U$39207 ( \39550 , \5881 , RI986e008_8);
and \U$39208 ( \39551 , RI986df18_6, \5879 );
nor \U$39209 ( \39552 , \39550 , \39551 );
and \U$39210 ( \39553 , \39552 , \5594 );
not \U$39211 ( \39554 , \39552 );
and \U$39212 ( \39555 , \39554 , \5885 );
nor \U$39213 ( \39556 , \39553 , \39555 );
xor \U$39214 ( \39557 , \39549 , \39556 );
and \U$39215 ( \39558 , \6453 , RI986de28_4);
and \U$39216 ( \39559 , RI986dd38_2, \6451 );
nor \U$39217 ( \39560 , \39558 , \39559 );
and \U$39218 ( \39561 , \39560 , \6190 );
not \U$39219 ( \39562 , \39560 );
and \U$39220 ( \39563 , \39562 , \6705 );
nor \U$39221 ( \39564 , \39561 , \39563 );
and \U$39222 ( \39565 , \39557 , \39564 );
and \U$39223 ( \39566 , \39549 , \39556 );
or \U$39224 ( \39567 , \39565 , \39566 );
and \U$39225 ( \39568 , \7729 , RI986e2d8_14);
and \U$39226 ( \39569 , RI986e3c8_16, \7727 );
nor \U$39227 ( \39570 , \39568 , \39569 );
and \U$39228 ( \39571 , \39570 , \7480 );
not \U$39229 ( \39572 , \39570 );
and \U$39230 ( \39573 , \39572 , \7733 );
nor \U$39231 ( \39574 , \39571 , \39573 );
xor \U$39232 ( \39575 , \39574 , \8050 );
and \U$39233 ( \39576 , \7079 , RI986e1e8_12);
and \U$39234 ( \39577 , RI986e0f8_10, \7077 );
nor \U$39235 ( \39578 , \39576 , \39577 );
and \U$39236 ( \39579 , \39578 , \6710 );
not \U$39237 ( \39580 , \39578 );
and \U$39238 ( \39581 , \39580 , \6709 );
nor \U$39239 ( \39582 , \39579 , \39581 );
and \U$39240 ( \39583 , \39575 , \39582 );
and \U$39241 ( \39584 , \39574 , \8050 );
or \U$39242 ( \39585 , \39583 , \39584 );
xor \U$39243 ( \39586 , \39567 , \39585 );
not \U$39244 ( \39587 , \4519 );
and \U$39245 ( \39588 , \4710 , RI986f4a8_52);
and \U$39246 ( \39589 , RI986f3b8_50, \4708 );
nor \U$39247 ( \39590 , \39588 , \39589 );
not \U$39248 ( \39591 , \39590 );
or \U$39249 ( \39592 , \39587 , \39591 );
or \U$39250 ( \39593 , \39590 , \4521 );
nand \U$39251 ( \39594 , \39592 , \39593 );
not \U$39252 ( \39595 , \3918 );
and \U$39253 ( \39596 , \3683 , RI986f868_60);
and \U$39254 ( \39597 , RI986f778_58, \3681 );
nor \U$39255 ( \39598 , \39596 , \39597 );
not \U$39256 ( \39599 , \39598 );
or \U$39257 ( \39600 , \39595 , \39599 );
or \U$39258 ( \39601 , \39598 , \3412 );
nand \U$39259 ( \39602 , \39600 , \39601 );
xor \U$39260 ( \39603 , \39594 , \39602 );
and \U$39261 ( \39604 , \4203 , RI986fa48_64);
and \U$39262 ( \39605 , RI986f958_62, \4201 );
nor \U$39263 ( \39606 , \39604 , \39605 );
and \U$39264 ( \39607 , \39606 , \4207 );
not \U$39265 ( \39608 , \39606 );
and \U$39266 ( \39609 , \39608 , \3923 );
nor \U$39267 ( \39610 , \39607 , \39609 );
and \U$39268 ( \39611 , \39603 , \39610 );
and \U$39269 ( \39612 , \39594 , \39602 );
or \U$39270 ( \39613 , \39611 , \39612 );
and \U$39271 ( \39614 , \39586 , \39613 );
and \U$39272 ( \39615 , \39567 , \39585 );
nor \U$39273 ( \39616 , \39614 , \39615 );
and \U$39274 ( \39617 , \2274 , RI986f2c8_48);
and \U$39275 ( \39618 , RI986f1d8_46, \2272 );
nor \U$39276 ( \39619 , \39617 , \39618 );
and \U$39277 ( \39620 , \39619 , \2031 );
not \U$39278 ( \39621 , \39619 );
and \U$39279 ( \39622 , \39621 , \2030 );
nor \U$39280 ( \39623 , \39620 , \39622 );
not \U$39281 ( \39624 , \39623 );
and \U$39282 ( \39625 , \3254 , RI986e788_24);
and \U$39283 ( \39626 , RI986e698_22, \3252 );
nor \U$39284 ( \39627 , \39625 , \39626 );
not \U$39285 ( \39628 , \39627 );
not \U$39286 ( \39629 , \3406 );
and \U$39287 ( \39630 , \39628 , \39629 );
and \U$39288 ( \39631 , \39627 , \3406 );
nor \U$39289 ( \39632 , \39630 , \39631 );
not \U$39290 ( \39633 , \39632 );
and \U$39291 ( \39634 , \39624 , \39633 );
and \U$39292 ( \39635 , \39632 , \39623 );
and \U$39293 ( \39636 , \2464 , RI986e5a8_20);
and \U$39294 ( \39637 , RI986e4b8_18, \2462 );
nor \U$39295 ( \39638 , \39636 , \39637 );
and \U$39296 ( \39639 , \39638 , \2263 );
not \U$39297 ( \39640 , \39638 );
and \U$39298 ( \39641 , \39640 , \2468 );
nor \U$39299 ( \39642 , \39639 , \39641 );
nor \U$39300 ( \39643 , \39635 , \39642 );
nor \U$39301 ( \39644 , \39634 , \39643 );
and \U$39302 ( \39645 , \438 , RI9871578_122);
and \U$39303 ( \39646 , RI9871668_124, \436 );
nor \U$39304 ( \39647 , \39645 , \39646 );
and \U$39305 ( \39648 , \39647 , \443 );
not \U$39306 ( \39649 , \39647 );
and \U$39307 ( \39650 , \39649 , \444 );
nor \U$39308 ( \39651 , \39648 , \39650 );
not \U$39309 ( \39652 , \39651 );
and \U$39310 ( \39653 , \1293 , RI986e968_28);
and \U$39311 ( \39654 , RI986e878_26, \1291 );
nor \U$39312 ( \39655 , \39653 , \39654 );
not \U$39313 ( \39656 , \39655 );
not \U$39314 ( \39657 , \1128 );
and \U$39315 ( \39658 , \39656 , \39657 );
and \U$39316 ( \39659 , \39655 , \1128 );
nor \U$39317 ( \39660 , \39658 , \39659 );
not \U$39318 ( \39661 , \39660 );
and \U$39319 ( \39662 , \39652 , \39661 );
and \U$39320 ( \39663 , \39660 , \39651 );
and \U$39321 ( \39664 , \776 , RI986eb48_32);
and \U$39322 ( \39665 , RI986ea58_30, \774 );
nor \U$39323 ( \39666 , \39664 , \39665 );
and \U$39324 ( \39667 , \39666 , \451 );
not \U$39325 ( \39668 , \39666 );
and \U$39326 ( \39669 , \39668 , \474 );
nor \U$39327 ( \39670 , \39667 , \39669 );
nor \U$39328 ( \39671 , \39663 , \39670 );
nor \U$39329 ( \39672 , \39662 , \39671 );
xor \U$39330 ( \39673 , \39644 , \39672 );
and \U$39331 ( \39674 , \1329 , RI986ef08_40);
and \U$39332 ( \39675 , RI986ee18_38, \1327 );
nor \U$39333 ( \39676 , \39674 , \39675 );
and \U$39334 ( \39677 , \39676 , \1337 );
not \U$39335 ( \39678 , \39676 );
and \U$39336 ( \39679 , \39678 , \1336 );
nor \U$39337 ( \39680 , \39677 , \39679 );
not \U$39338 ( \39681 , \39680 );
and \U$39339 ( \39682 , \1311 , RI986ec38_34);
and \U$39340 ( \39683 , RI986ed28_36, \1309 );
nor \U$39341 ( \39684 , \39682 , \39683 );
and \U$39342 ( \39685 , \39684 , \1315 );
not \U$39343 ( \39686 , \39684 );
and \U$39344 ( \39687 , \39686 , \1458 );
nor \U$39345 ( \39688 , \39685 , \39687 );
not \U$39346 ( \39689 , \39688 );
and \U$39347 ( \39690 , \39681 , \39689 );
and \U$39348 ( \39691 , \39688 , \39680 );
and \U$39349 ( \39692 , \2042 , RI986f0e8_44);
and \U$39350 ( \39693 , RI986eff8_42, \2040 );
nor \U$39351 ( \39694 , \39692 , \39693 );
not \U$39352 ( \39695 , \39694 );
not \U$39353 ( \39696 , \2034 );
and \U$39354 ( \39697 , \39695 , \39696 );
and \U$39355 ( \39698 , \39694 , \2034 );
nor \U$39356 ( \39699 , \39697 , \39698 );
nor \U$39357 ( \39700 , \39691 , \39699 );
nor \U$39358 ( \39701 , \39690 , \39700 );
and \U$39359 ( \39702 , \39673 , \39701 );
and \U$39360 ( \39703 , \39644 , \39672 );
or \U$39361 ( \39704 , \39702 , \39703 );
or \U$39362 ( \39705 , \39616 , \39704 );
not \U$39363 ( \39706 , \39616 );
not \U$39364 ( \39707 , \39704 );
or \U$39365 ( \39708 , \39706 , \39707 );
and \U$39366 ( \39709 , \354 , RI98710c8_112);
and \U$39367 ( \39710 , RI9870d08_104, \352 );
nor \U$39368 ( \39711 , \39709 , \39710 );
not \U$39369 ( \39712 , \39711 );
not \U$39370 ( \39713 , \361 );
and \U$39371 ( \39714 , \39712 , \39713 );
and \U$39372 ( \39715 , \39711 , \345 );
nor \U$39373 ( \39716 , \39714 , \39715 );
nand \U$39374 ( \39717 , RI9870a38_98, RI9871fc8_144);
or \U$39375 ( \39718 , \39716 , \39717 );
not \U$39376 ( \39719 , \39717 );
not \U$39377 ( \39720 , \39716 );
or \U$39378 ( \39721 , \39719 , \39720 );
and \U$39379 ( \39722 , \416 , RI9870ee8_108);
and \U$39380 ( \39723 , RI9870c18_102, \414 );
nor \U$39381 ( \39724 , \39722 , \39723 );
and \U$39382 ( \39725 , \39724 , \422 );
not \U$39383 ( \39726 , \39724 );
and \U$39384 ( \39727 , \39726 , \421 );
nor \U$39385 ( \39728 , \39725 , \39727 );
nand \U$39386 ( \39729 , \39721 , \39728 );
nand \U$39387 ( \39730 , \39718 , \39729 );
or \U$39388 ( \39731 , \39315 , \39308 );
nand \U$39389 ( \39732 , \39731 , \39316 );
xor \U$39390 ( \39733 , \39730 , \39732 );
not \U$39391 ( \39734 , \454 );
and \U$39392 ( \39735 , \465 , RI9871758_126);
and \U$39393 ( \39736 , RI9871848_128, \463 );
nor \U$39394 ( \39737 , \39735 , \39736 );
not \U$39395 ( \39738 , \39737 );
or \U$39396 ( \39739 , \39734 , \39738 );
or \U$39397 ( \39740 , \39737 , \456 );
nand \U$39398 ( \39741 , \39739 , \39740 );
not \U$39399 ( \39742 , \367 );
and \U$39400 ( \39743 , \376 , RI9871398_118);
and \U$39401 ( \39744 , RI9871488_120, \374 );
nor \U$39402 ( \39745 , \39743 , \39744 );
not \U$39403 ( \39746 , \39745 );
or \U$39404 ( \39747 , \39742 , \39746 );
or \U$39405 ( \39748 , \39745 , \367 );
nand \U$39406 ( \39749 , \39747 , \39748 );
xor \U$39407 ( \39750 , \39741 , \39749 );
not \U$39408 ( \39751 , \386 );
and \U$39409 ( \39752 , \395 , RI98712a8_116);
and \U$39410 ( \39753 , RI98711b8_114, \393 );
nor \U$39411 ( \39754 , \39752 , \39753 );
not \U$39412 ( \39755 , \39754 );
or \U$39413 ( \39756 , \39751 , \39755 );
or \U$39414 ( \39757 , \39754 , \386 );
nand \U$39415 ( \39758 , \39756 , \39757 );
and \U$39416 ( \39759 , \39750 , \39758 );
and \U$39417 ( \39760 , \39741 , \39749 );
or \U$39418 ( \39761 , \39759 , \39760 );
and \U$39419 ( \39762 , \39733 , \39761 );
and \U$39420 ( \39763 , \39730 , \39732 );
or \U$39421 ( \39764 , \39762 , \39763 );
nand \U$39422 ( \39765 , \39708 , \39764 );
nand \U$39423 ( \39766 , \39705 , \39765 );
xor \U$39424 ( \39767 , \39542 , \39766 );
xor \U$39425 ( \39768 , \39055 , \7480 );
xor \U$39426 ( \39769 , \39768 , \39063 );
xor \U$39427 ( \39770 , \39211 , \39213 );
xor \U$39428 ( \39771 , \39770 , \39216 );
and \U$39429 ( \39772 , \39769 , \39771 );
xor \U$39430 ( \39773 , \39000 , \39007 );
xor \U$39431 ( \39774 , \39773 , \39015 );
xor \U$39432 ( \39775 , \39199 , \39204 );
xor \U$39433 ( \39776 , \39774 , \39775 );
xor \U$39434 ( \39777 , \39211 , \39213 );
xor \U$39435 ( \39778 , \39777 , \39216 );
and \U$39436 ( \39779 , \39776 , \39778 );
and \U$39437 ( \39780 , \39769 , \39776 );
or \U$39438 ( \39781 , \39772 , \39779 , \39780 );
and \U$39439 ( \39782 , \39767 , \39781 );
and \U$39440 ( \39783 , \39542 , \39766 );
or \U$39441 ( \39784 , \39782 , \39783 );
xor \U$39442 ( \39785 , \38921 , \38923 );
xor \U$39443 ( \39786 , \39785 , \38936 );
xor \U$39444 ( \39787 , \39784 , \39786 );
xor \U$39445 ( \39788 , \39316 , \39323 );
xor \U$39446 ( \39789 , \39788 , \39352 );
xor \U$39447 ( \39790 , \39254 , \39277 );
xor \U$39448 ( \39791 , \39790 , \39304 );
and \U$39449 ( \39792 , \39789 , \39791 );
xor \U$39450 ( \39793 , \39382 , \39408 );
xor \U$39451 ( \39794 , \39793 , \39435 );
xor \U$39452 ( \39795 , \39254 , \39277 );
xor \U$39453 ( \39796 , \39795 , \39304 );
and \U$39454 ( \39797 , \39794 , \39796 );
and \U$39455 ( \39798 , \39789 , \39794 );
or \U$39456 ( \39799 , \39792 , \39797 , \39798 );
xor \U$39457 ( \39800 , \39048 , \39066 );
xor \U$39458 ( \39801 , \39800 , \39093 );
xor \U$39459 ( \39802 , \39799 , \39801 );
xor \U$39460 ( \39803 , \39125 , \38748 );
xor \U$39461 ( \39804 , \39803 , \39128 );
xor \U$39462 ( \39805 , \39444 , \39451 );
xor \U$39463 ( \39806 , \39804 , \39805 );
and \U$39464 ( \39807 , \39802 , \39806 );
and \U$39465 ( \39808 , \39799 , \39801 );
or \U$39466 ( \39809 , \39807 , \39808 );
and \U$39467 ( \39810 , \39787 , \39809 );
and \U$39468 ( \39811 , \39784 , \39786 );
or \U$39469 ( \39812 , \39810 , \39811 );
xor \U$39470 ( \39813 , \38882 , \38892 );
xor \U$39471 ( \39814 , \39813 , \38897 );
xor \U$39472 ( \39815 , \39157 , \39164 );
xor \U$39473 ( \39816 , \39814 , \39815 );
xor \U$39474 ( \39817 , \39812 , \39816 );
xor \U$39475 ( \39818 , \39021 , \39096 );
xor \U$39476 ( \39819 , \39818 , \39131 );
xor \U$39477 ( \39820 , \39464 , \39466 );
xor \U$39478 ( \39821 , \39820 , \39471 );
and \U$39479 ( \39822 , \39819 , \39821 );
xor \U$39480 ( \39823 , \39227 , \39441 );
xor \U$39481 ( \39824 , \39823 , \39456 );
xor \U$39482 ( \39825 , \39464 , \39466 );
xor \U$39483 ( \39826 , \39825 , \39471 );
and \U$39484 ( \39827 , \39824 , \39826 );
and \U$39485 ( \39828 , \39819 , \39824 );
or \U$39486 ( \39829 , \39822 , \39827 , \39828 );
and \U$39487 ( \39830 , \39817 , \39829 );
and \U$39488 ( \39831 , \39812 , \39816 );
or \U$39489 ( \39832 , \39830 , \39831 );
xor \U$39490 ( \39833 , \38939 , \39134 );
xor \U$39491 ( \39834 , \39833 , \39149 );
xor \U$39492 ( \39835 , \39459 , \39461 );
xor \U$39493 ( \39836 , \39835 , \39474 );
and \U$39494 ( \39837 , \39834 , \39836 );
xor \U$39495 ( \39838 , \39832 , \39837 );
xor \U$39496 ( \39839 , \39152 , \39154 );
xor \U$39497 ( \39840 , \39839 , \39169 );
xor \U$39498 ( \39841 , \39477 , \39484 );
xor \U$39499 ( \39842 , \39840 , \39841 );
and \U$39500 ( \39843 , \39838 , \39842 );
and \U$39501 ( \39844 , \39832 , \39837 );
or \U$39502 ( \39845 , \39843 , \39844 );
xor \U$39503 ( \39846 , \39489 , \39491 );
xor \U$39504 ( \39847 , \39846 , \39494 );
and \U$39505 ( \39848 , \39845 , \39847 );
not \U$39506 ( \39849 , \39848 );
xor \U$39507 ( \39850 , \39191 , \39192 );
xor \U$39508 ( \39851 , \39850 , \39195 );
xor \U$39509 ( \39852 , \39175 , \39497 );
xor \U$39510 ( \39853 , \39851 , \39852 );
not \U$39511 ( \39854 , \39853 );
or \U$39512 ( \39855 , \39849 , \39854 );
xor \U$39513 ( \39856 , \39845 , \39847 );
xor \U$39514 ( \39857 , \39832 , \39837 );
xor \U$39515 ( \39858 , \39857 , \39842 );
and \U$39516 ( \39859 , \1329 , RI986e878_26);
and \U$39517 ( \39860 , RI986ef08_40, \1327 );
nor \U$39518 ( \39861 , \39859 , \39860 );
and \U$39519 ( \39862 , \39861 , \1337 );
not \U$39520 ( \39863 , \39861 );
and \U$39521 ( \39864 , \39863 , \1336 );
nor \U$39522 ( \39865 , \39862 , \39864 );
and \U$39523 ( \39866 , \1311 , RI986ee18_38);
and \U$39524 ( \39867 , RI986ec38_34, \1309 );
nor \U$39525 ( \39868 , \39866 , \39867 );
and \U$39526 ( \39869 , \39868 , \1315 );
not \U$39527 ( \39870 , \39868 );
and \U$39528 ( \39871 , \39870 , \1319 );
nor \U$39529 ( \39872 , \39869 , \39871 );
xor \U$39530 ( \39873 , \39865 , \39872 );
and \U$39531 ( \39874 , \2042 , RI986ed28_36);
and \U$39532 ( \39875 , RI986f0e8_44, \2040 );
nor \U$39533 ( \39876 , \39874 , \39875 );
not \U$39534 ( \39877 , \39876 );
not \U$39535 ( \39878 , \2034 );
and \U$39536 ( \39879 , \39877 , \39878 );
and \U$39537 ( \39880 , \39876 , \1462 );
nor \U$39538 ( \39881 , \39879 , \39880 );
and \U$39539 ( \39882 , \39873 , \39881 );
and \U$39540 ( \39883 , \39865 , \39872 );
or \U$39541 ( \39884 , \39882 , \39883 );
and \U$39542 ( \39885 , \3254 , RI986e4b8_18);
and \U$39543 ( \39886 , RI986e788_24, \3252 );
nor \U$39544 ( \39887 , \39885 , \39886 );
not \U$39545 ( \39888 , \39887 );
not \U$39546 ( \39889 , \3406 );
and \U$39547 ( \39890 , \39888 , \39889 );
and \U$39548 ( \39891 , \39887 , \3406 );
nor \U$39549 ( \39892 , \39890 , \39891 );
and \U$39550 ( \39893 , \2274 , RI986eff8_42);
and \U$39551 ( \39894 , RI986f2c8_48, \2272 );
nor \U$39552 ( \39895 , \39893 , \39894 );
and \U$39553 ( \39896 , \39895 , \2031 );
not \U$39554 ( \39897 , \39895 );
and \U$39555 ( \39898 , \39897 , \2030 );
nor \U$39556 ( \39899 , \39896 , \39898 );
xor \U$39557 ( \39900 , \39892 , \39899 );
and \U$39558 ( \39901 , \2464 , RI986f1d8_46);
and \U$39559 ( \39902 , RI986e5a8_20, \2462 );
nor \U$39560 ( \39903 , \39901 , \39902 );
and \U$39561 ( \39904 , \39903 , \2263 );
not \U$39562 ( \39905 , \39903 );
and \U$39563 ( \39906 , \39905 , \2468 );
nor \U$39564 ( \39907 , \39904 , \39906 );
and \U$39565 ( \39908 , \39900 , \39907 );
and \U$39566 ( \39909 , \39892 , \39899 );
or \U$39567 ( \39910 , \39908 , \39909 );
xor \U$39568 ( \39911 , \39884 , \39910 );
and \U$39569 ( \39912 , \1293 , RI986ea58_30);
and \U$39570 ( \39913 , RI986e968_28, \1291 );
nor \U$39571 ( \39914 , \39912 , \39913 );
not \U$39572 ( \39915 , \39914 );
not \U$39573 ( \39916 , \1301 );
and \U$39574 ( \39917 , \39915 , \39916 );
and \U$39575 ( \39918 , \39914 , \1128 );
nor \U$39576 ( \39919 , \39917 , \39918 );
and \U$39577 ( \39920 , \776 , RI9871668_124);
and \U$39578 ( \39921 , RI986eb48_32, \774 );
nor \U$39579 ( \39922 , \39920 , \39921 );
and \U$39580 ( \39923 , \39922 , \451 );
not \U$39581 ( \39924 , \39922 );
and \U$39582 ( \39925 , \39924 , \474 );
nor \U$39583 ( \39926 , \39923 , \39925 );
xor \U$39584 ( \39927 , \39919 , \39926 );
and \U$39585 ( \39928 , \438 , RI9871848_128);
and \U$39586 ( \39929 , RI9871578_122, \436 );
nor \U$39587 ( \39930 , \39928 , \39929 );
and \U$39588 ( \39931 , \39930 , \443 );
not \U$39589 ( \39932 , \39930 );
and \U$39590 ( \39933 , \39932 , \444 );
nor \U$39591 ( \39934 , \39931 , \39933 );
and \U$39592 ( \39935 , \39927 , \39934 );
and \U$39593 ( \39936 , \39919 , \39926 );
or \U$39594 ( \39937 , \39935 , \39936 );
and \U$39595 ( \39938 , \39911 , \39937 );
and \U$39596 ( \39939 , \39884 , \39910 );
nor \U$39597 ( \39940 , \39938 , \39939 );
and \U$39598 ( \39941 , \7079 , RI986dd38_2);
and \U$39599 ( \39942 , RI986e1e8_12, \7077 );
nor \U$39600 ( \39943 , \39941 , \39942 );
and \U$39601 ( \39944 , \39943 , \6709 );
not \U$39602 ( \39945 , \39943 );
and \U$39603 ( \39946 , \39945 , \6710 );
nor \U$39604 ( \39947 , \39944 , \39946 );
nand \U$39605 ( \39948 , RI986e3c8_16, \8486 );
and \U$39606 ( \39949 , \39948 , \8051 );
not \U$39607 ( \39950 , \39948 );
and \U$39608 ( \39951 , \39950 , \8050 );
nor \U$39609 ( \39952 , \39949 , \39951 );
xor \U$39610 ( \39953 , \39947 , \39952 );
and \U$39611 ( \39954 , \7729 , RI986e0f8_10);
and \U$39612 ( \39955 , RI986e2d8_14, \7727 );
nor \U$39613 ( \39956 , \39954 , \39955 );
and \U$39614 ( \39957 , \39956 , \7733 );
not \U$39615 ( \39958 , \39956 );
and \U$39616 ( \39959 , \39958 , \7480 );
nor \U$39617 ( \39960 , \39957 , \39959 );
and \U$39618 ( \39961 , \39953 , \39960 );
and \U$39619 ( \39962 , \39947 , \39952 );
or \U$39620 ( \39963 , \39961 , \39962 );
and \U$39621 ( \39964 , \5318 , RI986f3b8_50);
and \U$39622 ( \39965 , RI986f598_54, \5316 );
nor \U$39623 ( \39966 , \39964 , \39965 );
and \U$39624 ( \39967 , \39966 , \5322 );
not \U$39625 ( \39968 , \39966 );
and \U$39626 ( \39969 , \39968 , \5052 );
nor \U$39627 ( \39970 , \39967 , \39969 );
not \U$39628 ( \39971 , \39970 );
and \U$39629 ( \39972 , \6453 , RI986df18_6);
and \U$39630 ( \39973 , RI986de28_4, \6451 );
nor \U$39631 ( \39974 , \39972 , \39973 );
and \U$39632 ( \39975 , \39974 , \6180 );
not \U$39633 ( \39976 , \39974 );
and \U$39634 ( \39977 , \39976 , \6190 );
nor \U$39635 ( \39978 , \39975 , \39977 );
not \U$39636 ( \39979 , \39978 );
and \U$39637 ( \39980 , \39971 , \39979 );
and \U$39638 ( \39981 , \39978 , \39970 );
and \U$39639 ( \39982 , \5881 , RI986f688_56);
and \U$39640 ( \39983 , RI986e008_8, \5879 );
nor \U$39641 ( \39984 , \39982 , \39983 );
and \U$39642 ( \39985 , \39984 , \5885 );
not \U$39643 ( \39986 , \39984 );
and \U$39644 ( \39987 , \39986 , \5594 );
nor \U$39645 ( \39988 , \39985 , \39987 );
nor \U$39646 ( \39989 , \39981 , \39988 );
nor \U$39647 ( \39990 , \39980 , \39989 );
xor \U$39648 ( \39991 , \39963 , \39990 );
and \U$39649 ( \39992 , \4203 , RI986f778_58);
and \U$39650 ( \39993 , RI986fa48_64, \4201 );
nor \U$39651 ( \39994 , \39992 , \39993 );
and \U$39652 ( \39995 , \39994 , \3923 );
not \U$39653 ( \39996 , \39994 );
and \U$39654 ( \39997 , \39996 , \4207 );
nor \U$39655 ( \39998 , \39995 , \39997 );
and \U$39656 ( \39999 , \3683 , RI986e698_22);
and \U$39657 ( \40000 , RI986f868_60, \3681 );
nor \U$39658 ( \40001 , \39999 , \40000 );
not \U$39659 ( \40002 , \40001 );
not \U$39660 ( \40003 , \3918 );
and \U$39661 ( \40004 , \40002 , \40003 );
and \U$39662 ( \40005 , \40001 , \3918 );
nor \U$39663 ( \40006 , \40004 , \40005 );
xor \U$39664 ( \40007 , \39998 , \40006 );
and \U$39665 ( \40008 , \4710 , RI986f958_62);
and \U$39666 ( \40009 , RI986f4a8_52, \4708 );
nor \U$39667 ( \40010 , \40008 , \40009 );
not \U$39668 ( \40011 , \40010 );
not \U$39669 ( \40012 , \4519 );
and \U$39670 ( \40013 , \40011 , \40012 );
and \U$39671 ( \40014 , \40010 , \4519 );
nor \U$39672 ( \40015 , \40013 , \40014 );
and \U$39673 ( \40016 , \40007 , \40015 );
and \U$39674 ( \40017 , \39998 , \40006 );
or \U$39675 ( \40018 , \40016 , \40017 );
and \U$39676 ( \40019 , \39991 , \40018 );
and \U$39677 ( \40020 , \39963 , \39990 );
nor \U$39678 ( \40021 , \40019 , \40020 );
xor \U$39679 ( \40022 , \39940 , \40021 );
not \U$39680 ( \40023 , \39716 );
not \U$39681 ( \40024 , \39728 );
or \U$39682 ( \40025 , \40023 , \40024 );
or \U$39683 ( \40026 , \39716 , \39728 );
nand \U$39684 ( \40027 , \40025 , \40026 );
not \U$39685 ( \40028 , \40027 );
not \U$39686 ( \40029 , \39717 );
and \U$39687 ( \40030 , \40028 , \40029 );
and \U$39688 ( \40031 , \40027 , \39717 );
nor \U$39689 ( \40032 , \40030 , \40031 );
and \U$39690 ( \40033 , \395 , RI9870d08_104);
and \U$39691 ( \40034 , RI98712a8_116, \393 );
nor \U$39692 ( \40035 , \40033 , \40034 );
not \U$39693 ( \40036 , \40035 );
not \U$39694 ( \40037 , \487 );
and \U$39695 ( \40038 , \40036 , \40037 );
and \U$39696 ( \40039 , \40035 , \386 );
nor \U$39697 ( \40040 , \40038 , \40039 );
and \U$39698 ( \40041 , \465 , RI9871488_120);
and \U$39699 ( \40042 , RI9871758_126, \463 );
nor \U$39700 ( \40043 , \40041 , \40042 );
not \U$39701 ( \40044 , \40043 );
not \U$39702 ( \40045 , \456 );
and \U$39703 ( \40046 , \40044 , \40045 );
and \U$39704 ( \40047 , \40043 , \454 );
nor \U$39705 ( \40048 , \40046 , \40047 );
xor \U$39706 ( \40049 , \40040 , \40048 );
and \U$39707 ( \40050 , \376 , RI98711b8_114);
and \U$39708 ( \40051 , RI9871398_118, \374 );
nor \U$39709 ( \40052 , \40050 , \40051 );
not \U$39710 ( \40053 , \40052 );
not \U$39711 ( \40054 , \367 );
and \U$39712 ( \40055 , \40053 , \40054 );
and \U$39713 ( \40056 , \40052 , \365 );
nor \U$39714 ( \40057 , \40055 , \40056 );
and \U$39715 ( \40058 , \40049 , \40057 );
and \U$39716 ( \40059 , \40040 , \40048 );
or \U$39717 ( \40060 , \40058 , \40059 );
or \U$39718 ( \40061 , \40032 , \40060 );
not \U$39719 ( \40062 , \40060 );
not \U$39720 ( \40063 , \40032 );
or \U$39721 ( \40064 , \40062 , \40063 );
and \U$39722 ( \40065 , \416 , RI9870a38_98);
and \U$39723 ( \40066 , RI9870ee8_108, \414 );
nor \U$39724 ( \40067 , \40065 , \40066 );
and \U$39725 ( \40068 , \40067 , \421 );
not \U$39726 ( \40069 , \40067 );
and \U$39727 ( \40070 , \40069 , \422 );
nor \U$39728 ( \40071 , \40068 , \40070 );
nand \U$39729 ( \40072 , RI9870df8_106, RI9871fc8_144);
or \U$39730 ( \40073 , \40071 , \40072 );
not \U$39731 ( \40074 , \40072 );
not \U$39732 ( \40075 , \40071 );
or \U$39733 ( \40076 , \40074 , \40075 );
not \U$39734 ( \40077 , \361 );
and \U$39735 ( \40078 , \354 , RI9870c18_102);
and \U$39736 ( \40079 , RI98710c8_112, \352 );
nor \U$39737 ( \40080 , \40078 , \40079 );
not \U$39738 ( \40081 , \40080 );
or \U$39739 ( \40082 , \40077 , \40081 );
or \U$39740 ( \40083 , \40080 , \361 );
nand \U$39741 ( \40084 , \40082 , \40083 );
nand \U$39742 ( \40085 , \40076 , \40084 );
nand \U$39743 ( \40086 , \40073 , \40085 );
nand \U$39744 ( \40087 , \40064 , \40086 );
nand \U$39745 ( \40088 , \40061 , \40087 );
and \U$39746 ( \40089 , \40022 , \40088 );
and \U$39747 ( \40090 , \39940 , \40021 );
or \U$39748 ( \40091 , \40089 , \40090 );
not \U$39749 ( \40092 , \40091 );
xor \U$39750 ( \40093 , \39730 , \39732 );
xor \U$39751 ( \40094 , \40093 , \39761 );
xor \U$39752 ( \40095 , \39531 , \39533 );
xor \U$39753 ( \40096 , \40095 , \39536 );
and \U$39754 ( \40097 , \40094 , \40096 );
xor \U$39755 ( \40098 , \39416 , \39423 );
xor \U$39756 ( \40099 , \40098 , \39432 );
xor \U$39757 ( \40100 , \39516 , \39521 );
xor \U$39758 ( \40101 , \40099 , \40100 );
xor \U$39759 ( \40102 , \39531 , \39533 );
xor \U$39760 ( \40103 , \40102 , \39536 );
and \U$39761 ( \40104 , \40101 , \40103 );
and \U$39762 ( \40105 , \40094 , \40101 );
or \U$39763 ( \40106 , \40097 , \40104 , \40105 );
not \U$39764 ( \40107 , \40106 );
or \U$39765 ( \40108 , \40092 , \40107 );
or \U$39766 ( \40109 , \40106 , \40091 );
not \U$39767 ( \40110 , \39680 );
xor \U$39768 ( \40111 , \39688 , \39699 );
not \U$39769 ( \40112 , \40111 );
or \U$39770 ( \40113 , \40110 , \40112 );
or \U$39771 ( \40114 , \40111 , \39680 );
nand \U$39772 ( \40115 , \40113 , \40114 );
xor \U$39773 ( \40116 , \39741 , \39749 );
xor \U$39774 ( \40117 , \40116 , \39758 );
xor \U$39775 ( \40118 , \40115 , \40117 );
not \U$39776 ( \40119 , \39651 );
xor \U$39777 ( \40120 , \39670 , \39660 );
not \U$39778 ( \40121 , \40120 );
or \U$39779 ( \40122 , \40119 , \40121 );
or \U$39780 ( \40123 , \40120 , \39651 );
nand \U$39781 ( \40124 , \40122 , \40123 );
and \U$39782 ( \40125 , \40118 , \40124 );
and \U$39783 ( \40126 , \40115 , \40117 );
or \U$39784 ( \40127 , \40125 , \40126 );
xor \U$39785 ( \40128 , \39261 , \39266 );
xor \U$39786 ( \40129 , \40128 , \39274 );
xor \U$39787 ( \40130 , \40127 , \40129 );
not \U$39788 ( \40131 , \39623 );
xor \U$39789 ( \40132 , \39642 , \39632 );
not \U$39790 ( \40133 , \40132 );
or \U$39791 ( \40134 , \40131 , \40133 );
or \U$39792 ( \40135 , \40132 , \39623 );
nand \U$39793 ( \40136 , \40134 , \40135 );
xor \U$39794 ( \40137 , \39594 , \39602 );
xor \U$39795 ( \40138 , \40137 , \39610 );
and \U$39796 ( \40139 , \40136 , \40138 );
xor \U$39797 ( \40140 , \39549 , \39556 );
xor \U$39798 ( \40141 , \40140 , \39564 );
xor \U$39799 ( \40142 , \39594 , \39602 );
xor \U$39800 ( \40143 , \40142 , \39610 );
and \U$39801 ( \40144 , \40141 , \40143 );
and \U$39802 ( \40145 , \40136 , \40141 );
or \U$39803 ( \40146 , \40139 , \40144 , \40145 );
and \U$39804 ( \40147 , \40130 , \40146 );
and \U$39805 ( \40148 , \40127 , \40129 );
or \U$39806 ( \40149 , \40147 , \40148 );
nand \U$39807 ( \40150 , \40109 , \40149 );
nand \U$39808 ( \40151 , \40108 , \40150 );
xor \U$39809 ( \40152 , \39209 , \39219 );
xor \U$39810 ( \40153 , \40152 , \39224 );
xor \U$39811 ( \40154 , \40151 , \40153 );
xor \U$39812 ( \40155 , \39254 , \39277 );
xor \U$39813 ( \40156 , \40155 , \39304 );
xor \U$39814 ( \40157 , \39789 , \39794 );
xor \U$39815 ( \40158 , \40156 , \40157 );
xor \U$39816 ( \40159 , \39526 , \39528 );
xor \U$39817 ( \40160 , \40159 , \39539 );
and \U$39818 ( \40161 , \40158 , \40160 );
xor \U$39819 ( \40162 , \39211 , \39213 );
xor \U$39820 ( \40163 , \40162 , \39216 );
xor \U$39821 ( \40164 , \39769 , \39776 );
xor \U$39822 ( \40165 , \40163 , \40164 );
xor \U$39823 ( \40166 , \39526 , \39528 );
xor \U$39824 ( \40167 , \40166 , \39539 );
and \U$39825 ( \40168 , \40165 , \40167 );
and \U$39826 ( \40169 , \40158 , \40165 );
or \U$39827 ( \40170 , \40161 , \40168 , \40169 );
and \U$39828 ( \40171 , \40154 , \40170 );
and \U$39829 ( \40172 , \40151 , \40153 );
or \U$39830 ( \40173 , \40171 , \40172 );
xor \U$39831 ( \40174 , \39307 , \39355 );
xor \U$39832 ( \40175 , \40174 , \39438 );
xor \U$39833 ( \40176 , \39542 , \39766 );
xor \U$39834 ( \40177 , \40176 , \39781 );
and \U$39835 ( \40178 , \40175 , \40177 );
xor \U$39836 ( \40179 , \39799 , \39801 );
xor \U$39837 ( \40180 , \40179 , \39806 );
xor \U$39838 ( \40181 , \39542 , \39766 );
xor \U$39839 ( \40182 , \40181 , \39781 );
and \U$39840 ( \40183 , \40180 , \40182 );
and \U$39841 ( \40184 , \40175 , \40180 );
or \U$39842 ( \40185 , \40178 , \40183 , \40184 );
xor \U$39843 ( \40186 , \40173 , \40185 );
xor \U$39844 ( \40187 , \39464 , \39466 );
xor \U$39845 ( \40188 , \40187 , \39471 );
xor \U$39846 ( \40189 , \39819 , \39824 );
xor \U$39847 ( \40190 , \40188 , \40189 );
and \U$39848 ( \40191 , \40186 , \40190 );
and \U$39849 ( \40192 , \40173 , \40185 );
or \U$39850 ( \40193 , \40191 , \40192 );
xor \U$39851 ( \40194 , \39834 , \39836 );
xor \U$39852 ( \40195 , \40193 , \40194 );
xor \U$39853 ( \40196 , \39812 , \39816 );
xor \U$39854 ( \40197 , \40196 , \39829 );
and \U$39855 ( \40198 , \40195 , \40197 );
and \U$39856 ( \40199 , \40193 , \40194 );
or \U$39857 ( \40200 , \40198 , \40199 );
and \U$39858 ( \40201 , \39858 , \40200 );
and \U$39859 ( \40202 , \39856 , \40201 );
xor \U$39860 ( \40203 , \40201 , \39856 );
xor \U$39861 ( \40204 , \39858 , \40200 );
not \U$39862 ( \40205 , \40204 );
xor \U$39863 ( \40206 , \39940 , \40021 );
xor \U$39864 ( \40207 , \40206 , \40088 );
xor \U$39865 ( \40208 , \40127 , \40129 );
xor \U$39866 ( \40209 , \40208 , \40146 );
and \U$39867 ( \40210 , \40207 , \40209 );
xor \U$39868 ( \40211 , \39531 , \39533 );
xor \U$39869 ( \40212 , \40211 , \39536 );
xor \U$39870 ( \40213 , \40094 , \40101 );
xor \U$39871 ( \40214 , \40212 , \40213 );
xor \U$39872 ( \40215 , \40127 , \40129 );
xor \U$39873 ( \40216 , \40215 , \40146 );
and \U$39874 ( \40217 , \40214 , \40216 );
and \U$39875 ( \40218 , \40207 , \40214 );
or \U$39876 ( \40219 , \40210 , \40217 , \40218 );
not \U$39877 ( \40220 , \40219 );
xor \U$39878 ( \40221 , \39567 , \39585 );
xor \U$39879 ( \40222 , \40221 , \39613 );
xor \U$39880 ( \40223 , \39644 , \39672 );
xor \U$39881 ( \40224 , \40223 , \39701 );
not \U$39882 ( \40225 , \40224 );
and \U$39883 ( \40226 , \40222 , \40225 );
not \U$39884 ( \40227 , \40222 );
not \U$39885 ( \40228 , \40225 );
and \U$39886 ( \40229 , \40227 , \40228 );
not \U$39887 ( \40230 , \40086 );
not \U$39888 ( \40231 , \40060 );
or \U$39889 ( \40232 , \40230 , \40231 );
or \U$39890 ( \40233 , \40060 , \40086 );
nand \U$39891 ( \40234 , \40232 , \40233 );
not \U$39892 ( \40235 , \40234 );
not \U$39893 ( \40236 , \40032 );
and \U$39894 ( \40237 , \40235 , \40236 );
and \U$39895 ( \40238 , \40234 , \40032 );
nor \U$39896 ( \40239 , \40237 , \40238 );
xor \U$39897 ( \40240 , \39963 , \39990 );
xor \U$39898 ( \40241 , \40240 , \40018 );
xor \U$39899 ( \40242 , \40239 , \40241 );
xor \U$39900 ( \40243 , \39884 , \39910 );
xor \U$39901 ( \40244 , \40243 , \39937 );
and \U$39902 ( \40245 , \40242 , \40244 );
and \U$39903 ( \40246 , \40239 , \40241 );
or \U$39904 ( \40247 , \40245 , \40246 );
nor \U$39905 ( \40248 , \40229 , \40247 );
nor \U$39906 ( \40249 , \40226 , \40248 );
or \U$39907 ( \40250 , \40220 , \40249 );
not \U$39908 ( \40251 , \40249 );
not \U$39909 ( \40252 , \40220 );
or \U$39910 ( \40253 , \40251 , \40252 );
xor \U$39911 ( \40254 , \40040 , \40048 );
xor \U$39912 ( \40255 , \40254 , \40057 );
xor \U$39913 ( \40256 , \39919 , \39926 );
xor \U$39914 ( \40257 , \40256 , \39934 );
xor \U$39915 ( \40258 , \40255 , \40257 );
not \U$39916 ( \40259 , \40071 );
not \U$39917 ( \40260 , \40084 );
or \U$39918 ( \40261 , \40259 , \40260 );
or \U$39919 ( \40262 , \40071 , \40084 );
nand \U$39920 ( \40263 , \40261 , \40262 );
not \U$39921 ( \40264 , \40263 );
not \U$39922 ( \40265 , \40072 );
and \U$39923 ( \40266 , \40264 , \40265 );
and \U$39924 ( \40267 , \40263 , \40072 );
nor \U$39925 ( \40268 , \40266 , \40267 );
and \U$39926 ( \40269 , \40258 , \40268 );
and \U$39927 ( \40270 , \40255 , \40257 );
nor \U$39928 ( \40271 , \40269 , \40270 );
not \U$39929 ( \40272 , \39970 );
xor \U$39930 ( \40273 , \39988 , \39978 );
not \U$39931 ( \40274 , \40273 );
or \U$39932 ( \40275 , \40272 , \40274 );
or \U$39933 ( \40276 , \40273 , \39970 );
nand \U$39934 ( \40277 , \40275 , \40276 );
not \U$39935 ( \40278 , \40277 );
xor \U$39936 ( \40279 , \39947 , \39952 );
xor \U$39937 ( \40280 , \40279 , \39960 );
nor \U$39938 ( \40281 , \40278 , \40280 );
xor \U$39939 ( \40282 , \40271 , \40281 );
xor \U$39940 ( \40283 , \39865 , \39872 );
xor \U$39941 ( \40284 , \40283 , \39881 );
xor \U$39942 ( \40285 , \39892 , \39899 );
xor \U$39943 ( \40286 , \40285 , \39907 );
xor \U$39944 ( \40287 , \40284 , \40286 );
xor \U$39945 ( \40288 , \39998 , \40006 );
xor \U$39946 ( \40289 , \40288 , \40015 );
and \U$39947 ( \40290 , \40287 , \40289 );
and \U$39948 ( \40291 , \40284 , \40286 );
nor \U$39949 ( \40292 , \40290 , \40291 );
and \U$39950 ( \40293 , \40282 , \40292 );
and \U$39951 ( \40294 , \40271 , \40281 );
or \U$39952 ( \40295 , \40293 , \40294 );
and \U$39953 ( \40296 , \465 , RI9871398_118);
and \U$39954 ( \40297 , RI9871488_120, \463 );
nor \U$39955 ( \40298 , \40296 , \40297 );
not \U$39956 ( \40299 , \40298 );
not \U$39957 ( \40300 , \454 );
and \U$39958 ( \40301 , \40299 , \40300 );
and \U$39959 ( \40302 , \40298 , \454 );
nor \U$39960 ( \40303 , \40301 , \40302 );
and \U$39961 ( \40304 , \438 , RI9871758_126);
and \U$39962 ( \40305 , RI9871848_128, \436 );
nor \U$39963 ( \40306 , \40304 , \40305 );
and \U$39964 ( \40307 , \40306 , \443 );
not \U$39965 ( \40308 , \40306 );
and \U$39966 ( \40309 , \40308 , \444 );
nor \U$39967 ( \40310 , \40307 , \40309 );
xor \U$39968 ( \40311 , \40303 , \40310 );
and \U$39969 ( \40312 , \376 , RI98712a8_116);
and \U$39970 ( \40313 , RI98711b8_114, \374 );
nor \U$39971 ( \40314 , \40312 , \40313 );
not \U$39972 ( \40315 , \40314 );
not \U$39973 ( \40316 , \365 );
and \U$39974 ( \40317 , \40315 , \40316 );
and \U$39975 ( \40318 , \40314 , \365 );
nor \U$39976 ( \40319 , \40317 , \40318 );
and \U$39977 ( \40320 , \40311 , \40319 );
and \U$39978 ( \40321 , \40303 , \40310 );
nor \U$39979 ( \40322 , \40320 , \40321 );
and \U$39980 ( \40323 , \395 , RI98710c8_112);
and \U$39981 ( \40324 , RI9870d08_104, \393 );
nor \U$39982 ( \40325 , \40323 , \40324 );
not \U$39983 ( \40326 , \40325 );
not \U$39984 ( \40327 , \487 );
and \U$39985 ( \40328 , \40326 , \40327 );
and \U$39986 ( \40329 , \40325 , \487 );
nor \U$39987 ( \40330 , \40328 , \40329 );
and \U$39988 ( \40331 , \354 , RI9870ee8_108);
and \U$39989 ( \40332 , RI9870c18_102, \352 );
nor \U$39990 ( \40333 , \40331 , \40332 );
not \U$39991 ( \40334 , \40333 );
not \U$39992 ( \40335 , \361 );
and \U$39993 ( \40336 , \40334 , \40335 );
and \U$39994 ( \40337 , \40333 , \361 );
nor \U$39995 ( \40338 , \40336 , \40337 );
xor \U$39996 ( \40339 , \40330 , \40338 );
and \U$39997 ( \40340 , \416 , RI9870df8_106);
and \U$39998 ( \40341 , RI9870a38_98, \414 );
nor \U$39999 ( \40342 , \40340 , \40341 );
and \U$40000 ( \40343 , \40342 , \421 );
not \U$40001 ( \40344 , \40342 );
and \U$40002 ( \40345 , \40344 , \422 );
nor \U$40003 ( \40346 , \40343 , \40345 );
and \U$40004 ( \40347 , \40339 , \40346 );
and \U$40005 ( \40348 , \40330 , \40338 );
nor \U$40006 ( \40349 , \40347 , \40348 );
nor \U$40007 ( \40350 , \40322 , \40349 );
not \U$40008 ( \40351 , \40350 );
not \U$40009 ( \40352 , \40351 );
not \U$40010 ( \40353 , \1301 );
and \U$40011 ( \40354 , \1293 , RI986eb48_32);
and \U$40012 ( \40355 , RI986ea58_30, \1291 );
nor \U$40013 ( \40356 , \40354 , \40355 );
not \U$40014 ( \40357 , \40356 );
or \U$40015 ( \40358 , \40353 , \40357 );
or \U$40016 ( \40359 , \40356 , \1301 );
nand \U$40017 ( \40360 , \40358 , \40359 );
and \U$40018 ( \40361 , \1329 , RI986e968_28);
and \U$40019 ( \40362 , RI986e878_26, \1327 );
nor \U$40020 ( \40363 , \40361 , \40362 );
and \U$40021 ( \40364 , \40363 , \1336 );
not \U$40022 ( \40365 , \40363 );
and \U$40023 ( \40366 , \40365 , \1337 );
nor \U$40024 ( \40367 , \40364 , \40366 );
xor \U$40025 ( \40368 , \40360 , \40367 );
and \U$40026 ( \40369 , \776 , RI9871578_122);
and \U$40027 ( \40370 , RI9871668_124, \774 );
nor \U$40028 ( \40371 , \40369 , \40370 );
and \U$40029 ( \40372 , \40371 , \474 );
not \U$40030 ( \40373 , \40371 );
and \U$40031 ( \40374 , \40373 , \451 );
nor \U$40032 ( \40375 , \40372 , \40374 );
and \U$40033 ( \40376 , \40368 , \40375 );
and \U$40034 ( \40377 , \40360 , \40367 );
nor \U$40035 ( \40378 , \40376 , \40377 );
and \U$40036 ( \40379 , \1311 , RI986ef08_40);
and \U$40037 ( \40380 , RI986ee18_38, \1309 );
nor \U$40038 ( \40381 , \40379 , \40380 );
and \U$40039 ( \40382 , \40381 , \1315 );
not \U$40040 ( \40383 , \40381 );
and \U$40041 ( \40384 , \40383 , \1458 );
nor \U$40042 ( \40385 , \40382 , \40384 );
not \U$40043 ( \40386 , \40385 );
and \U$40044 ( \40387 , \2042 , RI986ec38_34);
and \U$40045 ( \40388 , RI986ed28_36, \2040 );
nor \U$40046 ( \40389 , \40387 , \40388 );
not \U$40047 ( \40390 , \40389 );
not \U$40048 ( \40391 , \1462 );
and \U$40049 ( \40392 , \40390 , \40391 );
and \U$40050 ( \40393 , \40389 , \1462 );
nor \U$40051 ( \40394 , \40392 , \40393 );
not \U$40052 ( \40395 , \40394 );
and \U$40053 ( \40396 , \40386 , \40395 );
and \U$40054 ( \40397 , \40394 , \40385 );
and \U$40055 ( \40398 , \2274 , RI986f0e8_44);
and \U$40056 ( \40399 , RI986eff8_42, \2272 );
nor \U$40057 ( \40400 , \40398 , \40399 );
and \U$40058 ( \40401 , \40400 , \2031 );
not \U$40059 ( \40402 , \40400 );
and \U$40060 ( \40403 , \40402 , \2030 );
nor \U$40061 ( \40404 , \40401 , \40403 );
nor \U$40062 ( \40405 , \40397 , \40404 );
nor \U$40063 ( \40406 , \40396 , \40405 );
xor \U$40064 ( \40407 , \40378 , \40406 );
and \U$40065 ( \40408 , \2464 , RI986f2c8_48);
and \U$40066 ( \40409 , RI986f1d8_46, \2462 );
nor \U$40067 ( \40410 , \40408 , \40409 );
and \U$40068 ( \40411 , \40410 , \2263 );
not \U$40069 ( \40412 , \40410 );
and \U$40070 ( \40413 , \40412 , \2468 );
nor \U$40071 ( \40414 , \40411 , \40413 );
not \U$40072 ( \40415 , \40414 );
and \U$40073 ( \40416 , \3254 , RI986e5a8_20);
and \U$40074 ( \40417 , RI986e4b8_18, \3252 );
nor \U$40075 ( \40418 , \40416 , \40417 );
not \U$40076 ( \40419 , \40418 );
not \U$40077 ( \40420 , \2935 );
and \U$40078 ( \40421 , \40419 , \40420 );
and \U$40079 ( \40422 , \40418 , \2935 );
nor \U$40080 ( \40423 , \40421 , \40422 );
not \U$40081 ( \40424 , \40423 );
and \U$40082 ( \40425 , \40415 , \40424 );
and \U$40083 ( \40426 , \40423 , \40414 );
and \U$40084 ( \40427 , \3683 , RI986e788_24);
and \U$40085 ( \40428 , RI986e698_22, \3681 );
nor \U$40086 ( \40429 , \40427 , \40428 );
not \U$40087 ( \40430 , \40429 );
not \U$40088 ( \40431 , \3918 );
and \U$40089 ( \40432 , \40430 , \40431 );
and \U$40090 ( \40433 , \40429 , \3412 );
nor \U$40091 ( \40434 , \40432 , \40433 );
nor \U$40092 ( \40435 , \40426 , \40434 );
nor \U$40093 ( \40436 , \40425 , \40435 );
and \U$40094 ( \40437 , \40407 , \40436 );
and \U$40095 ( \40438 , \40378 , \40406 );
nor \U$40096 ( \40439 , \40437 , \40438 );
not \U$40097 ( \40440 , \40439 );
or \U$40098 ( \40441 , \40352 , \40440 );
or \U$40099 ( \40442 , \40439 , \40351 );
and \U$40100 ( \40443 , \7729 , RI986e1e8_12);
and \U$40101 ( \40444 , RI986e0f8_10, \7727 );
nor \U$40102 ( \40445 , \40443 , \40444 );
and \U$40103 ( \40446 , \40445 , \7733 );
not \U$40104 ( \40447 , \40445 );
and \U$40105 ( \40448 , \40447 , \7480 );
nor \U$40106 ( \40449 , \40446 , \40448 );
not \U$40107 ( \40450 , \40449 );
not \U$40108 ( \40451 , \8836 );
and \U$40109 ( \40452 , \40450 , \40451 );
and \U$40110 ( \40453 , \40449 , \8836 );
and \U$40111 ( \40454 , \8486 , RI986e2d8_14);
and \U$40112 ( \40455 , RI986e3c8_16, \8484 );
nor \U$40113 ( \40456 , \40454 , \40455 );
and \U$40114 ( \40457 , \40456 , \8051 );
not \U$40115 ( \40458 , \40456 );
and \U$40116 ( \40459 , \40458 , \8050 );
nor \U$40117 ( \40460 , \40457 , \40459 );
nor \U$40118 ( \40461 , \40453 , \40460 );
nor \U$40119 ( \40462 , \40452 , \40461 );
and \U$40120 ( \40463 , \5881 , RI986f598_54);
and \U$40121 ( \40464 , RI986f688_56, \5879 );
nor \U$40122 ( \40465 , \40463 , \40464 );
and \U$40123 ( \40466 , \40465 , \5885 );
not \U$40124 ( \40467 , \40465 );
and \U$40125 ( \40468 , \40467 , \5594 );
nor \U$40126 ( \40469 , \40466 , \40468 );
not \U$40127 ( \40470 , \40469 );
and \U$40128 ( \40471 , \6453 , RI986e008_8);
and \U$40129 ( \40472 , RI986df18_6, \6451 );
nor \U$40130 ( \40473 , \40471 , \40472 );
and \U$40131 ( \40474 , \40473 , \6180 );
not \U$40132 ( \40475 , \40473 );
and \U$40133 ( \40476 , \40475 , \6190 );
nor \U$40134 ( \40477 , \40474 , \40476 );
not \U$40135 ( \40478 , \40477 );
and \U$40136 ( \40479 , \40470 , \40478 );
and \U$40137 ( \40480 , \40477 , \40469 );
and \U$40138 ( \40481 , \7079 , RI986de28_4);
and \U$40139 ( \40482 , RI986dd38_2, \7077 );
nor \U$40140 ( \40483 , \40481 , \40482 );
and \U$40141 ( \40484 , \40483 , \6709 );
not \U$40142 ( \40485 , \40483 );
and \U$40143 ( \40486 , \40485 , \6710 );
nor \U$40144 ( \40487 , \40484 , \40486 );
nor \U$40145 ( \40488 , \40480 , \40487 );
nor \U$40146 ( \40489 , \40479 , \40488 );
xor \U$40147 ( \40490 , \40462 , \40489 );
not \U$40148 ( \40491 , \4519 );
and \U$40149 ( \40492 , \4710 , RI986fa48_64);
and \U$40150 ( \40493 , RI986f958_62, \4708 );
nor \U$40151 ( \40494 , \40492 , \40493 );
not \U$40152 ( \40495 , \40494 );
or \U$40153 ( \40496 , \40491 , \40495 );
or \U$40154 ( \40497 , \40494 , \4521 );
nand \U$40155 ( \40498 , \40496 , \40497 );
and \U$40156 ( \40499 , \5318 , RI986f4a8_52);
and \U$40157 ( \40500 , RI986f3b8_50, \5316 );
nor \U$40158 ( \40501 , \40499 , \40500 );
and \U$40159 ( \40502 , \40501 , \5052 );
not \U$40160 ( \40503 , \40501 );
and \U$40161 ( \40504 , \40503 , \5322 );
nor \U$40162 ( \40505 , \40502 , \40504 );
xor \U$40163 ( \40506 , \40498 , \40505 );
and \U$40164 ( \40507 , \4203 , RI986f868_60);
and \U$40165 ( \40508 , RI986f778_58, \4201 );
nor \U$40166 ( \40509 , \40507 , \40508 );
and \U$40167 ( \40510 , \40509 , \4207 );
not \U$40168 ( \40511 , \40509 );
and \U$40169 ( \40512 , \40511 , \3922 );
nor \U$40170 ( \40513 , \40510 , \40512 );
and \U$40171 ( \40514 , \40506 , \40513 );
and \U$40172 ( \40515 , \40498 , \40505 );
nor \U$40173 ( \40516 , \40514 , \40515 );
and \U$40174 ( \40517 , \40490 , \40516 );
and \U$40175 ( \40518 , \40462 , \40489 );
nor \U$40176 ( \40519 , \40517 , \40518 );
nand \U$40177 ( \40520 , \40442 , \40519 );
nand \U$40178 ( \40521 , \40441 , \40520 );
xor \U$40179 ( \40522 , \40295 , \40521 );
xor \U$40180 ( \40523 , \39574 , \8050 );
xor \U$40181 ( \40524 , \40523 , \39582 );
xor \U$40182 ( \40525 , \40115 , \40117 );
xor \U$40183 ( \40526 , \40525 , \40124 );
and \U$40184 ( \40527 , \40524 , \40526 );
xor \U$40185 ( \40528 , \39594 , \39602 );
xor \U$40186 ( \40529 , \40528 , \39610 );
xor \U$40187 ( \40530 , \40136 , \40141 );
xor \U$40188 ( \40531 , \40529 , \40530 );
xor \U$40189 ( \40532 , \40115 , \40117 );
xor \U$40190 ( \40533 , \40532 , \40124 );
and \U$40191 ( \40534 , \40531 , \40533 );
and \U$40192 ( \40535 , \40524 , \40531 );
or \U$40193 ( \40536 , \40527 , \40534 , \40535 );
and \U$40194 ( \40537 , \40522 , \40536 );
and \U$40195 ( \40538 , \40295 , \40521 );
or \U$40196 ( \40539 , \40537 , \40538 );
nand \U$40197 ( \40540 , \40253 , \40539 );
nand \U$40198 ( \40541 , \40250 , \40540 );
xnor \U$40199 ( \40542 , \40091 , \40149 );
not \U$40200 ( \40543 , \40542 );
not \U$40201 ( \40544 , \40106 );
and \U$40202 ( \40545 , \40543 , \40544 );
and \U$40203 ( \40546 , \40542 , \40106 );
nor \U$40204 ( \40547 , \40545 , \40546 );
xnor \U$40205 ( \40548 , \39616 , \39704 );
not \U$40206 ( \40549 , \40548 );
not \U$40207 ( \40550 , \39764 );
and \U$40208 ( \40551 , \40549 , \40550 );
and \U$40209 ( \40552 , \40548 , \39764 );
nor \U$40210 ( \40553 , \40551 , \40552 );
or \U$40211 ( \40554 , \40547 , \40553 );
not \U$40212 ( \40555 , \40553 );
not \U$40213 ( \40556 , \40547 );
or \U$40214 ( \40557 , \40555 , \40556 );
xor \U$40215 ( \40558 , \39526 , \39528 );
xor \U$40216 ( \40559 , \40558 , \39539 );
xor \U$40217 ( \40560 , \40158 , \40165 );
xor \U$40218 ( \40561 , \40559 , \40560 );
nand \U$40219 ( \40562 , \40557 , \40561 );
nand \U$40220 ( \40563 , \40554 , \40562 );
xor \U$40221 ( \40564 , \40541 , \40563 );
xor \U$40222 ( \40565 , \39542 , \39766 );
xor \U$40223 ( \40566 , \40565 , \39781 );
xor \U$40224 ( \40567 , \40175 , \40180 );
xor \U$40225 ( \40568 , \40566 , \40567 );
and \U$40226 ( \40569 , \40564 , \40568 );
and \U$40227 ( \40570 , \40541 , \40563 );
or \U$40228 ( \40571 , \40569 , \40570 );
xor \U$40229 ( \40572 , \39784 , \39786 );
xor \U$40230 ( \40573 , \40572 , \39809 );
xor \U$40231 ( \40574 , \40571 , \40573 );
xor \U$40232 ( \40575 , \40173 , \40185 );
xor \U$40233 ( \40576 , \40575 , \40190 );
and \U$40234 ( \40577 , \40574 , \40576 );
and \U$40235 ( \40578 , \40571 , \40573 );
or \U$40236 ( \40579 , \40577 , \40578 );
xor \U$40237 ( \40580 , \40193 , \40194 );
xor \U$40238 ( \40581 , \40580 , \40197 );
and \U$40239 ( \40582 , \40579 , \40581 );
not \U$40240 ( \40583 , \40582 );
or \U$40241 ( \40584 , \40205 , \40583 );
not \U$40242 ( \40585 , \40224 );
not \U$40243 ( \40586 , \40222 );
not \U$40244 ( \40587 , \40247 );
or \U$40245 ( \40588 , \40586 , \40587 );
or \U$40246 ( \40589 , \40247 , \40222 );
nand \U$40247 ( \40590 , \40588 , \40589 );
not \U$40248 ( \40591 , \40590 );
or \U$40249 ( \40592 , \40585 , \40591 );
or \U$40250 ( \40593 , \40590 , \40224 );
nand \U$40251 ( \40594 , \40592 , \40593 );
xor \U$40252 ( \40595 , \40295 , \40521 );
xor \U$40253 ( \40596 , \40595 , \40536 );
xor \U$40254 ( \40597 , \40594 , \40596 );
xor \U$40255 ( \40598 , \40127 , \40129 );
xor \U$40256 ( \40599 , \40598 , \40146 );
xor \U$40257 ( \40600 , \40207 , \40214 );
xor \U$40258 ( \40601 , \40599 , \40600 );
xor \U$40259 ( \40602 , \40597 , \40601 );
and \U$40260 ( \40603 , \7729 , RI986dd38_2);
and \U$40261 ( \40604 , RI986e1e8_12, \7727 );
nor \U$40262 ( \40605 , \40603 , \40604 );
and \U$40263 ( \40606 , \40605 , \7480 );
not \U$40264 ( \40607 , \40605 );
and \U$40265 ( \40608 , \40607 , \7733 );
nor \U$40266 ( \40609 , \40606 , \40608 );
nand \U$40267 ( \40610 , RI986e3c8_16, \9237 );
and \U$40268 ( \40611 , \40610 , \9241 );
not \U$40269 ( \40612 , \40610 );
and \U$40270 ( \40613 , \40612 , \8836 );
nor \U$40271 ( \40614 , \40611 , \40613 );
xor \U$40272 ( \40615 , \40609 , \40614 );
and \U$40273 ( \40616 , \8486 , RI986e0f8_10);
and \U$40274 ( \40617 , RI986e2d8_14, \8484 );
nor \U$40275 ( \40618 , \40616 , \40617 );
and \U$40276 ( \40619 , \40618 , \8050 );
not \U$40277 ( \40620 , \40618 );
and \U$40278 ( \40621 , \40620 , \8051 );
nor \U$40279 ( \40622 , \40619 , \40621 );
xor \U$40280 ( \40623 , \40615 , \40622 );
not \U$40281 ( \40624 , \4521 );
and \U$40282 ( \40625 , \4710 , RI986f778_58);
and \U$40283 ( \40626 , RI986fa48_64, \4708 );
nor \U$40284 ( \40627 , \40625 , \40626 );
not \U$40285 ( \40628 , \40627 );
or \U$40286 ( \40629 , \40624 , \40628 );
or \U$40287 ( \40630 , \40627 , \4521 );
nand \U$40288 ( \40631 , \40629 , \40630 );
and \U$40289 ( \40632 , \4203 , RI986e698_22);
and \U$40290 ( \40633 , RI986f868_60, \4201 );
nor \U$40291 ( \40634 , \40632 , \40633 );
and \U$40292 ( \40635 , \40634 , \4207 );
not \U$40293 ( \40636 , \40634 );
and \U$40294 ( \40637 , \40636 , \3922 );
nor \U$40295 ( \40638 , \40635 , \40637 );
xor \U$40296 ( \40639 , \40631 , \40638 );
and \U$40297 ( \40640 , \5318 , RI986f958_62);
and \U$40298 ( \40641 , RI986f4a8_52, \5316 );
nor \U$40299 ( \40642 , \40640 , \40641 );
and \U$40300 ( \40643 , \40642 , \5052 );
not \U$40301 ( \40644 , \40642 );
and \U$40302 ( \40645 , \40644 , \5322 );
nor \U$40303 ( \40646 , \40643 , \40645 );
xor \U$40304 ( \40647 , \40639 , \40646 );
and \U$40305 ( \40648 , \40623 , \40647 );
and \U$40306 ( \40649 , \5881 , RI986f3b8_50);
and \U$40307 ( \40650 , RI986f598_54, \5879 );
nor \U$40308 ( \40651 , \40649 , \40650 );
and \U$40309 ( \40652 , \40651 , \5594 );
not \U$40310 ( \40653 , \40651 );
and \U$40311 ( \40654 , \40653 , \5885 );
nor \U$40312 ( \40655 , \40652 , \40654 );
and \U$40313 ( \40656 , \6453 , RI986f688_56);
and \U$40314 ( \40657 , RI986e008_8, \6451 );
nor \U$40315 ( \40658 , \40656 , \40657 );
and \U$40316 ( \40659 , \40658 , \6190 );
not \U$40317 ( \40660 , \40658 );
and \U$40318 ( \40661 , \40660 , \6705 );
nor \U$40319 ( \40662 , \40659 , \40661 );
xor \U$40320 ( \40663 , \40655 , \40662 );
and \U$40321 ( \40664 , \7079 , RI986df18_6);
and \U$40322 ( \40665 , RI986de28_4, \7077 );
nor \U$40323 ( \40666 , \40664 , \40665 );
and \U$40324 ( \40667 , \40666 , \6710 );
not \U$40325 ( \40668 , \40666 );
and \U$40326 ( \40669 , \40668 , \6709 );
nor \U$40327 ( \40670 , \40667 , \40669 );
xor \U$40328 ( \40671 , \40663 , \40670 );
xor \U$40329 ( \40672 , \40631 , \40638 );
xor \U$40330 ( \40673 , \40672 , \40646 );
and \U$40331 ( \40674 , \40671 , \40673 );
and \U$40332 ( \40675 , \40623 , \40671 );
or \U$40333 ( \40676 , \40648 , \40674 , \40675 );
and \U$40334 ( \40677 , \416 , RI9870b28_100);
and \U$40335 ( \40678 , RI9870df8_106, \414 );
nor \U$40336 ( \40679 , \40677 , \40678 );
and \U$40337 ( \40680 , \40679 , \422 );
not \U$40338 ( \40681 , \40679 );
and \U$40339 ( \40682 , \40681 , \421 );
nor \U$40340 ( \40683 , \40680 , \40682 );
not \U$40341 ( \40684 , \487 );
and \U$40342 ( \40685 , \395 , RI9870c18_102);
and \U$40343 ( \40686 , RI98710c8_112, \393 );
nor \U$40344 ( \40687 , \40685 , \40686 );
not \U$40345 ( \40688 , \40687 );
or \U$40346 ( \40689 , \40684 , \40688 );
or \U$40347 ( \40690 , \40687 , \487 );
nand \U$40348 ( \40691 , \40689 , \40690 );
xor \U$40349 ( \40692 , \40683 , \40691 );
not \U$40350 ( \40693 , \345 );
and \U$40351 ( \40694 , \354 , RI9870a38_98);
and \U$40352 ( \40695 , RI9870ee8_108, \352 );
nor \U$40353 ( \40696 , \40694 , \40695 );
not \U$40354 ( \40697 , \40696 );
or \U$40355 ( \40698 , \40693 , \40697 );
or \U$40356 ( \40699 , \40696 , \361 );
nand \U$40357 ( \40700 , \40698 , \40699 );
xor \U$40358 ( \40701 , \40692 , \40700 );
nand \U$40359 ( \40702 , RI9870fd8_110, RI9871fc8_144);
xor \U$40360 ( \40703 , \40701 , \40702 );
and \U$40361 ( \40704 , \438 , RI9871488_120);
and \U$40362 ( \40705 , RI9871758_126, \436 );
nor \U$40363 ( \40706 , \40704 , \40705 );
and \U$40364 ( \40707 , \40706 , \444 );
not \U$40365 ( \40708 , \40706 );
and \U$40366 ( \40709 , \40708 , \443 );
nor \U$40367 ( \40710 , \40707 , \40709 );
not \U$40368 ( \40711 , \454 );
and \U$40369 ( \40712 , \465 , RI98711b8_114);
and \U$40370 ( \40713 , RI9871398_118, \463 );
nor \U$40371 ( \40714 , \40712 , \40713 );
not \U$40372 ( \40715 , \40714 );
or \U$40373 ( \40716 , \40711 , \40715 );
or \U$40374 ( \40717 , \40714 , \456 );
nand \U$40375 ( \40718 , \40716 , \40717 );
xor \U$40376 ( \40719 , \40710 , \40718 );
not \U$40377 ( \40720 , \367 );
and \U$40378 ( \40721 , \376 , RI9870d08_104);
and \U$40379 ( \40722 , RI98712a8_116, \374 );
nor \U$40380 ( \40723 , \40721 , \40722 );
not \U$40381 ( \40724 , \40723 );
or \U$40382 ( \40725 , \40720 , \40724 );
or \U$40383 ( \40726 , \40723 , \367 );
nand \U$40384 ( \40727 , \40725 , \40726 );
xor \U$40385 ( \40728 , \40719 , \40727 );
and \U$40386 ( \40729 , \40703 , \40728 );
and \U$40387 ( \40730 , \40701 , \40702 );
or \U$40388 ( \40731 , \40729 , \40730 );
xor \U$40389 ( \40732 , \40676 , \40731 );
not \U$40390 ( \40733 , \1128 );
and \U$40391 ( \40734 , \1293 , RI9871668_124);
and \U$40392 ( \40735 , RI986eb48_32, \1291 );
nor \U$40393 ( \40736 , \40734 , \40735 );
not \U$40394 ( \40737 , \40736 );
or \U$40395 ( \40738 , \40733 , \40737 );
or \U$40396 ( \40739 , \40736 , \1128 );
nand \U$40397 ( \40740 , \40738 , \40739 );
and \U$40398 ( \40741 , \776 , RI9871848_128);
and \U$40399 ( \40742 , RI9871578_122, \774 );
nor \U$40400 ( \40743 , \40741 , \40742 );
and \U$40401 ( \40744 , \40743 , \474 );
not \U$40402 ( \40745 , \40743 );
and \U$40403 ( \40746 , \40745 , \451 );
nor \U$40404 ( \40747 , \40744 , \40746 );
xor \U$40405 ( \40748 , \40740 , \40747 );
and \U$40406 ( \40749 , \1329 , RI986ea58_30);
and \U$40407 ( \40750 , RI986e968_28, \1327 );
nor \U$40408 ( \40751 , \40749 , \40750 );
and \U$40409 ( \40752 , \40751 , \1336 );
not \U$40410 ( \40753 , \40751 );
and \U$40411 ( \40754 , \40753 , \1337 );
nor \U$40412 ( \40755 , \40752 , \40754 );
xor \U$40413 ( \40756 , \40748 , \40755 );
and \U$40414 ( \40757 , \1311 , RI986e878_26);
and \U$40415 ( \40758 , RI986ef08_40, \1309 );
nor \U$40416 ( \40759 , \40757 , \40758 );
and \U$40417 ( \40760 , \40759 , \1458 );
not \U$40418 ( \40761 , \40759 );
and \U$40419 ( \40762 , \40761 , \1318 );
nor \U$40420 ( \40763 , \40760 , \40762 );
not \U$40421 ( \40764 , \1462 );
and \U$40422 ( \40765 , \2042 , RI986ee18_38);
and \U$40423 ( \40766 , RI986ec38_34, \2040 );
nor \U$40424 ( \40767 , \40765 , \40766 );
not \U$40425 ( \40768 , \40767 );
or \U$40426 ( \40769 , \40764 , \40768 );
or \U$40427 ( \40770 , \40767 , \2034 );
nand \U$40428 ( \40771 , \40769 , \40770 );
xor \U$40429 ( \40772 , \40763 , \40771 );
and \U$40430 ( \40773 , \2274 , RI986ed28_36);
and \U$40431 ( \40774 , RI986f0e8_44, \2272 );
nor \U$40432 ( \40775 , \40773 , \40774 );
and \U$40433 ( \40776 , \40775 , \2030 );
not \U$40434 ( \40777 , \40775 );
and \U$40435 ( \40778 , \40777 , \2031 );
nor \U$40436 ( \40779 , \40776 , \40778 );
xor \U$40437 ( \40780 , \40772 , \40779 );
and \U$40438 ( \40781 , \40756 , \40780 );
and \U$40439 ( \40782 , \2464 , RI986eff8_42);
and \U$40440 ( \40783 , RI986f2c8_48, \2462 );
nor \U$40441 ( \40784 , \40782 , \40783 );
and \U$40442 ( \40785 , \40784 , \2468 );
not \U$40443 ( \40786 , \40784 );
and \U$40444 ( \40787 , \40786 , \2263 );
nor \U$40445 ( \40788 , \40785 , \40787 );
not \U$40446 ( \40789 , \3406 );
and \U$40447 ( \40790 , \3254 , RI986f1d8_46);
and \U$40448 ( \40791 , RI986e5a8_20, \3252 );
nor \U$40449 ( \40792 , \40790 , \40791 );
not \U$40450 ( \40793 , \40792 );
or \U$40451 ( \40794 , \40789 , \40793 );
or \U$40452 ( \40795 , \40792 , \3406 );
nand \U$40453 ( \40796 , \40794 , \40795 );
xor \U$40454 ( \40797 , \40788 , \40796 );
not \U$40455 ( \40798 , \3918 );
and \U$40456 ( \40799 , \3683 , RI986e4b8_18);
and \U$40457 ( \40800 , RI986e788_24, \3681 );
nor \U$40458 ( \40801 , \40799 , \40800 );
not \U$40459 ( \40802 , \40801 );
or \U$40460 ( \40803 , \40798 , \40802 );
or \U$40461 ( \40804 , \40801 , \3918 );
nand \U$40462 ( \40805 , \40803 , \40804 );
xor \U$40463 ( \40806 , \40797 , \40805 );
xor \U$40464 ( \40807 , \40763 , \40771 );
xor \U$40465 ( \40808 , \40807 , \40779 );
and \U$40466 ( \40809 , \40806 , \40808 );
and \U$40467 ( \40810 , \40756 , \40806 );
or \U$40468 ( \40811 , \40781 , \40809 , \40810 );
and \U$40469 ( \40812 , \40732 , \40811 );
and \U$40470 ( \40813 , \40676 , \40731 );
or \U$40471 ( \40814 , \40812 , \40813 );
and \U$40472 ( \40815 , \5318 , RI986fa48_64);
and \U$40473 ( \40816 , RI986f958_62, \5316 );
nor \U$40474 ( \40817 , \40815 , \40816 );
and \U$40475 ( \40818 , \40817 , \5052 );
not \U$40476 ( \40819 , \40817 );
and \U$40477 ( \40820 , \40819 , \5322 );
nor \U$40478 ( \40821 , \40818 , \40820 );
not \U$40479 ( \40822 , \4521 );
and \U$40480 ( \40823 , \4710 , RI986f868_60);
and \U$40481 ( \40824 , RI986f778_58, \4708 );
nor \U$40482 ( \40825 , \40823 , \40824 );
not \U$40483 ( \40826 , \40825 );
or \U$40484 ( \40827 , \40822 , \40826 );
or \U$40485 ( \40828 , \40825 , \4519 );
nand \U$40486 ( \40829 , \40827 , \40828 );
xor \U$40487 ( \40830 , \40821 , \40829 );
and \U$40488 ( \40831 , \5881 , RI986f4a8_52);
and \U$40489 ( \40832 , RI986f3b8_50, \5879 );
nor \U$40490 ( \40833 , \40831 , \40832 );
and \U$40491 ( \40834 , \40833 , \5594 );
not \U$40492 ( \40835 , \40833 );
and \U$40493 ( \40836 , \40835 , \5885 );
nor \U$40494 ( \40837 , \40834 , \40836 );
and \U$40495 ( \40838 , \40830 , \40837 );
and \U$40496 ( \40839 , \40821 , \40829 );
or \U$40497 ( \40840 , \40838 , \40839 );
and \U$40498 ( \40841 , \9237 , RI986e2d8_14);
and \U$40499 ( \40842 , RI986e3c8_16, \9235 );
nor \U$40500 ( \40843 , \40841 , \40842 );
and \U$40501 ( \40844 , \40843 , \9241 );
not \U$40502 ( \40845 , \40843 );
and \U$40503 ( \40846 , \40845 , \8836 );
nor \U$40504 ( \40847 , \40844 , \40846 );
xor \U$40505 ( \40848 , \40847 , \9510 );
and \U$40506 ( \40849 , \8486 , RI986e1e8_12);
and \U$40507 ( \40850 , RI986e0f8_10, \8484 );
nor \U$40508 ( \40851 , \40849 , \40850 );
and \U$40509 ( \40852 , \40851 , \8050 );
not \U$40510 ( \40853 , \40851 );
and \U$40511 ( \40854 , \40853 , \8051 );
nor \U$40512 ( \40855 , \40852 , \40854 );
and \U$40513 ( \40856 , \40848 , \40855 );
and \U$40514 ( \40857 , \40847 , \9510 );
or \U$40515 ( \40858 , \40856 , \40857 );
xor \U$40516 ( \40859 , \40840 , \40858 );
and \U$40517 ( \40860 , \6453 , RI986f598_54);
and \U$40518 ( \40861 , RI986f688_56, \6451 );
nor \U$40519 ( \40862 , \40860 , \40861 );
and \U$40520 ( \40863 , \40862 , \6190 );
not \U$40521 ( \40864 , \40862 );
and \U$40522 ( \40865 , \40864 , \6180 );
nor \U$40523 ( \40866 , \40863 , \40865 );
and \U$40524 ( \40867 , \7079 , RI986e008_8);
and \U$40525 ( \40868 , RI986df18_6, \7077 );
nor \U$40526 ( \40869 , \40867 , \40868 );
and \U$40527 ( \40870 , \40869 , \6710 );
not \U$40528 ( \40871 , \40869 );
and \U$40529 ( \40872 , \40871 , \6709 );
nor \U$40530 ( \40873 , \40870 , \40872 );
xor \U$40531 ( \40874 , \40866 , \40873 );
and \U$40532 ( \40875 , \7729 , RI986de28_4);
and \U$40533 ( \40876 , RI986dd38_2, \7727 );
nor \U$40534 ( \40877 , \40875 , \40876 );
and \U$40535 ( \40878 , \40877 , \7480 );
not \U$40536 ( \40879 , \40877 );
and \U$40537 ( \40880 , \40879 , \7733 );
nor \U$40538 ( \40881 , \40878 , \40880 );
and \U$40539 ( \40882 , \40874 , \40881 );
and \U$40540 ( \40883 , \40866 , \40873 );
or \U$40541 ( \40884 , \40882 , \40883 );
and \U$40542 ( \40885 , \40859 , \40884 );
and \U$40543 ( \40886 , \40840 , \40858 );
or \U$40544 ( \40887 , \40885 , \40886 );
not \U$40545 ( \40888 , \367 );
and \U$40546 ( \40889 , \376 , RI98710c8_112);
and \U$40547 ( \40890 , RI9870d08_104, \374 );
nor \U$40548 ( \40891 , \40889 , \40890 );
not \U$40549 ( \40892 , \40891 );
or \U$40550 ( \40893 , \40888 , \40892 );
or \U$40551 ( \40894 , \40891 , \365 );
nand \U$40552 ( \40895 , \40893 , \40894 );
not \U$40553 ( \40896 , \487 );
and \U$40554 ( \40897 , \395 , RI9870ee8_108);
and \U$40555 ( \40898 , RI9870c18_102, \393 );
nor \U$40556 ( \40899 , \40897 , \40898 );
not \U$40557 ( \40900 , \40899 );
or \U$40558 ( \40901 , \40896 , \40900 );
or \U$40559 ( \40902 , \40899 , \386 );
nand \U$40560 ( \40903 , \40901 , \40902 );
xor \U$40561 ( \40904 , \40895 , \40903 );
not \U$40562 ( \40905 , \345 );
and \U$40563 ( \40906 , \354 , RI9870df8_106);
and \U$40564 ( \40907 , RI9870a38_98, \352 );
nor \U$40565 ( \40908 , \40906 , \40907 );
not \U$40566 ( \40909 , \40908 );
or \U$40567 ( \40910 , \40905 , \40909 );
or \U$40568 ( \40911 , \40908 , \361 );
nand \U$40569 ( \40912 , \40910 , \40911 );
and \U$40570 ( \40913 , \40904 , \40912 );
and \U$40571 ( \40914 , \40895 , \40903 );
or \U$40572 ( \40915 , \40913 , \40914 );
not \U$40573 ( \40916 , RI98701c8_80);
nor \U$40574 ( \40917 , \40916 , \407 );
and \U$40575 ( \40918 , \416 , RI9870fd8_110);
and \U$40576 ( \40919 , RI9870b28_100, \414 );
nor \U$40577 ( \40920 , \40918 , \40919 );
and \U$40578 ( \40921 , \40920 , \422 );
not \U$40579 ( \40922 , \40920 );
and \U$40580 ( \40923 , \40922 , \421 );
nor \U$40581 ( \40924 , \40921 , \40923 );
and \U$40582 ( \40925 , \40917 , \40924 );
xor \U$40583 ( \40926 , \40915 , \40925 );
and \U$40584 ( \40927 , \776 , RI9871758_126);
and \U$40585 ( \40928 , RI9871848_128, \774 );
nor \U$40586 ( \40929 , \40927 , \40928 );
and \U$40587 ( \40930 , \40929 , \474 );
not \U$40588 ( \40931 , \40929 );
and \U$40589 ( \40932 , \40931 , \451 );
nor \U$40590 ( \40933 , \40930 , \40932 );
and \U$40591 ( \40934 , \438 , RI9871398_118);
and \U$40592 ( \40935 , RI9871488_120, \436 );
nor \U$40593 ( \40936 , \40934 , \40935 );
and \U$40594 ( \40937 , \40936 , \444 );
not \U$40595 ( \40938 , \40936 );
and \U$40596 ( \40939 , \40938 , \443 );
nor \U$40597 ( \40940 , \40937 , \40939 );
xor \U$40598 ( \40941 , \40933 , \40940 );
not \U$40599 ( \40942 , \454 );
and \U$40600 ( \40943 , \465 , RI98712a8_116);
and \U$40601 ( \40944 , RI98711b8_114, \463 );
nor \U$40602 ( \40945 , \40943 , \40944 );
not \U$40603 ( \40946 , \40945 );
or \U$40604 ( \40947 , \40942 , \40946 );
or \U$40605 ( \40948 , \40945 , \456 );
nand \U$40606 ( \40949 , \40947 , \40948 );
and \U$40607 ( \40950 , \40941 , \40949 );
and \U$40608 ( \40951 , \40933 , \40940 );
or \U$40609 ( \40952 , \40950 , \40951 );
and \U$40610 ( \40953 , \40926 , \40952 );
and \U$40611 ( \40954 , \40915 , \40925 );
or \U$40612 ( \40955 , \40953 , \40954 );
xor \U$40613 ( \40956 , \40887 , \40955 );
and \U$40614 ( \40957 , \2464 , RI986f0e8_44);
and \U$40615 ( \40958 , RI986eff8_42, \2462 );
nor \U$40616 ( \40959 , \40957 , \40958 );
and \U$40617 ( \40960 , \40959 , \2468 );
not \U$40618 ( \40961 , \40959 );
and \U$40619 ( \40962 , \40961 , \2263 );
nor \U$40620 ( \40963 , \40960 , \40962 );
not \U$40621 ( \40964 , \1462 );
and \U$40622 ( \40965 , \2042 , RI986ef08_40);
and \U$40623 ( \40966 , RI986ee18_38, \2040 );
nor \U$40624 ( \40967 , \40965 , \40966 );
not \U$40625 ( \40968 , \40967 );
or \U$40626 ( \40969 , \40964 , \40968 );
or \U$40627 ( \40970 , \40967 , \1462 );
nand \U$40628 ( \40971 , \40969 , \40970 );
xor \U$40629 ( \40972 , \40963 , \40971 );
and \U$40630 ( \40973 , \2274 , RI986ec38_34);
and \U$40631 ( \40974 , RI986ed28_36, \2272 );
nor \U$40632 ( \40975 , \40973 , \40974 );
and \U$40633 ( \40976 , \40975 , \2030 );
not \U$40634 ( \40977 , \40975 );
and \U$40635 ( \40978 , \40977 , \2031 );
nor \U$40636 ( \40979 , \40976 , \40978 );
and \U$40637 ( \40980 , \40972 , \40979 );
and \U$40638 ( \40981 , \40963 , \40971 );
or \U$40639 ( \40982 , \40980 , \40981 );
and \U$40640 ( \40983 , \1311 , RI986e968_28);
and \U$40641 ( \40984 , RI986e878_26, \1309 );
nor \U$40642 ( \40985 , \40983 , \40984 );
and \U$40643 ( \40986 , \40985 , \1458 );
not \U$40644 ( \40987 , \40985 );
and \U$40645 ( \40988 , \40987 , \1318 );
nor \U$40646 ( \40989 , \40986 , \40988 );
not \U$40647 ( \40990 , \1128 );
and \U$40648 ( \40991 , \1293 , RI9871578_122);
and \U$40649 ( \40992 , RI9871668_124, \1291 );
nor \U$40650 ( \40993 , \40991 , \40992 );
not \U$40651 ( \40994 , \40993 );
or \U$40652 ( \40995 , \40990 , \40994 );
or \U$40653 ( \40996 , \40993 , \1128 );
nand \U$40654 ( \40997 , \40995 , \40996 );
xor \U$40655 ( \40998 , \40989 , \40997 );
and \U$40656 ( \40999 , \1329 , RI986eb48_32);
and \U$40657 ( \41000 , RI986ea58_30, \1327 );
nor \U$40658 ( \41001 , \40999 , \41000 );
and \U$40659 ( \41002 , \41001 , \1336 );
not \U$40660 ( \41003 , \41001 );
and \U$40661 ( \41004 , \41003 , \1337 );
nor \U$40662 ( \41005 , \41002 , \41004 );
and \U$40663 ( \41006 , \40998 , \41005 );
and \U$40664 ( \41007 , \40989 , \40997 );
or \U$40665 ( \41008 , \41006 , \41007 );
xor \U$40666 ( \41009 , \40982 , \41008 );
and \U$40667 ( \41010 , \4203 , RI986e788_24);
and \U$40668 ( \41011 , RI986e698_22, \4201 );
nor \U$40669 ( \41012 , \41010 , \41011 );
and \U$40670 ( \41013 , \41012 , \4207 );
not \U$40671 ( \41014 , \41012 );
and \U$40672 ( \41015 , \41014 , \3923 );
nor \U$40673 ( \41016 , \41013 , \41015 );
not \U$40674 ( \41017 , \3406 );
and \U$40675 ( \41018 , \3254 , RI986f2c8_48);
and \U$40676 ( \41019 , RI986f1d8_46, \3252 );
nor \U$40677 ( \41020 , \41018 , \41019 );
not \U$40678 ( \41021 , \41020 );
or \U$40679 ( \41022 , \41017 , \41021 );
or \U$40680 ( \41023 , \41020 , \3406 );
nand \U$40681 ( \41024 , \41022 , \41023 );
xor \U$40682 ( \41025 , \41016 , \41024 );
not \U$40683 ( \41026 , \3918 );
and \U$40684 ( \41027 , \3683 , RI986e5a8_20);
and \U$40685 ( \41028 , RI986e4b8_18, \3681 );
nor \U$40686 ( \41029 , \41027 , \41028 );
not \U$40687 ( \41030 , \41029 );
or \U$40688 ( \41031 , \41026 , \41030 );
or \U$40689 ( \41032 , \41029 , \3412 );
nand \U$40690 ( \41033 , \41031 , \41032 );
and \U$40691 ( \41034 , \41025 , \41033 );
and \U$40692 ( \41035 , \41016 , \41024 );
or \U$40693 ( \41036 , \41034 , \41035 );
and \U$40694 ( \41037 , \41009 , \41036 );
and \U$40695 ( \41038 , \40982 , \41008 );
or \U$40696 ( \41039 , \41037 , \41038 );
and \U$40697 ( \41040 , \40956 , \41039 );
and \U$40698 ( \41041 , \40887 , \40955 );
or \U$40699 ( \41042 , \41040 , \41041 );
xor \U$40700 ( \41043 , \40814 , \41042 );
xor \U$40701 ( \41044 , \40330 , \40338 );
xor \U$40702 ( \41045 , \41044 , \40346 );
not \U$40703 ( \41046 , \41045 );
nand \U$40704 ( \41047 , RI9870b28_100, RI9871fc8_144);
xor \U$40705 ( \41048 , \40303 , \40310 );
xor \U$40706 ( \41049 , \41048 , \40319 );
xor \U$40707 ( \41050 , \41047 , \41049 );
not \U$40708 ( \41051 , \41050 );
or \U$40709 ( \41052 , \41046 , \41051 );
or \U$40710 ( \41053 , \41050 , \41045 );
nand \U$40711 ( \41054 , \41052 , \41053 );
not \U$40712 ( \41055 , \40449 );
and \U$40713 ( \41056 , \40460 , \8836 );
not \U$40714 ( \41057 , \40460 );
and \U$40715 ( \41058 , \41057 , \9241 );
nor \U$40716 ( \41059 , \41056 , \41058 );
not \U$40717 ( \41060 , \41059 );
or \U$40718 ( \41061 , \41055 , \41060 );
or \U$40719 ( \41062 , \41059 , \40449 );
nand \U$40720 ( \41063 , \41061 , \41062 );
xor \U$40721 ( \41064 , \40498 , \40505 );
xor \U$40722 ( \41065 , \41064 , \40513 );
xor \U$40723 ( \41066 , \41063 , \41065 );
not \U$40724 ( \41067 , \40469 );
xor \U$40725 ( \41068 , \40477 , \40487 );
not \U$40726 ( \41069 , \41068 );
or \U$40727 ( \41070 , \41067 , \41069 );
or \U$40728 ( \41071 , \41068 , \40469 );
nand \U$40729 ( \41072 , \41070 , \41071 );
xor \U$40730 ( \41073 , \41066 , \41072 );
and \U$40731 ( \41074 , \41054 , \41073 );
xor \U$40732 ( \41075 , \40360 , \40367 );
xor \U$40733 ( \41076 , \41075 , \40375 );
not \U$40734 ( \41077 , \40385 );
xor \U$40735 ( \41078 , \40394 , \40404 );
not \U$40736 ( \41079 , \41078 );
or \U$40737 ( \41080 , \41077 , \41079 );
or \U$40738 ( \41081 , \41078 , \40385 );
nand \U$40739 ( \41082 , \41080 , \41081 );
xor \U$40740 ( \41083 , \41076 , \41082 );
not \U$40741 ( \41084 , \40414 );
xor \U$40742 ( \41085 , \40423 , \40434 );
not \U$40743 ( \41086 , \41085 );
or \U$40744 ( \41087 , \41084 , \41086 );
or \U$40745 ( \41088 , \41085 , \40414 );
nand \U$40746 ( \41089 , \41087 , \41088 );
xor \U$40747 ( \41090 , \41083 , \41089 );
xor \U$40748 ( \41091 , \41063 , \41065 );
xor \U$40749 ( \41092 , \41091 , \41072 );
and \U$40750 ( \41093 , \41090 , \41092 );
and \U$40751 ( \41094 , \41054 , \41090 );
or \U$40752 ( \41095 , \41074 , \41093 , \41094 );
and \U$40753 ( \41096 , \41043 , \41095 );
and \U$40754 ( \41097 , \40814 , \41042 );
or \U$40755 ( \41098 , \41096 , \41097 );
xor \U$40756 ( \41099 , \40788 , \40796 );
and \U$40757 ( \41100 , \41099 , \40805 );
and \U$40758 ( \41101 , \40788 , \40796 );
or \U$40759 ( \41102 , \41100 , \41101 );
xor \U$40760 ( \41103 , \40763 , \40771 );
and \U$40761 ( \41104 , \41103 , \40779 );
and \U$40762 ( \41105 , \40763 , \40771 );
or \U$40763 ( \41106 , \41104 , \41105 );
xor \U$40764 ( \41107 , \41102 , \41106 );
xor \U$40765 ( \41108 , \40740 , \40747 );
and \U$40766 ( \41109 , \41108 , \40755 );
and \U$40767 ( \41110 , \40740 , \40747 );
or \U$40768 ( \41111 , \41109 , \41110 );
and \U$40769 ( \41112 , \41107 , \41111 );
and \U$40770 ( \41113 , \41102 , \41106 );
or \U$40771 ( \41114 , \41112 , \41113 );
xor \U$40772 ( \41115 , \40683 , \40691 );
and \U$40773 ( \41116 , \41115 , \40700 );
and \U$40774 ( \41117 , \40683 , \40691 );
or \U$40775 ( \41118 , \41116 , \41117 );
not \U$40776 ( \41119 , \40702 );
xor \U$40777 ( \41120 , \41118 , \41119 );
xor \U$40778 ( \41121 , \40710 , \40718 );
and \U$40779 ( \41122 , \41121 , \40727 );
and \U$40780 ( \41123 , \40710 , \40718 );
or \U$40781 ( \41124 , \41122 , \41123 );
and \U$40782 ( \41125 , \41120 , \41124 );
and \U$40783 ( \41126 , \41118 , \41119 );
or \U$40784 ( \41127 , \41125 , \41126 );
xor \U$40785 ( \41128 , \41114 , \41127 );
xor \U$40786 ( \41129 , \40655 , \40662 );
and \U$40787 ( \41130 , \41129 , \40670 );
and \U$40788 ( \41131 , \40655 , \40662 );
or \U$40789 ( \41132 , \41130 , \41131 );
xor \U$40790 ( \41133 , \40609 , \40614 );
and \U$40791 ( \41134 , \41133 , \40622 );
and \U$40792 ( \41135 , \40609 , \40614 );
or \U$40793 ( \41136 , \41134 , \41135 );
xor \U$40794 ( \41137 , \41132 , \41136 );
xor \U$40795 ( \41138 , \40631 , \40638 );
and \U$40796 ( \41139 , \41138 , \40646 );
and \U$40797 ( \41140 , \40631 , \40638 );
or \U$40798 ( \41141 , \41139 , \41140 );
and \U$40799 ( \41142 , \41137 , \41141 );
and \U$40800 ( \41143 , \41132 , \41136 );
or \U$40801 ( \41144 , \41142 , \41143 );
xor \U$40802 ( \41145 , \41128 , \41144 );
not \U$40803 ( \41146 , \41045 );
not \U$40804 ( \41147 , \41047 );
and \U$40805 ( \41148 , \41146 , \41147 );
and \U$40806 ( \41149 , \41045 , \41047 );
nor \U$40807 ( \41150 , \41149 , \41049 );
nor \U$40808 ( \41151 , \41148 , \41150 );
not \U$40809 ( \41152 , \41151 );
xor \U$40810 ( \41153 , \41076 , \41082 );
and \U$40811 ( \41154 , \41153 , \41089 );
and \U$40812 ( \41155 , \41076 , \41082 );
or \U$40813 ( \41156 , \41154 , \41155 );
xor \U$40814 ( \41157 , \41063 , \41065 );
and \U$40815 ( \41158 , \41157 , \41072 );
and \U$40816 ( \41159 , \41063 , \41065 );
or \U$40817 ( \41160 , \41158 , \41159 );
xor \U$40818 ( \41161 , \41156 , \41160 );
not \U$40819 ( \41162 , \41161 );
or \U$40820 ( \41163 , \41152 , \41162 );
or \U$40821 ( \41164 , \41161 , \41151 );
nand \U$40822 ( \41165 , \41163 , \41164 );
and \U$40823 ( \41166 , \41145 , \41165 );
xor \U$40824 ( \41167 , \41098 , \41166 );
and \U$40825 ( \41168 , \40322 , \40349 );
nor \U$40826 ( \41169 , \41168 , \40350 );
not \U$40827 ( \41170 , \41169 );
xor \U$40828 ( \41171 , \40462 , \40489 );
xor \U$40829 ( \41172 , \41171 , \40516 );
xor \U$40830 ( \41173 , \40378 , \40406 );
xor \U$40831 ( \41174 , \41173 , \40436 );
xor \U$40832 ( \41175 , \41172 , \41174 );
not \U$40833 ( \41176 , \41175 );
or \U$40834 ( \41177 , \41170 , \41176 );
or \U$40835 ( \41178 , \41175 , \41169 );
nand \U$40836 ( \41179 , \41177 , \41178 );
xor \U$40837 ( \41180 , \41118 , \41119 );
xor \U$40838 ( \41181 , \41180 , \41124 );
xor \U$40839 ( \41182 , \41132 , \41136 );
xor \U$40840 ( \41183 , \41182 , \41141 );
xor \U$40841 ( \41184 , \41181 , \41183 );
xor \U$40842 ( \41185 , \41102 , \41106 );
xor \U$40843 ( \41186 , \41185 , \41111 );
and \U$40844 ( \41187 , \41184 , \41186 );
and \U$40845 ( \41188 , \41181 , \41183 );
or \U$40846 ( \41189 , \41187 , \41188 );
xor \U$40847 ( \41190 , \41179 , \41189 );
not \U$40848 ( \41191 , \40280 );
not \U$40849 ( \41192 , \40277 );
and \U$40850 ( \41193 , \41191 , \41192 );
and \U$40851 ( \41194 , \40280 , \40277 );
nor \U$40852 ( \41195 , \41193 , \41194 );
not \U$40853 ( \41196 , \41195 );
xor \U$40854 ( \41197 , \40284 , \40286 );
xor \U$40855 ( \41198 , \41197 , \40289 );
xor \U$40856 ( \41199 , \40255 , \40257 );
xor \U$40857 ( \41200 , \41199 , \40268 );
xor \U$40858 ( \41201 , \41198 , \41200 );
not \U$40859 ( \41202 , \41201 );
or \U$40860 ( \41203 , \41196 , \41202 );
or \U$40861 ( \41204 , \41201 , \41195 );
nand \U$40862 ( \41205 , \41203 , \41204 );
and \U$40863 ( \41206 , \41190 , \41205 );
and \U$40864 ( \41207 , \41179 , \41189 );
or \U$40865 ( \41208 , \41206 , \41207 );
and \U$40866 ( \41209 , \41167 , \41208 );
and \U$40867 ( \41210 , \41098 , \41166 );
or \U$40868 ( \41211 , \41209 , \41210 );
and \U$40869 ( \41212 , \40602 , \41211 );
not \U$40870 ( \41213 , \40602 );
not \U$40871 ( \41214 , \41211 );
and \U$40872 ( \41215 , \41213 , \41214 );
xor \U$40873 ( \41216 , \40271 , \40281 );
xor \U$40874 ( \41217 , \41216 , \40292 );
not \U$40875 ( \41218 , \41217 );
xnor \U$40876 ( \41219 , \40439 , \40519 );
not \U$40877 ( \41220 , \41219 );
not \U$40878 ( \41221 , \40351 );
and \U$40879 ( \41222 , \41220 , \41221 );
and \U$40880 ( \41223 , \41219 , \40351 );
nor \U$40881 ( \41224 , \41222 , \41223 );
not \U$40882 ( \41225 , \41224 );
and \U$40883 ( \41226 , \41218 , \41225 );
and \U$40884 ( \41227 , \41217 , \41224 );
nor \U$40885 ( \41228 , \41226 , \41227 );
and \U$40886 ( \41229 , \41160 , \41156 );
not \U$40887 ( \41230 , \41156 );
not \U$40888 ( \41231 , \41160 );
and \U$40889 ( \41232 , \41230 , \41231 );
nor \U$40890 ( \41233 , \41232 , \41151 );
nor \U$40891 ( \41234 , \41229 , \41233 );
xor \U$40892 ( \41235 , \41114 , \41127 );
and \U$40893 ( \41236 , \41235 , \41144 );
and \U$40894 ( \41237 , \41114 , \41127 );
nor \U$40895 ( \41238 , \41236 , \41237 );
xor \U$40896 ( \41239 , \41234 , \41238 );
not \U$40897 ( \41240 , \41200 );
not \U$40898 ( \41241 , \41195 );
and \U$40899 ( \41242 , \41240 , \41241 );
and \U$40900 ( \41243 , \41200 , \41195 );
nor \U$40901 ( \41244 , \41243 , \41198 );
nor \U$40902 ( \41245 , \41242 , \41244 );
xor \U$40903 ( \41246 , \41239 , \41245 );
and \U$40904 ( \41247 , \41228 , \41246 );
not \U$40905 ( \41248 , \41174 );
not \U$40906 ( \41249 , \41169 );
and \U$40907 ( \41250 , \41248 , \41249 );
and \U$40908 ( \41251 , \41174 , \41169 );
nor \U$40909 ( \41252 , \41251 , \41172 );
nor \U$40910 ( \41253 , \41250 , \41252 );
not \U$40911 ( \41254 , \41253 );
xor \U$40912 ( \41255 , \40115 , \40117 );
xor \U$40913 ( \41256 , \41255 , \40124 );
xor \U$40914 ( \41257 , \40524 , \40531 );
xor \U$40915 ( \41258 , \41256 , \41257 );
not \U$40916 ( \41259 , \41258 );
or \U$40917 ( \41260 , \41254 , \41259 );
or \U$40918 ( \41261 , \41258 , \41253 );
nand \U$40919 ( \41262 , \41260 , \41261 );
not \U$40920 ( \41263 , \41262 );
xor \U$40921 ( \41264 , \40239 , \40241 );
xor \U$40922 ( \41265 , \41264 , \40244 );
not \U$40923 ( \41266 , \41265 );
and \U$40924 ( \41267 , \41263 , \41266 );
and \U$40925 ( \41268 , \41262 , \41265 );
nor \U$40926 ( \41269 , \41267 , \41268 );
xor \U$40927 ( \41270 , \41234 , \41238 );
xor \U$40928 ( \41271 , \41270 , \41245 );
and \U$40929 ( \41272 , \41269 , \41271 );
and \U$40930 ( \41273 , \41228 , \41269 );
or \U$40931 ( \41274 , \41247 , \41272 , \41273 );
nor \U$40932 ( \41275 , \41215 , \41274 );
nor \U$40933 ( \41276 , \41212 , \41275 );
not \U$40934 ( \41277 , \40249 );
not \U$40935 ( \41278 , \40539 );
or \U$40936 ( \41279 , \41277 , \41278 );
or \U$40937 ( \41280 , \40539 , \40249 );
nand \U$40938 ( \41281 , \41279 , \41280 );
not \U$40939 ( \41282 , \41281 );
not \U$40940 ( \41283 , \40220 );
and \U$40941 ( \41284 , \41282 , \41283 );
and \U$40942 ( \41285 , \41281 , \40220 );
nor \U$40943 ( \41286 , \41284 , \41285 );
xor \U$40944 ( \41287 , \41276 , \41286 );
xor \U$40945 ( \41288 , \40594 , \40596 );
and \U$40946 ( \41289 , \41288 , \40601 );
and \U$40947 ( \41290 , \40594 , \40596 );
nor \U$40948 ( \41291 , \41289 , \41290 );
or \U$40949 ( \41292 , \41265 , \41253 );
not \U$40950 ( \41293 , \41253 );
not \U$40951 ( \41294 , \41265 );
or \U$40952 ( \41295 , \41293 , \41294 );
nand \U$40953 ( \41296 , \41295 , \41258 );
nand \U$40954 ( \41297 , \41292 , \41296 );
not \U$40955 ( \41298 , \41224 );
nand \U$40956 ( \41299 , \41298 , \41217 );
not \U$40957 ( \41300 , \41299 );
and \U$40958 ( \41301 , \41297 , \41300 );
not \U$40959 ( \41302 , \41297 );
not \U$40960 ( \41303 , \41300 );
and \U$40961 ( \41304 , \41302 , \41303 );
xor \U$40962 ( \41305 , \41234 , \41238 );
and \U$40963 ( \41306 , \41305 , \41245 );
and \U$40964 ( \41307 , \41234 , \41238 );
or \U$40965 ( \41308 , \41306 , \41307 );
nor \U$40966 ( \41309 , \41304 , \41308 );
nor \U$40967 ( \41310 , \41301 , \41309 );
xor \U$40968 ( \41311 , \41291 , \41310 );
xnor \U$40969 ( \41312 , \40553 , \40547 );
not \U$40970 ( \41313 , \41312 );
not \U$40971 ( \41314 , \40561 );
and \U$40972 ( \41315 , \41313 , \41314 );
and \U$40973 ( \41316 , \41312 , \40561 );
nor \U$40974 ( \41317 , \41315 , \41316 );
xor \U$40975 ( \41318 , \41311 , \41317 );
and \U$40976 ( \41319 , \41287 , \41318 );
and \U$40977 ( \41320 , \41276 , \41286 );
or \U$40978 ( \41321 , \41319 , \41320 );
not \U$40979 ( \41322 , \41321 );
xor \U$40980 ( \41323 , \40541 , \40563 );
xor \U$40981 ( \41324 , \41323 , \40568 );
not \U$40982 ( \41325 , \41324 );
xor \U$40983 ( \41326 , \41291 , \41310 );
and \U$40984 ( \41327 , \41326 , \41317 );
and \U$40985 ( \41328 , \41291 , \41310 );
or \U$40986 ( \41329 , \41327 , \41328 );
not \U$40987 ( \41330 , \41329 );
xor \U$40988 ( \41331 , \40151 , \40153 );
xor \U$40989 ( \41332 , \41331 , \40170 );
not \U$40990 ( \41333 , \41332 );
and \U$40991 ( \41334 , \41330 , \41333 );
and \U$40992 ( \41335 , \41329 , \41332 );
nor \U$40993 ( \41336 , \41334 , \41335 );
not \U$40994 ( \41337 , \41336 );
or \U$40995 ( \41338 , \41325 , \41337 );
or \U$40996 ( \41339 , \41336 , \41324 );
nand \U$40997 ( \41340 , \41338 , \41339 );
not \U$40998 ( \41341 , \41340 );
or \U$40999 ( \41342 , \41322 , \41341 );
or \U$41000 ( \41343 , \41340 , \41321 );
nand \U$41001 ( \41344 , \41342 , \41343 );
not \U$41002 ( \41345 , \41299 );
not \U$41003 ( \41346 , \41308 );
not \U$41004 ( \41347 , \41297 );
or \U$41005 ( \41348 , \41346 , \41347 );
or \U$41006 ( \41349 , \41297 , \41308 );
nand \U$41007 ( \41350 , \41348 , \41349 );
not \U$41008 ( \41351 , \41350 );
or \U$41009 ( \41352 , \41345 , \41351 );
or \U$41010 ( \41353 , \41350 , \41299 );
nand \U$41011 ( \41354 , \41352 , \41353 );
not \U$41012 ( \41355 , \41354 );
not \U$41013 ( \41356 , \40602 );
not \U$41014 ( \41357 , \41274 );
not \U$41015 ( \41358 , \41211 );
and \U$41016 ( \41359 , \41357 , \41358 );
and \U$41017 ( \41360 , \41274 , \41211 );
nor \U$41018 ( \41361 , \41359 , \41360 );
not \U$41019 ( \41362 , \41361 );
or \U$41020 ( \41363 , \41356 , \41362 );
or \U$41021 ( \41364 , \41361 , \40602 );
nand \U$41022 ( \41365 , \41363 , \41364 );
not \U$41023 ( \41366 , \41365 );
or \U$41024 ( \41367 , \41355 , \41366 );
or \U$41025 ( \41368 , \41365 , \41354 );
xor \U$41026 ( \41369 , \41145 , \41165 );
xor \U$41027 ( \41370 , \40814 , \41042 );
xor \U$41028 ( \41371 , \41370 , \41095 );
and \U$41029 ( \41372 , \41369 , \41371 );
xor \U$41030 ( \41373 , \41179 , \41189 );
xor \U$41031 ( \41374 , \41373 , \41205 );
xor \U$41032 ( \41375 , \40814 , \41042 );
xor \U$41033 ( \41376 , \41375 , \41095 );
and \U$41034 ( \41377 , \41374 , \41376 );
and \U$41035 ( \41378 , \41369 , \41374 );
or \U$41036 ( \41379 , \41372 , \41377 , \41378 );
xor \U$41037 ( \41380 , \40847 , \9510 );
xor \U$41038 ( \41381 , \41380 , \40855 );
xor \U$41039 ( \41382 , \40821 , \40829 );
xor \U$41040 ( \41383 , \41382 , \40837 );
and \U$41041 ( \41384 , \41381 , \41383 );
xor \U$41042 ( \41385 , \40866 , \40873 );
xor \U$41043 ( \41386 , \41385 , \40881 );
xor \U$41044 ( \41387 , \40821 , \40829 );
xor \U$41045 ( \41388 , \41387 , \40837 );
and \U$41046 ( \41389 , \41386 , \41388 );
and \U$41047 ( \41390 , \41381 , \41386 );
or \U$41048 ( \41391 , \41384 , \41389 , \41390 );
xor \U$41049 ( \41392 , \40917 , \40924 );
xor \U$41050 ( \41393 , \40895 , \40903 );
xor \U$41051 ( \41394 , \41393 , \40912 );
and \U$41052 ( \41395 , \41392 , \41394 );
xor \U$41053 ( \41396 , \40933 , \40940 );
xor \U$41054 ( \41397 , \41396 , \40949 );
xor \U$41055 ( \41398 , \40895 , \40903 );
xor \U$41056 ( \41399 , \41398 , \40912 );
and \U$41057 ( \41400 , \41397 , \41399 );
and \U$41058 ( \41401 , \41392 , \41397 );
or \U$41059 ( \41402 , \41395 , \41400 , \41401 );
xor \U$41060 ( \41403 , \41391 , \41402 );
xor \U$41061 ( \41404 , \41016 , \41024 );
xor \U$41062 ( \41405 , \41404 , \41033 );
xor \U$41063 ( \41406 , \40989 , \40997 );
xor \U$41064 ( \41407 , \41406 , \41005 );
xor \U$41065 ( \41408 , \41405 , \41407 );
xor \U$41066 ( \41409 , \40963 , \40971 );
xor \U$41067 ( \41410 , \41409 , \40979 );
and \U$41068 ( \41411 , \41408 , \41410 );
and \U$41069 ( \41412 , \41405 , \41407 );
or \U$41070 ( \41413 , \41411 , \41412 );
and \U$41071 ( \41414 , \41403 , \41413 );
and \U$41072 ( \41415 , \41391 , \41402 );
or \U$41073 ( \41416 , \41414 , \41415 );
and \U$41074 ( \41417 , \5318 , RI986f778_58);
and \U$41075 ( \41418 , RI986fa48_64, \5316 );
nor \U$41076 ( \41419 , \41417 , \41418 );
and \U$41077 ( \41420 , \41419 , \5052 );
not \U$41078 ( \41421 , \41419 );
and \U$41079 ( \41422 , \41421 , \5322 );
nor \U$41080 ( \41423 , \41420 , \41422 );
not \U$41081 ( \41424 , \4519 );
and \U$41082 ( \41425 , \4710 , RI986e698_22);
and \U$41083 ( \41426 , RI986f868_60, \4708 );
nor \U$41084 ( \41427 , \41425 , \41426 );
not \U$41085 ( \41428 , \41427 );
or \U$41086 ( \41429 , \41424 , \41428 );
or \U$41087 ( \41430 , \41427 , \4519 );
nand \U$41088 ( \41431 , \41429 , \41430 );
xor \U$41089 ( \41432 , \41423 , \41431 );
and \U$41090 ( \41433 , \5881 , RI986f958_62);
and \U$41091 ( \41434 , RI986f4a8_52, \5879 );
nor \U$41092 ( \41435 , \41433 , \41434 );
and \U$41093 ( \41436 , \41435 , \5594 );
not \U$41094 ( \41437 , \41435 );
and \U$41095 ( \41438 , \41437 , \5885 );
nor \U$41096 ( \41439 , \41436 , \41438 );
and \U$41097 ( \41440 , \41432 , \41439 );
and \U$41098 ( \41441 , \41423 , \41431 );
or \U$41099 ( \41442 , \41440 , \41441 );
and \U$41100 ( \41443 , \8486 , RI986dd38_2);
and \U$41101 ( \41444 , RI986e1e8_12, \8484 );
nor \U$41102 ( \41445 , \41443 , \41444 );
and \U$41103 ( \41446 , \41445 , \8050 );
not \U$41104 ( \41447 , \41445 );
and \U$41105 ( \41448 , \41447 , \8051 );
nor \U$41106 ( \41449 , \41446 , \41448 );
nand \U$41107 ( \41450 , RI986e3c8_16, \9505 );
and \U$41108 ( \41451 , \41450 , \9510 );
not \U$41109 ( \41452 , \41450 );
and \U$41110 ( \41453 , \41452 , \9513 );
nor \U$41111 ( \41454 , \41451 , \41453 );
xor \U$41112 ( \41455 , \41449 , \41454 );
and \U$41113 ( \41456 , \9237 , RI986e0f8_10);
and \U$41114 ( \41457 , RI986e2d8_14, \9235 );
nor \U$41115 ( \41458 , \41456 , \41457 );
and \U$41116 ( \41459 , \41458 , \9241 );
not \U$41117 ( \41460 , \41458 );
and \U$41118 ( \41461 , \41460 , \8836 );
nor \U$41119 ( \41462 , \41459 , \41461 );
and \U$41120 ( \41463 , \41455 , \41462 );
and \U$41121 ( \41464 , \41449 , \41454 );
or \U$41122 ( \41465 , \41463 , \41464 );
xor \U$41123 ( \41466 , \41442 , \41465 );
and \U$41124 ( \41467 , \7729 , RI986df18_6);
and \U$41125 ( \41468 , RI986de28_4, \7727 );
nor \U$41126 ( \41469 , \41467 , \41468 );
and \U$41127 ( \41470 , \41469 , \7480 );
not \U$41128 ( \41471 , \41469 );
and \U$41129 ( \41472 , \41471 , \7733 );
nor \U$41130 ( \41473 , \41470 , \41472 );
and \U$41131 ( \41474 , \6453 , RI986f3b8_50);
and \U$41132 ( \41475 , RI986f598_54, \6451 );
nor \U$41133 ( \41476 , \41474 , \41475 );
and \U$41134 ( \41477 , \41476 , \6190 );
not \U$41135 ( \41478 , \41476 );
and \U$41136 ( \41479 , \41478 , \6180 );
nor \U$41137 ( \41480 , \41477 , \41479 );
xor \U$41138 ( \41481 , \41473 , \41480 );
and \U$41139 ( \41482 , \7079 , RI986f688_56);
and \U$41140 ( \41483 , RI986e008_8, \7077 );
nor \U$41141 ( \41484 , \41482 , \41483 );
and \U$41142 ( \41485 , \41484 , \6710 );
not \U$41143 ( \41486 , \41484 );
and \U$41144 ( \41487 , \41486 , \6709 );
nor \U$41145 ( \41488 , \41485 , \41487 );
and \U$41146 ( \41489 , \41481 , \41488 );
and \U$41147 ( \41490 , \41473 , \41480 );
or \U$41148 ( \41491 , \41489 , \41490 );
and \U$41149 ( \41492 , \41466 , \41491 );
and \U$41150 ( \41493 , \41442 , \41465 );
or \U$41151 ( \41494 , \41492 , \41493 );
not \U$41152 ( \41495 , \345 );
and \U$41153 ( \41496 , \354 , RI9870b28_100);
and \U$41154 ( \41497 , RI9870df8_106, \352 );
nor \U$41155 ( \41498 , \41496 , \41497 );
not \U$41156 ( \41499 , \41498 );
or \U$41157 ( \41500 , \41495 , \41499 );
or \U$41158 ( \41501 , \41498 , \345 );
nand \U$41159 ( \41502 , \41500 , \41501 );
not \U$41160 ( \41503 , \365 );
and \U$41161 ( \41504 , \376 , RI9870c18_102);
and \U$41162 ( \41505 , RI98710c8_112, \374 );
nor \U$41163 ( \41506 , \41504 , \41505 );
not \U$41164 ( \41507 , \41506 );
or \U$41165 ( \41508 , \41503 , \41507 );
or \U$41166 ( \41509 , \41506 , \367 );
nand \U$41167 ( \41510 , \41508 , \41509 );
xor \U$41168 ( \41511 , \41502 , \41510 );
not \U$41169 ( \41512 , \386 );
and \U$41170 ( \41513 , \395 , RI9870a38_98);
and \U$41171 ( \41514 , RI9870ee8_108, \393 );
nor \U$41172 ( \41515 , \41513 , \41514 );
not \U$41173 ( \41516 , \41515 );
or \U$41174 ( \41517 , \41512 , \41516 );
or \U$41175 ( \41518 , \41515 , \386 );
nand \U$41176 ( \41519 , \41517 , \41518 );
and \U$41177 ( \41520 , \41511 , \41519 );
and \U$41178 ( \41521 , \41502 , \41510 );
or \U$41179 ( \41522 , \41520 , \41521 );
nand \U$41180 ( \41523 , RI98700d8_78, RI9871fc8_144);
and \U$41181 ( \41524 , \416 , RI98701c8_80);
and \U$41182 ( \41525 , RI9870fd8_110, \414 );
nor \U$41183 ( \41526 , \41524 , \41525 );
and \U$41184 ( \41527 , \41526 , \421 );
not \U$41185 ( \41528 , \41526 );
and \U$41186 ( \41529 , \41528 , \422 );
nor \U$41187 ( \41530 , \41527 , \41529 );
nand \U$41188 ( \41531 , \41523 , \41530 );
xor \U$41189 ( \41532 , \41522 , \41531 );
not \U$41190 ( \41533 , \456 );
and \U$41191 ( \41534 , \465 , RI9870d08_104);
and \U$41192 ( \41535 , RI98712a8_116, \463 );
nor \U$41193 ( \41536 , \41534 , \41535 );
not \U$41194 ( \41537 , \41536 );
or \U$41195 ( \41538 , \41533 , \41537 );
or \U$41196 ( \41539 , \41536 , \454 );
nand \U$41197 ( \41540 , \41538 , \41539 );
and \U$41198 ( \41541 , \776 , RI9871488_120);
and \U$41199 ( \41542 , RI9871758_126, \774 );
nor \U$41200 ( \41543 , \41541 , \41542 );
and \U$41201 ( \41544 , \41543 , \474 );
not \U$41202 ( \41545 , \41543 );
and \U$41203 ( \41546 , \41545 , \451 );
nor \U$41204 ( \41547 , \41544 , \41546 );
xor \U$41205 ( \41548 , \41540 , \41547 );
and \U$41206 ( \41549 , \438 , RI98711b8_114);
and \U$41207 ( \41550 , RI9871398_118, \436 );
nor \U$41208 ( \41551 , \41549 , \41550 );
and \U$41209 ( \41552 , \41551 , \444 );
not \U$41210 ( \41553 , \41551 );
and \U$41211 ( \41554 , \41553 , \443 );
nor \U$41212 ( \41555 , \41552 , \41554 );
and \U$41213 ( \41556 , \41548 , \41555 );
and \U$41214 ( \41557 , \41540 , \41547 );
or \U$41215 ( \41558 , \41556 , \41557 );
and \U$41216 ( \41559 , \41532 , \41558 );
and \U$41217 ( \41560 , \41522 , \41531 );
or \U$41218 ( \41561 , \41559 , \41560 );
xor \U$41219 ( \41562 , \41494 , \41561 );
not \U$41220 ( \41563 , \3412 );
and \U$41221 ( \41564 , \3683 , RI986f1d8_46);
and \U$41222 ( \41565 , RI986e5a8_20, \3681 );
nor \U$41223 ( \41566 , \41564 , \41565 );
not \U$41224 ( \41567 , \41566 );
or \U$41225 ( \41568 , \41563 , \41567 );
or \U$41226 ( \41569 , \41566 , \3918 );
nand \U$41227 ( \41570 , \41568 , \41569 );
not \U$41228 ( \41571 , \2935 );
and \U$41229 ( \41572 , \3254 , RI986eff8_42);
and \U$41230 ( \41573 , RI986f2c8_48, \3252 );
nor \U$41231 ( \41574 , \41572 , \41573 );
not \U$41232 ( \41575 , \41574 );
or \U$41233 ( \41576 , \41571 , \41575 );
or \U$41234 ( \41577 , \41574 , \2935 );
nand \U$41235 ( \41578 , \41576 , \41577 );
xor \U$41236 ( \41579 , \41570 , \41578 );
and \U$41237 ( \41580 , \4203 , RI986e4b8_18);
and \U$41238 ( \41581 , RI986e788_24, \4201 );
nor \U$41239 ( \41582 , \41580 , \41581 );
and \U$41240 ( \41583 , \41582 , \4207 );
not \U$41241 ( \41584 , \41582 );
and \U$41242 ( \41585 , \41584 , \3923 );
nor \U$41243 ( \41586 , \41583 , \41585 );
and \U$41244 ( \41587 , \41579 , \41586 );
and \U$41245 ( \41588 , \41570 , \41578 );
or \U$41246 ( \41589 , \41587 , \41588 );
not \U$41247 ( \41590 , \2034 );
and \U$41248 ( \41591 , \2042 , RI986e878_26);
and \U$41249 ( \41592 , RI986ef08_40, \2040 );
nor \U$41250 ( \41593 , \41591 , \41592 );
not \U$41251 ( \41594 , \41593 );
or \U$41252 ( \41595 , \41590 , \41594 );
or \U$41253 ( \41596 , \41593 , \2034 );
nand \U$41254 ( \41597 , \41595 , \41596 );
and \U$41255 ( \41598 , \2274 , RI986ee18_38);
and \U$41256 ( \41599 , RI986ec38_34, \2272 );
nor \U$41257 ( \41600 , \41598 , \41599 );
and \U$41258 ( \41601 , \41600 , \2030 );
not \U$41259 ( \41602 , \41600 );
and \U$41260 ( \41603 , \41602 , \2031 );
nor \U$41261 ( \41604 , \41601 , \41603 );
xor \U$41262 ( \41605 , \41597 , \41604 );
and \U$41263 ( \41606 , \2464 , RI986ed28_36);
and \U$41264 ( \41607 , RI986f0e8_44, \2462 );
nor \U$41265 ( \41608 , \41606 , \41607 );
and \U$41266 ( \41609 , \41608 , \2468 );
not \U$41267 ( \41610 , \41608 );
and \U$41268 ( \41611 , \41610 , \2263 );
nor \U$41269 ( \41612 , \41609 , \41611 );
and \U$41270 ( \41613 , \41605 , \41612 );
and \U$41271 ( \41614 , \41597 , \41604 );
or \U$41272 ( \41615 , \41613 , \41614 );
xor \U$41273 ( \41616 , \41589 , \41615 );
and \U$41274 ( \41617 , \1311 , RI986ea58_30);
and \U$41275 ( \41618 , RI986e968_28, \1309 );
nor \U$41276 ( \41619 , \41617 , \41618 );
and \U$41277 ( \41620 , \41619 , \1458 );
not \U$41278 ( \41621 , \41619 );
and \U$41279 ( \41622 , \41621 , \1318 );
nor \U$41280 ( \41623 , \41620 , \41622 );
not \U$41281 ( \41624 , \1128 );
and \U$41282 ( \41625 , \1293 , RI9871848_128);
and \U$41283 ( \41626 , RI9871578_122, \1291 );
nor \U$41284 ( \41627 , \41625 , \41626 );
not \U$41285 ( \41628 , \41627 );
or \U$41286 ( \41629 , \41624 , \41628 );
or \U$41287 ( \41630 , \41627 , \1301 );
nand \U$41288 ( \41631 , \41629 , \41630 );
xor \U$41289 ( \41632 , \41623 , \41631 );
and \U$41290 ( \41633 , \1329 , RI9871668_124);
and \U$41291 ( \41634 , RI986eb48_32, \1327 );
nor \U$41292 ( \41635 , \41633 , \41634 );
and \U$41293 ( \41636 , \41635 , \1336 );
not \U$41294 ( \41637 , \41635 );
and \U$41295 ( \41638 , \41637 , \1337 );
nor \U$41296 ( \41639 , \41636 , \41638 );
and \U$41297 ( \41640 , \41632 , \41639 );
and \U$41298 ( \41641 , \41623 , \41631 );
or \U$41299 ( \41642 , \41640 , \41641 );
and \U$41300 ( \41643 , \41616 , \41642 );
and \U$41301 ( \41644 , \41589 , \41615 );
or \U$41302 ( \41645 , \41643 , \41644 );
and \U$41303 ( \41646 , \41562 , \41645 );
and \U$41304 ( \41647 , \41494 , \41561 );
or \U$41305 ( \41648 , \41646 , \41647 );
xor \U$41306 ( \41649 , \41416 , \41648 );
xor \U$41307 ( \41650 , \40763 , \40771 );
xor \U$41308 ( \41651 , \41650 , \40779 );
xor \U$41309 ( \41652 , \40756 , \40806 );
xor \U$41310 ( \41653 , \41651 , \41652 );
xor \U$41311 ( \41654 , \40701 , \40702 );
xor \U$41312 ( \41655 , \41654 , \40728 );
and \U$41313 ( \41656 , \41653 , \41655 );
xor \U$41314 ( \41657 , \40631 , \40638 );
xor \U$41315 ( \41658 , \41657 , \40646 );
xor \U$41316 ( \41659 , \40623 , \40671 );
xor \U$41317 ( \41660 , \41658 , \41659 );
xor \U$41318 ( \41661 , \40701 , \40702 );
xor \U$41319 ( \41662 , \41661 , \40728 );
and \U$41320 ( \41663 , \41660 , \41662 );
and \U$41321 ( \41664 , \41653 , \41660 );
or \U$41322 ( \41665 , \41656 , \41663 , \41664 );
and \U$41323 ( \41666 , \41649 , \41665 );
and \U$41324 ( \41667 , \41416 , \41648 );
or \U$41325 ( \41668 , \41666 , \41667 );
xor \U$41326 ( \41669 , \40887 , \40955 );
xor \U$41327 ( \41670 , \41669 , \41039 );
xor \U$41328 ( \41671 , \40676 , \40731 );
xor \U$41329 ( \41672 , \41671 , \40811 );
and \U$41330 ( \41673 , \41670 , \41672 );
xor \U$41331 ( \41674 , \41668 , \41673 );
xor \U$41332 ( \41675 , \40840 , \40858 );
xor \U$41333 ( \41676 , \41675 , \40884 );
xor \U$41334 ( \41677 , \40982 , \41008 );
xor \U$41335 ( \41678 , \41677 , \41036 );
xor \U$41336 ( \41679 , \41676 , \41678 );
xor \U$41337 ( \41680 , \40915 , \40925 );
xor \U$41338 ( \41681 , \41680 , \40952 );
and \U$41339 ( \41682 , \41679 , \41681 );
and \U$41340 ( \41683 , \41676 , \41678 );
or \U$41341 ( \41684 , \41682 , \41683 );
xor \U$41342 ( \41685 , \41181 , \41183 );
xor \U$41343 ( \41686 , \41685 , \41186 );
and \U$41344 ( \41687 , \41684 , \41686 );
xor \U$41345 ( \41688 , \41063 , \41065 );
xor \U$41346 ( \41689 , \41688 , \41072 );
xor \U$41347 ( \41690 , \41054 , \41090 );
xor \U$41348 ( \41691 , \41689 , \41690 );
xor \U$41349 ( \41692 , \41181 , \41183 );
xor \U$41350 ( \41693 , \41692 , \41186 );
and \U$41351 ( \41694 , \41691 , \41693 );
and \U$41352 ( \41695 , \41684 , \41691 );
or \U$41353 ( \41696 , \41687 , \41694 , \41695 );
and \U$41354 ( \41697 , \41674 , \41696 );
and \U$41355 ( \41698 , \41668 , \41673 );
or \U$41356 ( \41699 , \41697 , \41698 );
and \U$41357 ( \41700 , \41379 , \41699 );
not \U$41358 ( \41701 , \41379 );
not \U$41359 ( \41702 , \41699 );
and \U$41360 ( \41703 , \41701 , \41702 );
xor \U$41361 ( \41704 , \41234 , \41238 );
xor \U$41362 ( \41705 , \41704 , \41245 );
xor \U$41363 ( \41706 , \41228 , \41269 );
xor \U$41364 ( \41707 , \41705 , \41706 );
nor \U$41365 ( \41708 , \41703 , \41707 );
nor \U$41366 ( \41709 , \41700 , \41708 );
not \U$41367 ( \41710 , \41709 );
nand \U$41368 ( \41711 , \41368 , \41710 );
nand \U$41369 ( \41712 , \41367 , \41711 );
not \U$41370 ( \41713 , \41712 );
xor \U$41371 ( \41714 , \41276 , \41286 );
xor \U$41372 ( \41715 , \41714 , \41318 );
nor \U$41373 ( \41716 , \41713 , \41715 );
and \U$41374 ( \41717 , \41344 , \41716 );
xor \U$41375 ( \41718 , \41716 , \41344 );
not \U$41376 ( \41719 , \41715 );
not \U$41377 ( \41720 , \41712 );
and \U$41378 ( \41721 , \41719 , \41720 );
and \U$41379 ( \41722 , \41715 , \41712 );
nor \U$41380 ( \41723 , \41721 , \41722 );
not \U$41381 ( \41724 , \41709 );
not \U$41382 ( \41725 , \41354 );
and \U$41383 ( \41726 , \41724 , \41725 );
and \U$41384 ( \41727 , \41709 , \41354 );
nor \U$41385 ( \41728 , \41726 , \41727 );
not \U$41386 ( \41729 , \41728 );
not \U$41387 ( \41730 , \41365 );
and \U$41388 ( \41731 , \41729 , \41730 );
and \U$41389 ( \41732 , \41728 , \41365 );
nor \U$41390 ( \41733 , \41731 , \41732 );
not \U$41391 ( \41734 , \41733 );
not \U$41392 ( \41735 , \41707 );
xor \U$41393 ( \41736 , \41699 , \41379 );
not \U$41394 ( \41737 , \41736 );
or \U$41395 ( \41738 , \41735 , \41737 );
or \U$41396 ( \41739 , \41736 , \41707 );
nand \U$41397 ( \41740 , \41738 , \41739 );
xor \U$41398 ( \41741 , \41098 , \41166 );
xor \U$41399 ( \41742 , \41741 , \41208 );
xor \U$41400 ( \41743 , \41740 , \41742 );
xor \U$41401 ( \41744 , \41449 , \41454 );
xor \U$41402 ( \41745 , \41744 , \41462 );
xor \U$41403 ( \41746 , \41423 , \41431 );
xor \U$41404 ( \41747 , \41746 , \41439 );
and \U$41405 ( \41748 , \41745 , \41747 );
xor \U$41406 ( \41749 , \41473 , \41480 );
xor \U$41407 ( \41750 , \41749 , \41488 );
xor \U$41408 ( \41751 , \41423 , \41431 );
xor \U$41409 ( \41752 , \41751 , \41439 );
and \U$41410 ( \41753 , \41750 , \41752 );
and \U$41411 ( \41754 , \41745 , \41750 );
or \U$41412 ( \41755 , \41748 , \41753 , \41754 );
xor \U$41413 ( \41756 , \41540 , \41547 );
xor \U$41414 ( \41757 , \41756 , \41555 );
or \U$41415 ( \41758 , \41530 , \41523 );
nand \U$41416 ( \41759 , \41758 , \41531 );
xor \U$41417 ( \41760 , \41757 , \41759 );
xor \U$41418 ( \41761 , \41502 , \41510 );
xor \U$41419 ( \41762 , \41761 , \41519 );
and \U$41420 ( \41763 , \41760 , \41762 );
and \U$41421 ( \41764 , \41757 , \41759 );
or \U$41422 ( \41765 , \41763 , \41764 );
xor \U$41423 ( \41766 , \41755 , \41765 );
xor \U$41424 ( \41767 , \41623 , \41631 );
xor \U$41425 ( \41768 , \41767 , \41639 );
xor \U$41426 ( \41769 , \41597 , \41604 );
xor \U$41427 ( \41770 , \41769 , \41612 );
and \U$41428 ( \41771 , \41768 , \41770 );
xor \U$41429 ( \41772 , \41570 , \41578 );
xor \U$41430 ( \41773 , \41772 , \41586 );
xor \U$41431 ( \41774 , \41597 , \41604 );
xor \U$41432 ( \41775 , \41774 , \41612 );
and \U$41433 ( \41776 , \41773 , \41775 );
and \U$41434 ( \41777 , \41768 , \41773 );
or \U$41435 ( \41778 , \41771 , \41776 , \41777 );
and \U$41436 ( \41779 , \41766 , \41778 );
and \U$41437 ( \41780 , \41755 , \41765 );
or \U$41438 ( \41781 , \41779 , \41780 );
and \U$41439 ( \41782 , \6453 , RI986f4a8_52);
and \U$41440 ( \41783 , RI986f3b8_50, \6451 );
nor \U$41441 ( \41784 , \41782 , \41783 );
and \U$41442 ( \41785 , \41784 , \6190 );
not \U$41443 ( \41786 , \41784 );
and \U$41444 ( \41787 , \41786 , \6705 );
nor \U$41445 ( \41788 , \41785 , \41787 );
and \U$41446 ( \41789 , \5318 , RI986f868_60);
and \U$41447 ( \41790 , RI986f778_58, \5316 );
nor \U$41448 ( \41791 , \41789 , \41790 );
and \U$41449 ( \41792 , \41791 , \5052 );
not \U$41450 ( \41793 , \41791 );
and \U$41451 ( \41794 , \41793 , \5322 );
nor \U$41452 ( \41795 , \41792 , \41794 );
xor \U$41453 ( \41796 , \41788 , \41795 );
and \U$41454 ( \41797 , \5881 , RI986fa48_64);
and \U$41455 ( \41798 , RI986f958_62, \5879 );
nor \U$41456 ( \41799 , \41797 , \41798 );
and \U$41457 ( \41800 , \41799 , \5594 );
not \U$41458 ( \41801 , \41799 );
and \U$41459 ( \41802 , \41801 , \5885 );
nor \U$41460 ( \41803 , \41800 , \41802 );
and \U$41461 ( \41804 , \41796 , \41803 );
and \U$41462 ( \41805 , \41788 , \41795 );
or \U$41463 ( \41806 , \41804 , \41805 );
and \U$41464 ( \41807 , \9505 , RI986e2d8_14);
and \U$41465 ( \41808 , RI986e3c8_16, \9503 );
nor \U$41466 ( \41809 , \41807 , \41808 );
and \U$41467 ( \41810 , \41809 , \9510 );
not \U$41468 ( \41811 , \41809 );
and \U$41469 ( \41812 , \41811 , \9513 );
nor \U$41470 ( \41813 , \41810 , \41812 );
xor \U$41471 ( \41814 , \41813 , \9840 );
and \U$41472 ( \41815 , \9237 , RI986e1e8_12);
and \U$41473 ( \41816 , RI986e0f8_10, \9235 );
nor \U$41474 ( \41817 , \41815 , \41816 );
and \U$41475 ( \41818 , \41817 , \9241 );
not \U$41476 ( \41819 , \41817 );
and \U$41477 ( \41820 , \41819 , \8836 );
nor \U$41478 ( \41821 , \41818 , \41820 );
and \U$41479 ( \41822 , \41814 , \41821 );
and \U$41480 ( \41823 , \41813 , \9840 );
or \U$41481 ( \41824 , \41822 , \41823 );
xor \U$41482 ( \41825 , \41806 , \41824 );
and \U$41483 ( \41826 , \7079 , RI986f598_54);
and \U$41484 ( \41827 , RI986f688_56, \7077 );
nor \U$41485 ( \41828 , \41826 , \41827 );
and \U$41486 ( \41829 , \41828 , \6710 );
not \U$41487 ( \41830 , \41828 );
and \U$41488 ( \41831 , \41830 , \6709 );
nor \U$41489 ( \41832 , \41829 , \41831 );
and \U$41490 ( \41833 , \7729 , RI986e008_8);
and \U$41491 ( \41834 , RI986df18_6, \7727 );
nor \U$41492 ( \41835 , \41833 , \41834 );
and \U$41493 ( \41836 , \41835 , \7480 );
not \U$41494 ( \41837 , \41835 );
and \U$41495 ( \41838 , \41837 , \7733 );
nor \U$41496 ( \41839 , \41836 , \41838 );
xor \U$41497 ( \41840 , \41832 , \41839 );
and \U$41498 ( \41841 , \8486 , RI986de28_4);
and \U$41499 ( \41842 , RI986dd38_2, \8484 );
nor \U$41500 ( \41843 , \41841 , \41842 );
and \U$41501 ( \41844 , \41843 , \8050 );
not \U$41502 ( \41845 , \41843 );
and \U$41503 ( \41846 , \41845 , \8051 );
nor \U$41504 ( \41847 , \41844 , \41846 );
and \U$41505 ( \41848 , \41840 , \41847 );
and \U$41506 ( \41849 , \41832 , \41839 );
or \U$41507 ( \41850 , \41848 , \41849 );
and \U$41508 ( \41851 , \41825 , \41850 );
and \U$41509 ( \41852 , \41806 , \41824 );
or \U$41510 ( \41853 , \41851 , \41852 );
not \U$41511 ( \41854 , \454 );
and \U$41512 ( \41855 , \465 , RI98710c8_112);
and \U$41513 ( \41856 , RI9870d08_104, \463 );
nor \U$41514 ( \41857 , \41855 , \41856 );
not \U$41515 ( \41858 , \41857 );
or \U$41516 ( \41859 , \41854 , \41858 );
or \U$41517 ( \41860 , \41857 , \456 );
nand \U$41518 ( \41861 , \41859 , \41860 );
not \U$41519 ( \41862 , \365 );
and \U$41520 ( \41863 , \376 , RI9870ee8_108);
and \U$41521 ( \41864 , RI9870c18_102, \374 );
nor \U$41522 ( \41865 , \41863 , \41864 );
not \U$41523 ( \41866 , \41865 );
or \U$41524 ( \41867 , \41862 , \41866 );
or \U$41525 ( \41868 , \41865 , \365 );
nand \U$41526 ( \41869 , \41867 , \41868 );
xor \U$41527 ( \41870 , \41861 , \41869 );
not \U$41528 ( \41871 , \386 );
and \U$41529 ( \41872 , \395 , RI9870df8_106);
and \U$41530 ( \41873 , RI9870a38_98, \393 );
nor \U$41531 ( \41874 , \41872 , \41873 );
not \U$41532 ( \41875 , \41874 );
or \U$41533 ( \41876 , \41871 , \41875 );
or \U$41534 ( \41877 , \41874 , \386 );
nand \U$41535 ( \41878 , \41876 , \41877 );
and \U$41536 ( \41879 , \41870 , \41878 );
and \U$41537 ( \41880 , \41861 , \41869 );
or \U$41538 ( \41881 , \41879 , \41880 );
and \U$41539 ( \41882 , \416 , RI98700d8_78);
and \U$41540 ( \41883 , RI98701c8_80, \414 );
nor \U$41541 ( \41884 , \41882 , \41883 );
and \U$41542 ( \41885 , \41884 , \422 );
not \U$41543 ( \41886 , \41884 );
and \U$41544 ( \41887 , \41886 , \421 );
nor \U$41545 ( \41888 , \41885 , \41887 );
not \U$41546 ( \41889 , RI986fef8_74);
nor \U$41547 ( \41890 , \41889 , \407 );
xor \U$41548 ( \41891 , \41888 , \41890 );
not \U$41549 ( \41892 , \345 );
and \U$41550 ( \41893 , \354 , RI9870fd8_110);
and \U$41551 ( \41894 , RI9870b28_100, \352 );
nor \U$41552 ( \41895 , \41893 , \41894 );
not \U$41553 ( \41896 , \41895 );
or \U$41554 ( \41897 , \41892 , \41896 );
or \U$41555 ( \41898 , \41895 , \361 );
nand \U$41556 ( \41899 , \41897 , \41898 );
and \U$41557 ( \41900 , \41891 , \41899 );
and \U$41558 ( \41901 , \41888 , \41890 );
or \U$41559 ( \41902 , \41900 , \41901 );
xor \U$41560 ( \41903 , \41881 , \41902 );
and \U$41561 ( \41904 , \438 , RI98712a8_116);
and \U$41562 ( \41905 , RI98711b8_114, \436 );
nor \U$41563 ( \41906 , \41904 , \41905 );
and \U$41564 ( \41907 , \41906 , \444 );
not \U$41565 ( \41908 , \41906 );
and \U$41566 ( \41909 , \41908 , \443 );
nor \U$41567 ( \41910 , \41907 , \41909 );
and \U$41568 ( \41911 , \776 , RI9871398_118);
and \U$41569 ( \41912 , RI9871488_120, \774 );
nor \U$41570 ( \41913 , \41911 , \41912 );
and \U$41571 ( \41914 , \41913 , \474 );
not \U$41572 ( \41915 , \41913 );
and \U$41573 ( \41916 , \41915 , \451 );
nor \U$41574 ( \41917 , \41914 , \41916 );
xor \U$41575 ( \41918 , \41910 , \41917 );
not \U$41576 ( \41919 , \1128 );
and \U$41577 ( \41920 , \1293 , RI9871758_126);
and \U$41578 ( \41921 , RI9871848_128, \1291 );
nor \U$41579 ( \41922 , \41920 , \41921 );
not \U$41580 ( \41923 , \41922 );
or \U$41581 ( \41924 , \41919 , \41923 );
or \U$41582 ( \41925 , \41922 , \1128 );
nand \U$41583 ( \41926 , \41924 , \41925 );
and \U$41584 ( \41927 , \41918 , \41926 );
and \U$41585 ( \41928 , \41910 , \41917 );
or \U$41586 ( \41929 , \41927 , \41928 );
and \U$41587 ( \41930 , \41903 , \41929 );
and \U$41588 ( \41931 , \41881 , \41902 );
or \U$41589 ( \41932 , \41930 , \41931 );
xor \U$41590 ( \41933 , \41853 , \41932 );
and \U$41591 ( \41934 , \2274 , RI986ef08_40);
and \U$41592 ( \41935 , RI986ee18_38, \2272 );
nor \U$41593 ( \41936 , \41934 , \41935 );
and \U$41594 ( \41937 , \41936 , \2030 );
not \U$41595 ( \41938 , \41936 );
and \U$41596 ( \41939 , \41938 , \2031 );
nor \U$41597 ( \41940 , \41937 , \41939 );
and \U$41598 ( \41941 , \2464 , RI986ec38_34);
and \U$41599 ( \41942 , RI986ed28_36, \2462 );
nor \U$41600 ( \41943 , \41941 , \41942 );
and \U$41601 ( \41944 , \41943 , \2468 );
not \U$41602 ( \41945 , \41943 );
and \U$41603 ( \41946 , \41945 , \2263 );
nor \U$41604 ( \41947 , \41944 , \41946 );
xor \U$41605 ( \41948 , \41940 , \41947 );
not \U$41606 ( \41949 , \3406 );
and \U$41607 ( \41950 , \3254 , RI986f0e8_44);
and \U$41608 ( \41951 , RI986eff8_42, \3252 );
nor \U$41609 ( \41952 , \41950 , \41951 );
not \U$41610 ( \41953 , \41952 );
or \U$41611 ( \41954 , \41949 , \41953 );
or \U$41612 ( \41955 , \41952 , \3406 );
nand \U$41613 ( \41956 , \41954 , \41955 );
and \U$41614 ( \41957 , \41948 , \41956 );
and \U$41615 ( \41958 , \41940 , \41947 );
or \U$41616 ( \41959 , \41957 , \41958 );
not \U$41617 ( \41960 , \2034 );
and \U$41618 ( \41961 , \2042 , RI986e968_28);
and \U$41619 ( \41962 , RI986e878_26, \2040 );
nor \U$41620 ( \41963 , \41961 , \41962 );
not \U$41621 ( \41964 , \41963 );
or \U$41622 ( \41965 , \41960 , \41964 );
or \U$41623 ( \41966 , \41963 , \1462 );
nand \U$41624 ( \41967 , \41965 , \41966 );
and \U$41625 ( \41968 , \1329 , RI9871578_122);
and \U$41626 ( \41969 , RI9871668_124, \1327 );
nor \U$41627 ( \41970 , \41968 , \41969 );
and \U$41628 ( \41971 , \41970 , \1336 );
not \U$41629 ( \41972 , \41970 );
and \U$41630 ( \41973 , \41972 , \1337 );
nor \U$41631 ( \41974 , \41971 , \41973 );
xor \U$41632 ( \41975 , \41967 , \41974 );
and \U$41633 ( \41976 , \1311 , RI986eb48_32);
and \U$41634 ( \41977 , RI986ea58_30, \1309 );
nor \U$41635 ( \41978 , \41976 , \41977 );
and \U$41636 ( \41979 , \41978 , \1458 );
not \U$41637 ( \41980 , \41978 );
and \U$41638 ( \41981 , \41980 , \1318 );
nor \U$41639 ( \41982 , \41979 , \41981 );
and \U$41640 ( \41983 , \41975 , \41982 );
and \U$41641 ( \41984 , \41967 , \41974 );
or \U$41642 ( \41985 , \41983 , \41984 );
xor \U$41643 ( \41986 , \41959 , \41985 );
not \U$41644 ( \41987 , \4519 );
and \U$41645 ( \41988 , \4710 , RI986e788_24);
and \U$41646 ( \41989 , RI986e698_22, \4708 );
nor \U$41647 ( \41990 , \41988 , \41989 );
not \U$41648 ( \41991 , \41990 );
or \U$41649 ( \41992 , \41987 , \41991 );
or \U$41650 ( \41993 , \41990 , \4519 );
nand \U$41651 ( \41994 , \41992 , \41993 );
not \U$41652 ( \41995 , \3412 );
and \U$41653 ( \41996 , \3683 , RI986f2c8_48);
and \U$41654 ( \41997 , RI986f1d8_46, \3681 );
nor \U$41655 ( \41998 , \41996 , \41997 );
not \U$41656 ( \41999 , \41998 );
or \U$41657 ( \42000 , \41995 , \41999 );
or \U$41658 ( \42001 , \41998 , \3918 );
nand \U$41659 ( \42002 , \42000 , \42001 );
xor \U$41660 ( \42003 , \41994 , \42002 );
and \U$41661 ( \42004 , \4203 , RI986e5a8_20);
and \U$41662 ( \42005 , RI986e4b8_18, \4201 );
nor \U$41663 ( \42006 , \42004 , \42005 );
and \U$41664 ( \42007 , \42006 , \4207 );
not \U$41665 ( \42008 , \42006 );
and \U$41666 ( \42009 , \42008 , \3923 );
nor \U$41667 ( \42010 , \42007 , \42009 );
and \U$41668 ( \42011 , \42003 , \42010 );
and \U$41669 ( \42012 , \41994 , \42002 );
or \U$41670 ( \42013 , \42011 , \42012 );
and \U$41671 ( \42014 , \41986 , \42013 );
and \U$41672 ( \42015 , \41959 , \41985 );
or \U$41673 ( \42016 , \42014 , \42015 );
and \U$41674 ( \42017 , \41933 , \42016 );
and \U$41675 ( \42018 , \41853 , \41932 );
or \U$41676 ( \42019 , \42017 , \42018 );
xor \U$41677 ( \42020 , \41781 , \42019 );
xor \U$41678 ( \42021 , \40895 , \40903 );
xor \U$41679 ( \42022 , \42021 , \40912 );
xor \U$41680 ( \42023 , \41392 , \41397 );
xor \U$41681 ( \42024 , \42022 , \42023 );
xor \U$41682 ( \42025 , \41405 , \41407 );
xor \U$41683 ( \42026 , \42025 , \41410 );
and \U$41684 ( \42027 , \42024 , \42026 );
xor \U$41685 ( \42028 , \40821 , \40829 );
xor \U$41686 ( \42029 , \42028 , \40837 );
xor \U$41687 ( \42030 , \41381 , \41386 );
xor \U$41688 ( \42031 , \42029 , \42030 );
xor \U$41689 ( \42032 , \41405 , \41407 );
xor \U$41690 ( \42033 , \42032 , \41410 );
and \U$41691 ( \42034 , \42031 , \42033 );
and \U$41692 ( \42035 , \42024 , \42031 );
or \U$41693 ( \42036 , \42027 , \42034 , \42035 );
and \U$41694 ( \42037 , \42020 , \42036 );
and \U$41695 ( \42038 , \41781 , \42019 );
or \U$41696 ( \42039 , \42037 , \42038 );
xor \U$41697 ( \42040 , \41494 , \41561 );
xor \U$41698 ( \42041 , \42040 , \41645 );
xor \U$41699 ( \42042 , \41391 , \41402 );
xor \U$41700 ( \42043 , \42042 , \41413 );
and \U$41701 ( \42044 , \42041 , \42043 );
xor \U$41702 ( \42045 , \42039 , \42044 );
xor \U$41703 ( \42046 , \41589 , \41615 );
xor \U$41704 ( \42047 , \42046 , \41642 );
xor \U$41705 ( \42048 , \41522 , \41531 );
xor \U$41706 ( \42049 , \42048 , \41558 );
xor \U$41707 ( \42050 , \42047 , \42049 );
xor \U$41708 ( \42051 , \41442 , \41465 );
xor \U$41709 ( \42052 , \42051 , \41491 );
and \U$41710 ( \42053 , \42050 , \42052 );
and \U$41711 ( \42054 , \42047 , \42049 );
or \U$41712 ( \42055 , \42053 , \42054 );
xor \U$41713 ( \42056 , \41676 , \41678 );
xor \U$41714 ( \42057 , \42056 , \41681 );
and \U$41715 ( \42058 , \42055 , \42057 );
xor \U$41716 ( \42059 , \40701 , \40702 );
xor \U$41717 ( \42060 , \42059 , \40728 );
xor \U$41718 ( \42061 , \41653 , \41660 );
xor \U$41719 ( \42062 , \42060 , \42061 );
xor \U$41720 ( \42063 , \41676 , \41678 );
xor \U$41721 ( \42064 , \42063 , \41681 );
and \U$41722 ( \42065 , \42062 , \42064 );
and \U$41723 ( \42066 , \42055 , \42062 );
or \U$41724 ( \42067 , \42058 , \42065 , \42066 );
and \U$41725 ( \42068 , \42045 , \42067 );
and \U$41726 ( \42069 , \42039 , \42044 );
or \U$41727 ( \42070 , \42068 , \42069 );
xor \U$41728 ( \42071 , \41670 , \41672 );
xor \U$41729 ( \42072 , \41416 , \41648 );
xor \U$41730 ( \42073 , \42072 , \41665 );
and \U$41731 ( \42074 , \42071 , \42073 );
xor \U$41732 ( \42075 , \41181 , \41183 );
xor \U$41733 ( \42076 , \42075 , \41186 );
xor \U$41734 ( \42077 , \41684 , \41691 );
xor \U$41735 ( \42078 , \42076 , \42077 );
xor \U$41736 ( \42079 , \41416 , \41648 );
xor \U$41737 ( \42080 , \42079 , \41665 );
and \U$41738 ( \42081 , \42078 , \42080 );
and \U$41739 ( \42082 , \42071 , \42078 );
or \U$41740 ( \42083 , \42074 , \42081 , \42082 );
xor \U$41741 ( \42084 , \42070 , \42083 );
xor \U$41742 ( \42085 , \40814 , \41042 );
xor \U$41743 ( \42086 , \42085 , \41095 );
xor \U$41744 ( \42087 , \41369 , \41374 );
xor \U$41745 ( \42088 , \42086 , \42087 );
and \U$41746 ( \42089 , \42084 , \42088 );
and \U$41747 ( \42090 , \42070 , \42083 );
or \U$41748 ( \42091 , \42089 , \42090 );
and \U$41749 ( \42092 , \41743 , \42091 );
and \U$41750 ( \42093 , \41740 , \41742 );
or \U$41751 ( \42094 , \42092 , \42093 );
nand \U$41752 ( \42095 , \41734 , \42094 );
or \U$41753 ( \42096 , \41723 , \42095 );
xnor \U$41754 ( \42097 , \42095 , \41723 );
not \U$41755 ( \42098 , \3412 );
and \U$41756 ( \42099 , \3683 , RI986eff8_42);
and \U$41757 ( \42100 , RI986f2c8_48, \3681 );
nor \U$41758 ( \42101 , \42099 , \42100 );
not \U$41759 ( \42102 , \42101 );
or \U$41760 ( \42103 , \42098 , \42102 );
or \U$41761 ( \42104 , \42101 , \3918 );
nand \U$41762 ( \42105 , \42103 , \42104 );
and \U$41763 ( \42106 , \4203 , RI986f1d8_46);
and \U$41764 ( \42107 , RI986e5a8_20, \4201 );
nor \U$41765 ( \42108 , \42106 , \42107 );
and \U$41766 ( \42109 , \42108 , \4207 );
not \U$41767 ( \42110 , \42108 );
and \U$41768 ( \42111 , \42110 , \3922 );
nor \U$41769 ( \42112 , \42109 , \42111 );
xor \U$41770 ( \42113 , \42105 , \42112 );
not \U$41771 ( \42114 , \4519 );
and \U$41772 ( \42115 , \4710 , RI986e4b8_18);
and \U$41773 ( \42116 , RI986e788_24, \4708 );
nor \U$41774 ( \42117 , \42115 , \42116 );
not \U$41775 ( \42118 , \42117 );
or \U$41776 ( \42119 , \42114 , \42118 );
or \U$41777 ( \42120 , \42117 , \4521 );
nand \U$41778 ( \42121 , \42119 , \42120 );
xor \U$41779 ( \42122 , \42113 , \42121 );
and \U$41780 ( \42123 , \7079 , RI986f3b8_50);
and \U$41781 ( \42124 , RI986f598_54, \7077 );
nor \U$41782 ( \42125 , \42123 , \42124 );
and \U$41783 ( \42126 , \42125 , \6710 );
not \U$41784 ( \42127 , \42125 );
and \U$41785 ( \42128 , \42127 , \6709 );
nor \U$41786 ( \42129 , \42126 , \42128 );
and \U$41787 ( \42130 , \7729 , RI986f688_56);
and \U$41788 ( \42131 , RI986e008_8, \7727 );
nor \U$41789 ( \42132 , \42130 , \42131 );
and \U$41790 ( \42133 , \42132 , \7480 );
not \U$41791 ( \42134 , \42132 );
and \U$41792 ( \42135 , \42134 , \7733 );
nor \U$41793 ( \42136 , \42133 , \42135 );
xor \U$41794 ( \42137 , \42129 , \42136 );
and \U$41795 ( \42138 , \8486 , RI986df18_6);
and \U$41796 ( \42139 , RI986de28_4, \8484 );
nor \U$41797 ( \42140 , \42138 , \42139 );
and \U$41798 ( \42141 , \42140 , \8050 );
not \U$41799 ( \42142 , \42140 );
and \U$41800 ( \42143 , \42142 , \8051 );
nor \U$41801 ( \42144 , \42141 , \42143 );
xor \U$41802 ( \42145 , \42137 , \42144 );
and \U$41803 ( \42146 , \42122 , \42145 );
and \U$41804 ( \42147 , \5318 , RI986e698_22);
and \U$41805 ( \42148 , RI986f868_60, \5316 );
nor \U$41806 ( \42149 , \42147 , \42148 );
and \U$41807 ( \42150 , \42149 , \5052 );
not \U$41808 ( \42151 , \42149 );
and \U$41809 ( \42152 , \42151 , \5322 );
nor \U$41810 ( \42153 , \42150 , \42152 );
and \U$41811 ( \42154 , \5881 , RI986f778_58);
and \U$41812 ( \42155 , RI986fa48_64, \5879 );
nor \U$41813 ( \42156 , \42154 , \42155 );
and \U$41814 ( \42157 , \42156 , \5594 );
not \U$41815 ( \42158 , \42156 );
and \U$41816 ( \42159 , \42158 , \5885 );
nor \U$41817 ( \42160 , \42157 , \42159 );
xor \U$41818 ( \42161 , \42153 , \42160 );
and \U$41819 ( \42162 , \6453 , RI986f958_62);
and \U$41820 ( \42163 , RI986f4a8_52, \6451 );
nor \U$41821 ( \42164 , \42162 , \42163 );
and \U$41822 ( \42165 , \42164 , \6190 );
not \U$41823 ( \42166 , \42164 );
and \U$41824 ( \42167 , \42166 , \6705 );
nor \U$41825 ( \42168 , \42165 , \42167 );
xor \U$41826 ( \42169 , \42161 , \42168 );
xor \U$41827 ( \42170 , \42129 , \42136 );
xor \U$41828 ( \42171 , \42170 , \42144 );
and \U$41829 ( \42172 , \42169 , \42171 );
and \U$41830 ( \42173 , \42122 , \42169 );
or \U$41831 ( \42174 , \42146 , \42172 , \42173 );
and \U$41832 ( \42175 , \354 , RI98701c8_80);
and \U$41833 ( \42176 , RI9870fd8_110, \352 );
nor \U$41834 ( \42177 , \42175 , \42176 );
not \U$41835 ( \42178 , \42177 );
not \U$41836 ( \42179 , \345 );
and \U$41837 ( \42180 , \42178 , \42179 );
and \U$41838 ( \42181 , \42177 , \345 );
nor \U$41839 ( \42182 , \42180 , \42181 );
not \U$41840 ( \42183 , \42182 );
and \U$41841 ( \42184 , \416 , RI986fef8_74);
and \U$41842 ( \42185 , RI98700d8_78, \414 );
nor \U$41843 ( \42186 , \42184 , \42185 );
and \U$41844 ( \42187 , \42186 , \422 );
not \U$41845 ( \42188 , \42186 );
and \U$41846 ( \42189 , \42188 , \421 );
nor \U$41847 ( \42190 , \42187 , \42189 );
not \U$41848 ( \42191 , \42190 );
or \U$41849 ( \42192 , \42183 , \42191 );
or \U$41850 ( \42193 , \42182 , \42190 );
nand \U$41851 ( \42194 , \42192 , \42193 );
not \U$41852 ( \42195 , \42194 );
nand \U$41853 ( \42196 , RI986ffe8_76, RI9871fc8_144);
not \U$41854 ( \42197 , \42196 );
and \U$41855 ( \42198 , \42195 , \42197 );
and \U$41856 ( \42199 , \42194 , \42196 );
nor \U$41857 ( \42200 , \42198 , \42199 );
and \U$41858 ( \42201 , \376 , RI9870a38_98);
and \U$41859 ( \42202 , RI9870ee8_108, \374 );
nor \U$41860 ( \42203 , \42201 , \42202 );
not \U$41861 ( \42204 , \42203 );
not \U$41862 ( \42205 , \365 );
and \U$41863 ( \42206 , \42204 , \42205 );
and \U$41864 ( \42207 , \42203 , \367 );
nor \U$41865 ( \42208 , \42206 , \42207 );
not \U$41866 ( \42209 , \42208 );
not \U$41867 ( \42210 , \454 );
and \U$41868 ( \42211 , \465 , RI9870c18_102);
and \U$41869 ( \42212 , RI98710c8_112, \463 );
nor \U$41870 ( \42213 , \42211 , \42212 );
not \U$41871 ( \42214 , \42213 );
or \U$41872 ( \42215 , \42210 , \42214 );
or \U$41873 ( \42216 , \42213 , \454 );
nand \U$41874 ( \42217 , \42215 , \42216 );
not \U$41875 ( \42218 , \42217 );
or \U$41876 ( \42219 , \42209 , \42218 );
or \U$41877 ( \42220 , \42208 , \42217 );
nand \U$41878 ( \42221 , \42219 , \42220 );
not \U$41879 ( \42222 , \42221 );
and \U$41880 ( \42223 , \395 , RI9870b28_100);
and \U$41881 ( \42224 , RI9870df8_106, \393 );
nor \U$41882 ( \42225 , \42223 , \42224 );
not \U$41883 ( \42226 , \42225 );
not \U$41884 ( \42227 , \487 );
and \U$41885 ( \42228 , \42226 , \42227 );
and \U$41886 ( \42229 , \42225 , \386 );
nor \U$41887 ( \42230 , \42228 , \42229 );
not \U$41888 ( \42231 , \42230 );
and \U$41889 ( \42232 , \42222 , \42231 );
and \U$41890 ( \42233 , \42221 , \42230 );
nor \U$41891 ( \42234 , \42232 , \42233 );
nand \U$41892 ( \42235 , \42200 , \42234 );
xor \U$41893 ( \42236 , \42174 , \42235 );
and \U$41894 ( \42237 , \2274 , RI986e878_26);
and \U$41895 ( \42238 , RI986ef08_40, \2272 );
nor \U$41896 ( \42239 , \42237 , \42238 );
and \U$41897 ( \42240 , \42239 , \2030 );
not \U$41898 ( \42241 , \42239 );
and \U$41899 ( \42242 , \42241 , \2031 );
nor \U$41900 ( \42243 , \42240 , \42242 );
and \U$41901 ( \42244 , \2464 , RI986ee18_38);
and \U$41902 ( \42245 , RI986ec38_34, \2462 );
nor \U$41903 ( \42246 , \42244 , \42245 );
and \U$41904 ( \42247 , \42246 , \2468 );
not \U$41905 ( \42248 , \42246 );
and \U$41906 ( \42249 , \42248 , \2263 );
nor \U$41907 ( \42250 , \42247 , \42249 );
xor \U$41908 ( \42251 , \42243 , \42250 );
not \U$41909 ( \42252 , \2935 );
and \U$41910 ( \42253 , \3254 , RI986ed28_36);
and \U$41911 ( \42254 , RI986f0e8_44, \3252 );
nor \U$41912 ( \42255 , \42253 , \42254 );
not \U$41913 ( \42256 , \42255 );
or \U$41914 ( \42257 , \42252 , \42256 );
or \U$41915 ( \42258 , \42255 , \3406 );
nand \U$41916 ( \42259 , \42257 , \42258 );
xor \U$41917 ( \42260 , \42251 , \42259 );
not \U$41918 ( \42261 , \1301 );
and \U$41919 ( \42262 , \1293 , RI9871488_120);
and \U$41920 ( \42263 , RI9871758_126, \1291 );
nor \U$41921 ( \42264 , \42262 , \42263 );
not \U$41922 ( \42265 , \42264 );
or \U$41923 ( \42266 , \42261 , \42265 );
or \U$41924 ( \42267 , \42264 , \1301 );
nand \U$41925 ( \42268 , \42266 , \42267 );
and \U$41926 ( \42269 , \776 , RI98711b8_114);
and \U$41927 ( \42270 , RI9871398_118, \774 );
nor \U$41928 ( \42271 , \42269 , \42270 );
and \U$41929 ( \42272 , \42271 , \474 );
not \U$41930 ( \42273 , \42271 );
and \U$41931 ( \42274 , \42273 , \451 );
nor \U$41932 ( \42275 , \42272 , \42274 );
xor \U$41933 ( \42276 , \42268 , \42275 );
and \U$41934 ( \42277 , \438 , RI9870d08_104);
and \U$41935 ( \42278 , RI98712a8_116, \436 );
nor \U$41936 ( \42279 , \42277 , \42278 );
and \U$41937 ( \42280 , \42279 , \444 );
not \U$41938 ( \42281 , \42279 );
and \U$41939 ( \42282 , \42281 , \443 );
nor \U$41940 ( \42283 , \42280 , \42282 );
xor \U$41941 ( \42284 , \42276 , \42283 );
xor \U$41942 ( \42285 , \42260 , \42284 );
not \U$41943 ( \42286 , \1462 );
and \U$41944 ( \42287 , \2042 , RI986ea58_30);
and \U$41945 ( \42288 , RI986e968_28, \2040 );
nor \U$41946 ( \42289 , \42287 , \42288 );
not \U$41947 ( \42290 , \42289 );
or \U$41948 ( \42291 , \42286 , \42290 );
or \U$41949 ( \42292 , \42289 , \2034 );
nand \U$41950 ( \42293 , \42291 , \42292 );
and \U$41951 ( \42294 , \1329 , RI9871848_128);
and \U$41952 ( \42295 , RI9871578_122, \1327 );
nor \U$41953 ( \42296 , \42294 , \42295 );
and \U$41954 ( \42297 , \42296 , \1336 );
not \U$41955 ( \42298 , \42296 );
and \U$41956 ( \42299 , \42298 , \1337 );
nor \U$41957 ( \42300 , \42297 , \42299 );
xor \U$41958 ( \42301 , \42293 , \42300 );
and \U$41959 ( \42302 , \1311 , RI9871668_124);
and \U$41960 ( \42303 , RI986eb48_32, \1309 );
nor \U$41961 ( \42304 , \42302 , \42303 );
and \U$41962 ( \42305 , \42304 , \1458 );
not \U$41963 ( \42306 , \42304 );
and \U$41964 ( \42307 , \42306 , \1315 );
nor \U$41965 ( \42308 , \42305 , \42307 );
xor \U$41966 ( \42309 , \42301 , \42308 );
and \U$41967 ( \42310 , \42285 , \42309 );
and \U$41968 ( \42311 , \42260 , \42284 );
or \U$41969 ( \42312 , \42310 , \42311 );
and \U$41970 ( \42313 , \42236 , \42312 );
and \U$41971 ( \42314 , \42174 , \42235 );
or \U$41972 ( \42315 , \42313 , \42314 );
not \U$41973 ( \42316 , \487 );
and \U$41974 ( \42317 , \395 , RI9870fd8_110);
and \U$41975 ( \42318 , RI9870b28_100, \393 );
nor \U$41976 ( \42319 , \42317 , \42318 );
not \U$41977 ( \42320 , \42319 );
or \U$41978 ( \42321 , \42316 , \42320 );
or \U$41979 ( \42322 , \42319 , \487 );
nand \U$41980 ( \42323 , \42321 , \42322 );
not \U$41981 ( \42324 , \361 );
and \U$41982 ( \42325 , \354 , RI98700d8_78);
and \U$41983 ( \42326 , RI98701c8_80, \352 );
nor \U$41984 ( \42327 , \42325 , \42326 );
not \U$41985 ( \42328 , \42327 );
or \U$41986 ( \42329 , \42324 , \42328 );
or \U$41987 ( \42330 , \42327 , \345 );
nand \U$41988 ( \42331 , \42329 , \42330 );
xor \U$41989 ( \42332 , \42323 , \42331 );
and \U$41990 ( \42333 , \416 , RI986ffe8_76);
and \U$41991 ( \42334 , RI986fef8_74, \414 );
nor \U$41992 ( \42335 , \42333 , \42334 );
and \U$41993 ( \42336 , \42335 , \422 );
not \U$41994 ( \42337 , \42335 );
and \U$41995 ( \42338 , \42337 , \421 );
nor \U$41996 ( \42339 , \42336 , \42338 );
and \U$41997 ( \42340 , \42332 , \42339 );
and \U$41998 ( \42341 , \42323 , \42331 );
or \U$41999 ( \42342 , \42340 , \42341 );
and \U$42000 ( \42343 , \438 , RI98710c8_112);
and \U$42001 ( \42344 , RI9870d08_104, \436 );
nor \U$42002 ( \42345 , \42343 , \42344 );
and \U$42003 ( \42346 , \42345 , \444 );
not \U$42004 ( \42347 , \42345 );
and \U$42005 ( \42348 , \42347 , \443 );
nor \U$42006 ( \42349 , \42346 , \42348 );
not \U$42007 ( \42350 , \454 );
and \U$42008 ( \42351 , \465 , RI9870ee8_108);
and \U$42009 ( \42352 , RI9870c18_102, \463 );
nor \U$42010 ( \42353 , \42351 , \42352 );
not \U$42011 ( \42354 , \42353 );
or \U$42012 ( \42355 , \42350 , \42354 );
or \U$42013 ( \42356 , \42353 , \456 );
nand \U$42014 ( \42357 , \42355 , \42356 );
xor \U$42015 ( \42358 , \42349 , \42357 );
not \U$42016 ( \42359 , \367 );
and \U$42017 ( \42360 , \376 , RI9870df8_106);
and \U$42018 ( \42361 , RI9870a38_98, \374 );
nor \U$42019 ( \42362 , \42360 , \42361 );
not \U$42020 ( \42363 , \42362 );
or \U$42021 ( \42364 , \42359 , \42363 );
or \U$42022 ( \42365 , \42362 , \365 );
nand \U$42023 ( \42366 , \42364 , \42365 );
and \U$42024 ( \42367 , \42358 , \42366 );
and \U$42025 ( \42368 , \42349 , \42357 );
or \U$42026 ( \42369 , \42367 , \42368 );
xor \U$42027 ( \42370 , \42342 , \42369 );
not \U$42028 ( \42371 , \1301 );
and \U$42029 ( \42372 , \1293 , RI9871398_118);
and \U$42030 ( \42373 , RI9871488_120, \1291 );
nor \U$42031 ( \42374 , \42372 , \42373 );
not \U$42032 ( \42375 , \42374 );
or \U$42033 ( \42376 , \42371 , \42375 );
or \U$42034 ( \42377 , \42374 , \1128 );
nand \U$42035 ( \42378 , \42376 , \42377 );
and \U$42036 ( \42379 , \776 , RI98712a8_116);
and \U$42037 ( \42380 , RI98711b8_114, \774 );
nor \U$42038 ( \42381 , \42379 , \42380 );
and \U$42039 ( \42382 , \42381 , \474 );
not \U$42040 ( \42383 , \42381 );
and \U$42041 ( \42384 , \42383 , \451 );
nor \U$42042 ( \42385 , \42382 , \42384 );
xor \U$42043 ( \42386 , \42378 , \42385 );
and \U$42044 ( \42387 , \1329 , RI9871758_126);
and \U$42045 ( \42388 , RI9871848_128, \1327 );
nor \U$42046 ( \42389 , \42387 , \42388 );
and \U$42047 ( \42390 , \42389 , \1336 );
not \U$42048 ( \42391 , \42389 );
and \U$42049 ( \42392 , \42391 , \1337 );
nor \U$42050 ( \42393 , \42390 , \42392 );
and \U$42051 ( \42394 , \42386 , \42393 );
and \U$42052 ( \42395 , \42378 , \42385 );
or \U$42053 ( \42396 , \42394 , \42395 );
and \U$42054 ( \42397 , \42370 , \42396 );
and \U$42055 ( \42398 , \42342 , \42369 );
or \U$42056 ( \42399 , \42397 , \42398 );
and \U$42057 ( \42400 , \9237 , RI986de28_4);
and \U$42058 ( \42401 , RI986dd38_2, \9235 );
nor \U$42059 ( \42402 , \42400 , \42401 );
and \U$42060 ( \42403 , \42402 , \9241 );
not \U$42061 ( \42404 , \42402 );
and \U$42062 ( \42405 , \42404 , \8836 );
nor \U$42063 ( \42406 , \42403 , \42405 );
and \U$42064 ( \42407 , \7729 , RI986f598_54);
and \U$42065 ( \42408 , RI986f688_56, \7727 );
nor \U$42066 ( \42409 , \42407 , \42408 );
and \U$42067 ( \42410 , \42409 , \7480 );
not \U$42068 ( \42411 , \42409 );
and \U$42069 ( \42412 , \42411 , \7733 );
nor \U$42070 ( \42413 , \42410 , \42412 );
xor \U$42071 ( \42414 , \42406 , \42413 );
and \U$42072 ( \42415 , \8486 , RI986e008_8);
and \U$42073 ( \42416 , RI986df18_6, \8484 );
nor \U$42074 ( \42417 , \42415 , \42416 );
and \U$42075 ( \42418 , \42417 , \8050 );
not \U$42076 ( \42419 , \42417 );
and \U$42077 ( \42420 , \42419 , \8051 );
nor \U$42078 ( \42421 , \42418 , \42420 );
and \U$42079 ( \42422 , \42414 , \42421 );
and \U$42080 ( \42423 , \42406 , \42413 );
or \U$42081 ( \42424 , \42422 , \42423 );
and \U$42082 ( \42425 , \9505 , RI986e1e8_12);
and \U$42083 ( \42426 , RI986e0f8_10, \9503 );
nor \U$42084 ( \42427 , \42425 , \42426 );
and \U$42085 ( \42428 , \42427 , \9510 );
not \U$42086 ( \42429 , \42427 );
and \U$42087 ( \42430 , \42429 , \9513 );
nor \U$42088 ( \42431 , \42428 , \42430 );
xor \U$42089 ( \42432 , \42431 , \10965 );
and \U$42090 ( \42433 , \10424 , RI986e2d8_14);
and \U$42091 ( \42434 , RI986e3c8_16, \10422 );
nor \U$42092 ( \42435 , \42433 , \42434 );
and \U$42093 ( \42436 , \42435 , \9840 );
not \U$42094 ( \42437 , \42435 );
and \U$42095 ( \42438 , \42437 , \10428 );
nor \U$42096 ( \42439 , \42436 , \42438 );
and \U$42097 ( \42440 , \42432 , \42439 );
and \U$42098 ( \42441 , \42431 , \10965 );
or \U$42099 ( \42442 , \42440 , \42441 );
xor \U$42100 ( \42443 , \42424 , \42442 );
and \U$42101 ( \42444 , \5881 , RI986f868_60);
and \U$42102 ( \42445 , RI986f778_58, \5879 );
nor \U$42103 ( \42446 , \42444 , \42445 );
and \U$42104 ( \42447 , \42446 , \5594 );
not \U$42105 ( \42448 , \42446 );
and \U$42106 ( \42449 , \42448 , \5885 );
nor \U$42107 ( \42450 , \42447 , \42449 );
and \U$42108 ( \42451 , \6453 , RI986fa48_64);
and \U$42109 ( \42452 , RI986f958_62, \6451 );
nor \U$42110 ( \42453 , \42451 , \42452 );
and \U$42111 ( \42454 , \42453 , \6190 );
not \U$42112 ( \42455 , \42453 );
and \U$42113 ( \42456 , \42455 , \6705 );
nor \U$42114 ( \42457 , \42454 , \42456 );
xor \U$42115 ( \42458 , \42450 , \42457 );
and \U$42116 ( \42459 , \7079 , RI986f4a8_52);
and \U$42117 ( \42460 , RI986f3b8_50, \7077 );
nor \U$42118 ( \42461 , \42459 , \42460 );
and \U$42119 ( \42462 , \42461 , \6710 );
not \U$42120 ( \42463 , \42461 );
and \U$42121 ( \42464 , \42463 , \6709 );
nor \U$42122 ( \42465 , \42462 , \42464 );
and \U$42123 ( \42466 , \42458 , \42465 );
and \U$42124 ( \42467 , \42450 , \42457 );
or \U$42125 ( \42468 , \42466 , \42467 );
and \U$42126 ( \42469 , \42443 , \42468 );
and \U$42127 ( \42470 , \42424 , \42442 );
or \U$42128 ( \42471 , \42469 , \42470 );
xor \U$42129 ( \42472 , \42399 , \42471 );
and \U$42130 ( \42473 , \5318 , RI986e788_24);
and \U$42131 ( \42474 , RI986e698_22, \5316 );
nor \U$42132 ( \42475 , \42473 , \42474 );
and \U$42133 ( \42476 , \42475 , \5052 );
not \U$42134 ( \42477 , \42475 );
and \U$42135 ( \42478 , \42477 , \5322 );
nor \U$42136 ( \42479 , \42476 , \42478 );
and \U$42137 ( \42480 , \4203 , RI986f2c8_48);
and \U$42138 ( \42481 , RI986f1d8_46, \4201 );
nor \U$42139 ( \42482 , \42480 , \42481 );
and \U$42140 ( \42483 , \42482 , \4207 );
not \U$42141 ( \42484 , \42482 );
and \U$42142 ( \42485 , \42484 , \3922 );
nor \U$42143 ( \42486 , \42483 , \42485 );
xor \U$42144 ( \42487 , \42479 , \42486 );
not \U$42145 ( \42488 , \4521 );
and \U$42146 ( \42489 , \4710 , RI986e5a8_20);
and \U$42147 ( \42490 , RI986e4b8_18, \4708 );
nor \U$42148 ( \42491 , \42489 , \42490 );
not \U$42149 ( \42492 , \42491 );
or \U$42150 ( \42493 , \42488 , \42492 );
or \U$42151 ( \42494 , \42491 , \4519 );
nand \U$42152 ( \42495 , \42493 , \42494 );
and \U$42153 ( \42496 , \42487 , \42495 );
and \U$42154 ( \42497 , \42479 , \42486 );
or \U$42155 ( \42498 , \42496 , \42497 );
not \U$42156 ( \42499 , \3918 );
and \U$42157 ( \42500 , \3683 , RI986f0e8_44);
and \U$42158 ( \42501 , RI986eff8_42, \3681 );
nor \U$42159 ( \42502 , \42500 , \42501 );
not \U$42160 ( \42503 , \42502 );
or \U$42161 ( \42504 , \42499 , \42503 );
or \U$42162 ( \42505 , \42502 , \3918 );
nand \U$42163 ( \42506 , \42504 , \42505 );
and \U$42164 ( \42507 , \2464 , RI986ef08_40);
and \U$42165 ( \42508 , RI986ee18_38, \2462 );
nor \U$42166 ( \42509 , \42507 , \42508 );
and \U$42167 ( \42510 , \42509 , \2468 );
not \U$42168 ( \42511 , \42509 );
and \U$42169 ( \42512 , \42511 , \2263 );
nor \U$42170 ( \42513 , \42510 , \42512 );
xor \U$42171 ( \42514 , \42506 , \42513 );
not \U$42172 ( \42515 , \3406 );
and \U$42173 ( \42516 , \3254 , RI986ec38_34);
and \U$42174 ( \42517 , RI986ed28_36, \3252 );
nor \U$42175 ( \42518 , \42516 , \42517 );
not \U$42176 ( \42519 , \42518 );
or \U$42177 ( \42520 , \42515 , \42519 );
or \U$42178 ( \42521 , \42518 , \3406 );
nand \U$42179 ( \42522 , \42520 , \42521 );
and \U$42180 ( \42523 , \42514 , \42522 );
and \U$42181 ( \42524 , \42506 , \42513 );
or \U$42182 ( \42525 , \42523 , \42524 );
xor \U$42183 ( \42526 , \42498 , \42525 );
and \U$42184 ( \42527 , \2274 , RI986e968_28);
and \U$42185 ( \42528 , RI986e878_26, \2272 );
nor \U$42186 ( \42529 , \42527 , \42528 );
and \U$42187 ( \42530 , \42529 , \2030 );
not \U$42188 ( \42531 , \42529 );
and \U$42189 ( \42532 , \42531 , \2031 );
nor \U$42190 ( \42533 , \42530 , \42532 );
and \U$42191 ( \42534 , \1311 , RI9871578_122);
and \U$42192 ( \42535 , RI9871668_124, \1309 );
nor \U$42193 ( \42536 , \42534 , \42535 );
and \U$42194 ( \42537 , \42536 , \1458 );
not \U$42195 ( \42538 , \42536 );
and \U$42196 ( \42539 , \42538 , \1318 );
nor \U$42197 ( \42540 , \42537 , \42539 );
xor \U$42198 ( \42541 , \42533 , \42540 );
not \U$42199 ( \42542 , \2034 );
and \U$42200 ( \42543 , \2042 , RI986eb48_32);
and \U$42201 ( \42544 , RI986ea58_30, \2040 );
nor \U$42202 ( \42545 , \42543 , \42544 );
not \U$42203 ( \42546 , \42545 );
or \U$42204 ( \42547 , \42542 , \42546 );
or \U$42205 ( \42548 , \42545 , \2034 );
nand \U$42206 ( \42549 , \42547 , \42548 );
and \U$42207 ( \42550 , \42541 , \42549 );
and \U$42208 ( \42551 , \42533 , \42540 );
or \U$42209 ( \42552 , \42550 , \42551 );
and \U$42210 ( \42553 , \42526 , \42552 );
and \U$42211 ( \42554 , \42498 , \42525 );
or \U$42212 ( \42555 , \42553 , \42554 );
and \U$42213 ( \42556 , \42472 , \42555 );
and \U$42214 ( \42557 , \42399 , \42471 );
or \U$42215 ( \42558 , \42556 , \42557 );
xor \U$42216 ( \42559 , \42315 , \42558 );
xor \U$42217 ( \42560 , \41861 , \41869 );
xor \U$42218 ( \42561 , \42560 , \41878 );
xor \U$42219 ( \42562 , \41888 , \41890 );
xor \U$42220 ( \42563 , \42562 , \41899 );
xor \U$42221 ( \42564 , \41910 , \41917 );
xor \U$42222 ( \42565 , \42564 , \41926 );
xor \U$42223 ( \42566 , \42563 , \42565 );
xor \U$42224 ( \42567 , \42561 , \42566 );
xor \U$42225 ( \42568 , \41940 , \41947 );
xor \U$42226 ( \42569 , \42568 , \41956 );
xor \U$42227 ( \42570 , \41967 , \41974 );
xor \U$42228 ( \42571 , \42570 , \41982 );
xor \U$42229 ( \42572 , \42569 , \42571 );
xor \U$42230 ( \42573 , \41994 , \42002 );
xor \U$42231 ( \42574 , \42573 , \42010 );
xor \U$42232 ( \42575 , \42572 , \42574 );
and \U$42233 ( \42576 , \42567 , \42575 );
xor \U$42234 ( \42577 , \41788 , \41795 );
xor \U$42235 ( \42578 , \42577 , \41803 );
xor \U$42236 ( \42579 , \41813 , \9840 );
xor \U$42237 ( \42580 , \42579 , \41821 );
xor \U$42238 ( \42581 , \41832 , \41839 );
xor \U$42239 ( \42582 , \42581 , \41847 );
xor \U$42240 ( \42583 , \42580 , \42582 );
xor \U$42241 ( \42584 , \42578 , \42583 );
xor \U$42242 ( \42585 , \42569 , \42571 );
xor \U$42243 ( \42586 , \42585 , \42574 );
and \U$42244 ( \42587 , \42584 , \42586 );
and \U$42245 ( \42588 , \42567 , \42584 );
or \U$42246 ( \42589 , \42576 , \42587 , \42588 );
and \U$42247 ( \42590 , \42559 , \42589 );
and \U$42248 ( \42591 , \42315 , \42558 );
or \U$42249 ( \42592 , \42590 , \42591 );
xor \U$42250 ( \42593 , \42105 , \42112 );
and \U$42251 ( \42594 , \42593 , \42121 );
and \U$42252 ( \42595 , \42105 , \42112 );
or \U$42253 ( \42596 , \42594 , \42595 );
xor \U$42254 ( \42597 , \42243 , \42250 );
and \U$42255 ( \42598 , \42597 , \42259 );
and \U$42256 ( \42599 , \42243 , \42250 );
or \U$42257 ( \42600 , \42598 , \42599 );
xor \U$42258 ( \42601 , \42596 , \42600 );
xor \U$42259 ( \42602 , \42293 , \42300 );
and \U$42260 ( \42603 , \42602 , \42308 );
and \U$42261 ( \42604 , \42293 , \42300 );
or \U$42262 ( \42605 , \42603 , \42604 );
and \U$42263 ( \42606 , \42601 , \42605 );
and \U$42264 ( \42607 , \42596 , \42600 );
or \U$42265 ( \42608 , \42606 , \42607 );
or \U$42266 ( \42609 , \42208 , \42230 );
not \U$42267 ( \42610 , \42230 );
not \U$42268 ( \42611 , \42208 );
or \U$42269 ( \42612 , \42610 , \42611 );
nand \U$42270 ( \42613 , \42612 , \42217 );
nand \U$42271 ( \42614 , \42609 , \42613 );
or \U$42272 ( \42615 , \42182 , \42196 );
not \U$42273 ( \42616 , \42196 );
not \U$42274 ( \42617 , \42182 );
or \U$42275 ( \42618 , \42616 , \42617 );
nand \U$42276 ( \42619 , \42618 , \42190 );
nand \U$42277 ( \42620 , \42615 , \42619 );
xor \U$42278 ( \42621 , \42614 , \42620 );
xor \U$42279 ( \42622 , \42268 , \42275 );
and \U$42280 ( \42623 , \42622 , \42283 );
and \U$42281 ( \42624 , \42268 , \42275 );
or \U$42282 ( \42625 , \42623 , \42624 );
and \U$42283 ( \42626 , \42621 , \42625 );
and \U$42284 ( \42627 , \42614 , \42620 );
or \U$42285 ( \42628 , \42626 , \42627 );
xor \U$42286 ( \42629 , \42608 , \42628 );
xor \U$42287 ( \42630 , \42153 , \42160 );
and \U$42288 ( \42631 , \42630 , \42168 );
and \U$42289 ( \42632 , \42153 , \42160 );
or \U$42290 ( \42633 , \42631 , \42632 );
and \U$42291 ( \42634 , \9237 , RI986dd38_2);
and \U$42292 ( \42635 , RI986e1e8_12, \9235 );
nor \U$42293 ( \42636 , \42634 , \42635 );
and \U$42294 ( \42637 , \42636 , \9241 );
not \U$42295 ( \42638 , \42636 );
and \U$42296 ( \42639 , \42638 , \8836 );
nor \U$42297 ( \42640 , \42637 , \42639 );
nand \U$42298 ( \42641 , RI986e3c8_16, \10424 );
and \U$42299 ( \42642 , \42641 , \9840 );
not \U$42300 ( \42643 , \42641 );
and \U$42301 ( \42644 , \42643 , \10428 );
nor \U$42302 ( \42645 , \42642 , \42644 );
xor \U$42303 ( \42646 , \42640 , \42645 );
and \U$42304 ( \42647 , \9505 , RI986e0f8_10);
and \U$42305 ( \42648 , RI986e2d8_14, \9503 );
nor \U$42306 ( \42649 , \42647 , \42648 );
and \U$42307 ( \42650 , \42649 , \9510 );
not \U$42308 ( \42651 , \42649 );
and \U$42309 ( \42652 , \42651 , \9513 );
nor \U$42310 ( \42653 , \42650 , \42652 );
and \U$42311 ( \42654 , \42646 , \42653 );
and \U$42312 ( \42655 , \42640 , \42645 );
or \U$42313 ( \42656 , \42654 , \42655 );
xor \U$42314 ( \42657 , \42633 , \42656 );
xor \U$42315 ( \42658 , \42129 , \42136 );
and \U$42316 ( \42659 , \42658 , \42144 );
and \U$42317 ( \42660 , \42129 , \42136 );
or \U$42318 ( \42661 , \42659 , \42660 );
and \U$42319 ( \42662 , \42657 , \42661 );
and \U$42320 ( \42663 , \42633 , \42656 );
or \U$42321 ( \42664 , \42662 , \42663 );
xor \U$42322 ( \42665 , \42629 , \42664 );
xor \U$42323 ( \42666 , \41788 , \41795 );
xor \U$42324 ( \42667 , \42666 , \41803 );
and \U$42325 ( \42668 , \42580 , \42667 );
xor \U$42326 ( \42669 , \41788 , \41795 );
xor \U$42327 ( \42670 , \42669 , \41803 );
and \U$42328 ( \42671 , \42582 , \42670 );
and \U$42329 ( \42672 , \42580 , \42582 );
or \U$42330 ( \42673 , \42668 , \42671 , \42672 );
xor \U$42331 ( \42674 , \41861 , \41869 );
xor \U$42332 ( \42675 , \42674 , \41878 );
and \U$42333 ( \42676 , \42563 , \42675 );
xor \U$42334 ( \42677 , \41861 , \41869 );
xor \U$42335 ( \42678 , \42677 , \41878 );
and \U$42336 ( \42679 , \42565 , \42678 );
and \U$42337 ( \42680 , \42563 , \42565 );
or \U$42338 ( \42681 , \42676 , \42679 , \42680 );
xor \U$42339 ( \42682 , \42673 , \42681 );
xor \U$42340 ( \42683 , \42569 , \42571 );
and \U$42341 ( \42684 , \42683 , \42574 );
and \U$42342 ( \42685 , \42569 , \42571 );
or \U$42343 ( \42686 , \42684 , \42685 );
xor \U$42344 ( \42687 , \42682 , \42686 );
and \U$42345 ( \42688 , \42665 , \42687 );
xor \U$42346 ( \42689 , \42592 , \42688 );
xor \U$42347 ( \42690 , \42596 , \42600 );
xor \U$42348 ( \42691 , \42690 , \42605 );
xor \U$42349 ( \42692 , \42633 , \42656 );
xor \U$42350 ( \42693 , \42692 , \42661 );
xor \U$42351 ( \42694 , \42691 , \42693 );
xor \U$42352 ( \42695 , \42614 , \42620 );
xor \U$42353 ( \42696 , \42695 , \42625 );
and \U$42354 ( \42697 , \42694 , \42696 );
and \U$42355 ( \42698 , \42691 , \42693 );
or \U$42356 ( \42699 , \42697 , \42698 );
xor \U$42357 ( \42700 , \41881 , \41902 );
xor \U$42358 ( \42701 , \42700 , \41929 );
xor \U$42359 ( \42702 , \41806 , \41824 );
xor \U$42360 ( \42703 , \42702 , \41850 );
xor \U$42361 ( \42704 , \42701 , \42703 );
xor \U$42362 ( \42705 , \41959 , \41985 );
xor \U$42363 ( \42706 , \42705 , \42013 );
xor \U$42364 ( \42707 , \42704 , \42706 );
and \U$42365 ( \42708 , \42699 , \42707 );
xor \U$42366 ( \42709 , \41757 , \41759 );
xor \U$42367 ( \42710 , \42709 , \41762 );
xor \U$42368 ( \42711 , \41423 , \41431 );
xor \U$42369 ( \42712 , \42711 , \41439 );
xor \U$42370 ( \42713 , \41745 , \41750 );
xor \U$42371 ( \42714 , \42712 , \42713 );
xor \U$42372 ( \42715 , \41597 , \41604 );
xor \U$42373 ( \42716 , \42715 , \41612 );
xor \U$42374 ( \42717 , \41768 , \41773 );
xor \U$42375 ( \42718 , \42716 , \42717 );
xor \U$42376 ( \42719 , \42714 , \42718 );
xor \U$42377 ( \42720 , \42710 , \42719 );
xor \U$42378 ( \42721 , \42701 , \42703 );
xor \U$42379 ( \42722 , \42721 , \42706 );
and \U$42380 ( \42723 , \42720 , \42722 );
and \U$42381 ( \42724 , \42699 , \42720 );
or \U$42382 ( \42725 , \42708 , \42723 , \42724 );
and \U$42383 ( \42726 , \42689 , \42725 );
and \U$42384 ( \42727 , \42592 , \42688 );
or \U$42385 ( \42728 , \42726 , \42727 );
xor \U$42386 ( \42729 , \41853 , \41932 );
xor \U$42387 ( \42730 , \42729 , \42016 );
xor \U$42388 ( \42731 , \41755 , \41765 );
xor \U$42389 ( \42732 , \42731 , \41778 );
xor \U$42390 ( \42733 , \42730 , \42732 );
xor \U$42391 ( \42734 , \42673 , \42681 );
and \U$42392 ( \42735 , \42734 , \42686 );
and \U$42393 ( \42736 , \42673 , \42681 );
or \U$42394 ( \42737 , \42735 , \42736 );
xor \U$42395 ( \42738 , \42608 , \42628 );
and \U$42396 ( \42739 , \42738 , \42664 );
and \U$42397 ( \42740 , \42608 , \42628 );
or \U$42398 ( \42741 , \42739 , \42740 );
xor \U$42399 ( \42742 , \42737 , \42741 );
xor \U$42400 ( \42743 , \41757 , \41759 );
xor \U$42401 ( \42744 , \42743 , \41762 );
and \U$42402 ( \42745 , \42714 , \42744 );
xor \U$42403 ( \42746 , \41757 , \41759 );
xor \U$42404 ( \42747 , \42746 , \41762 );
and \U$42405 ( \42748 , \42718 , \42747 );
and \U$42406 ( \42749 , \42714 , \42718 );
or \U$42407 ( \42750 , \42745 , \42748 , \42749 );
xor \U$42408 ( \42751 , \42742 , \42750 );
and \U$42409 ( \42752 , \42733 , \42751 );
xor \U$42410 ( \42753 , \42047 , \42049 );
xor \U$42411 ( \42754 , \42753 , \42052 );
xor \U$42412 ( \42755 , \42701 , \42703 );
and \U$42413 ( \42756 , \42755 , \42706 );
and \U$42414 ( \42757 , \42701 , \42703 );
or \U$42415 ( \42758 , \42756 , \42757 );
xor \U$42416 ( \42759 , \41405 , \41407 );
xor \U$42417 ( \42760 , \42759 , \41410 );
xor \U$42418 ( \42761 , \42024 , \42031 );
xor \U$42419 ( \42762 , \42760 , \42761 );
xor \U$42420 ( \42763 , \42758 , \42762 );
xor \U$42421 ( \42764 , \42754 , \42763 );
xor \U$42422 ( \42765 , \42737 , \42741 );
xor \U$42423 ( \42766 , \42765 , \42750 );
and \U$42424 ( \42767 , \42764 , \42766 );
and \U$42425 ( \42768 , \42733 , \42764 );
or \U$42426 ( \42769 , \42752 , \42767 , \42768 );
xor \U$42427 ( \42770 , \42728 , \42769 );
xor \U$42428 ( \42771 , \41781 , \42019 );
xor \U$42429 ( \42772 , \42771 , \42036 );
xor \U$42430 ( \42773 , \42041 , \42043 );
xor \U$42431 ( \42774 , \41676 , \41678 );
xor \U$42432 ( \42775 , \42774 , \41681 );
xor \U$42433 ( \42776 , \42055 , \42062 );
xor \U$42434 ( \42777 , \42775 , \42776 );
xor \U$42435 ( \42778 , \42773 , \42777 );
xor \U$42436 ( \42779 , \42772 , \42778 );
and \U$42437 ( \42780 , \42770 , \42779 );
and \U$42438 ( \42781 , \42728 , \42769 );
or \U$42439 ( \42782 , \42780 , \42781 );
xor \U$42440 ( \42783 , \42039 , \42044 );
xor \U$42441 ( \42784 , \42783 , \42067 );
xor \U$42442 ( \42785 , \42782 , \42784 );
xor \U$42443 ( \42786 , \42737 , \42741 );
and \U$42444 ( \42787 , \42786 , \42750 );
and \U$42445 ( \42788 , \42737 , \42741 );
or \U$42446 ( \42789 , \42787 , \42788 );
and \U$42447 ( \42790 , \42730 , \42732 );
xor \U$42448 ( \42791 , \42789 , \42790 );
xor \U$42449 ( \42792 , \42047 , \42049 );
xor \U$42450 ( \42793 , \42792 , \42052 );
and \U$42451 ( \42794 , \42758 , \42793 );
xor \U$42452 ( \42795 , \42047 , \42049 );
xor \U$42453 ( \42796 , \42795 , \42052 );
and \U$42454 ( \42797 , \42762 , \42796 );
and \U$42455 ( \42798 , \42758 , \42762 );
or \U$42456 ( \42799 , \42794 , \42797 , \42798 );
and \U$42457 ( \42800 , \42791 , \42799 );
and \U$42458 ( \42801 , \42789 , \42790 );
or \U$42459 ( \42802 , \42800 , \42801 );
xor \U$42460 ( \42803 , \41781 , \42019 );
xor \U$42461 ( \42804 , \42803 , \42036 );
and \U$42462 ( \42805 , \42773 , \42804 );
xor \U$42463 ( \42806 , \41781 , \42019 );
xor \U$42464 ( \42807 , \42806 , \42036 );
and \U$42465 ( \42808 , \42777 , \42807 );
and \U$42466 ( \42809 , \42773 , \42777 );
or \U$42467 ( \42810 , \42805 , \42808 , \42809 );
xor \U$42468 ( \42811 , \42802 , \42810 );
xor \U$42469 ( \42812 , \41416 , \41648 );
xor \U$42470 ( \42813 , \42812 , \41665 );
xor \U$42471 ( \42814 , \42071 , \42078 );
xor \U$42472 ( \42815 , \42813 , \42814 );
xor \U$42473 ( \42816 , \42811 , \42815 );
and \U$42474 ( \42817 , \42785 , \42816 );
and \U$42475 ( \42818 , \42782 , \42784 );
or \U$42476 ( \42819 , \42817 , \42818 );
xor \U$42477 ( \42820 , \42802 , \42810 );
and \U$42478 ( \42821 , \42820 , \42815 );
and \U$42479 ( \42822 , \42802 , \42810 );
or \U$42480 ( \42823 , \42821 , \42822 );
xor \U$42481 ( \42824 , \41668 , \41673 );
xor \U$42482 ( \42825 , \42824 , \41696 );
xor \U$42483 ( \42826 , \42823 , \42825 );
xor \U$42484 ( \42827 , \42070 , \42083 );
xor \U$42485 ( \42828 , \42827 , \42088 );
xor \U$42486 ( \42829 , \42826 , \42828 );
and \U$42487 ( \42830 , \42819 , \42829 );
not \U$42488 ( \42831 , \42830 );
xor \U$42489 ( \42832 , \42823 , \42825 );
and \U$42490 ( \42833 , \42832 , \42828 );
and \U$42491 ( \42834 , \42823 , \42825 );
or \U$42492 ( \42835 , \42833 , \42834 );
xor \U$42493 ( \42836 , \41740 , \41742 );
xor \U$42494 ( \42837 , \42836 , \42091 );
xor \U$42495 ( \42838 , \42835 , \42837 );
not \U$42496 ( \42839 , \42838 );
or \U$42497 ( \42840 , \42831 , \42839 );
xor \U$42498 ( \42841 , \42592 , \42688 );
xor \U$42499 ( \42842 , \42841 , \42725 );
xor \U$42500 ( \42843 , \42665 , \42687 );
xor \U$42501 ( \42844 , \42315 , \42558 );
xor \U$42502 ( \42845 , \42844 , \42589 );
and \U$42503 ( \42846 , \42843 , \42845 );
xor \U$42504 ( \42847 , \42701 , \42703 );
xor \U$42505 ( \42848 , \42847 , \42706 );
xor \U$42506 ( \42849 , \42699 , \42720 );
xor \U$42507 ( \42850 , \42848 , \42849 );
xor \U$42508 ( \42851 , \42315 , \42558 );
xor \U$42509 ( \42852 , \42851 , \42589 );
and \U$42510 ( \42853 , \42850 , \42852 );
and \U$42511 ( \42854 , \42843 , \42850 );
or \U$42512 ( \42855 , \42846 , \42853 , \42854 );
xor \U$42513 ( \42856 , \42378 , \42385 );
xor \U$42514 ( \42857 , \42856 , \42393 );
xor \U$42515 ( \42858 , \42533 , \42540 );
xor \U$42516 ( \42859 , \42858 , \42549 );
and \U$42517 ( \42860 , \42857 , \42859 );
xor \U$42518 ( \42861 , \42506 , \42513 );
xor \U$42519 ( \42862 , \42861 , \42522 );
xor \U$42520 ( \42863 , \42533 , \42540 );
xor \U$42521 ( \42864 , \42863 , \42549 );
and \U$42522 ( \42865 , \42862 , \42864 );
and \U$42523 ( \42866 , \42857 , \42862 );
or \U$42524 ( \42867 , \42860 , \42865 , \42866 );
not \U$42525 ( \42868 , RI986fd18_70);
nor \U$42526 ( \42869 , \42868 , \407 );
xor \U$42527 ( \42870 , \42349 , \42357 );
xor \U$42528 ( \42871 , \42870 , \42366 );
and \U$42529 ( \42872 , \42869 , \42871 );
xor \U$42530 ( \42873 , \42323 , \42331 );
xor \U$42531 ( \42874 , \42873 , \42339 );
xor \U$42532 ( \42875 , \42349 , \42357 );
xor \U$42533 ( \42876 , \42875 , \42366 );
and \U$42534 ( \42877 , \42874 , \42876 );
and \U$42535 ( \42878 , \42869 , \42874 );
or \U$42536 ( \42879 , \42872 , \42877 , \42878 );
xor \U$42537 ( \42880 , \42867 , \42879 );
xor \U$42538 ( \42881 , \42406 , \42413 );
xor \U$42539 ( \42882 , \42881 , \42421 );
xor \U$42540 ( \42883 , \42479 , \42486 );
xor \U$42541 ( \42884 , \42883 , \42495 );
xor \U$42542 ( \42885 , \42882 , \42884 );
xor \U$42543 ( \42886 , \42450 , \42457 );
xor \U$42544 ( \42887 , \42886 , \42465 );
and \U$42545 ( \42888 , \42885 , \42887 );
and \U$42546 ( \42889 , \42882 , \42884 );
or \U$42547 ( \42890 , \42888 , \42889 );
and \U$42548 ( \42891 , \42880 , \42890 );
and \U$42549 ( \42892 , \42867 , \42879 );
or \U$42550 ( \42893 , \42891 , \42892 );
and \U$42551 ( \42894 , \8486 , RI986f688_56);
and \U$42552 ( \42895 , RI986e008_8, \8484 );
nor \U$42553 ( \42896 , \42894 , \42895 );
and \U$42554 ( \42897 , \42896 , \8050 );
not \U$42555 ( \42898 , \42896 );
and \U$42556 ( \42899 , \42898 , \8051 );
nor \U$42557 ( \42900 , \42897 , \42899 );
and \U$42558 ( \42901 , \7729 , RI986f3b8_50);
and \U$42559 ( \42902 , RI986f598_54, \7727 );
nor \U$42560 ( \42903 , \42901 , \42902 );
and \U$42561 ( \42904 , \42903 , \7480 );
not \U$42562 ( \42905 , \42903 );
and \U$42563 ( \42906 , \42905 , \7733 );
nor \U$42564 ( \42907 , \42904 , \42906 );
xor \U$42565 ( \42908 , \42900 , \42907 );
and \U$42566 ( \42909 , \9237 , RI986df18_6);
and \U$42567 ( \42910 , RI986de28_4, \9235 );
nor \U$42568 ( \42911 , \42909 , \42910 );
and \U$42569 ( \42912 , \42911 , \9241 );
not \U$42570 ( \42913 , \42911 );
and \U$42571 ( \42914 , \42913 , \8836 );
nor \U$42572 ( \42915 , \42912 , \42914 );
and \U$42573 ( \42916 , \42908 , \42915 );
and \U$42574 ( \42917 , \42900 , \42907 );
or \U$42575 ( \42918 , \42916 , \42917 );
and \U$42576 ( \42919 , \9505 , RI986dd38_2);
and \U$42577 ( \42920 , RI986e1e8_12, \9503 );
nor \U$42578 ( \42921 , \42919 , \42920 );
and \U$42579 ( \42922 , \42921 , \9510 );
not \U$42580 ( \42923 , \42921 );
and \U$42581 ( \42924 , \42923 , \9513 );
nor \U$42582 ( \42925 , \42922 , \42924 );
nand \U$42583 ( \42926 , RI986e3c8_16, \11696 );
and \U$42584 ( \42927 , \42926 , \10965 );
not \U$42585 ( \42928 , \42926 );
and \U$42586 ( \42929 , \42928 , \11702 );
nor \U$42587 ( \42930 , \42927 , \42929 );
xor \U$42588 ( \42931 , \42925 , \42930 );
and \U$42589 ( \42932 , \10424 , RI986e0f8_10);
and \U$42590 ( \42933 , RI986e2d8_14, \10422 );
nor \U$42591 ( \42934 , \42932 , \42933 );
and \U$42592 ( \42935 , \42934 , \9840 );
not \U$42593 ( \42936 , \42934 );
and \U$42594 ( \42937 , \42936 , \10428 );
nor \U$42595 ( \42938 , \42935 , \42937 );
and \U$42596 ( \42939 , \42931 , \42938 );
and \U$42597 ( \42940 , \42925 , \42930 );
or \U$42598 ( \42941 , \42939 , \42940 );
xor \U$42599 ( \42942 , \42918 , \42941 );
and \U$42600 ( \42943 , \5881 , RI986e698_22);
and \U$42601 ( \42944 , RI986f868_60, \5879 );
nor \U$42602 ( \42945 , \42943 , \42944 );
and \U$42603 ( \42946 , \42945 , \5594 );
not \U$42604 ( \42947 , \42945 );
and \U$42605 ( \42948 , \42947 , \5885 );
nor \U$42606 ( \42949 , \42946 , \42948 );
and \U$42607 ( \42950 , \6453 , RI986f778_58);
and \U$42608 ( \42951 , RI986fa48_64, \6451 );
nor \U$42609 ( \42952 , \42950 , \42951 );
and \U$42610 ( \42953 , \42952 , \6190 );
not \U$42611 ( \42954 , \42952 );
and \U$42612 ( \42955 , \42954 , \6705 );
nor \U$42613 ( \42956 , \42953 , \42955 );
xor \U$42614 ( \42957 , \42949 , \42956 );
and \U$42615 ( \42958 , \7079 , RI986f958_62);
and \U$42616 ( \42959 , RI986f4a8_52, \7077 );
nor \U$42617 ( \42960 , \42958 , \42959 );
and \U$42618 ( \42961 , \42960 , \6710 );
not \U$42619 ( \42962 , \42960 );
and \U$42620 ( \42963 , \42962 , \6709 );
nor \U$42621 ( \42964 , \42961 , \42963 );
and \U$42622 ( \42965 , \42957 , \42964 );
and \U$42623 ( \42966 , \42949 , \42956 );
or \U$42624 ( \42967 , \42965 , \42966 );
and \U$42625 ( \42968 , \42942 , \42967 );
and \U$42626 ( \42969 , \42918 , \42941 );
or \U$42627 ( \42970 , \42968 , \42969 );
and \U$42628 ( \42971 , \438 , RI9870c18_102);
and \U$42629 ( \42972 , RI98710c8_112, \436 );
nor \U$42630 ( \42973 , \42971 , \42972 );
and \U$42631 ( \42974 , \42973 , \444 );
not \U$42632 ( \42975 , \42973 );
and \U$42633 ( \42976 , \42975 , \443 );
nor \U$42634 ( \42977 , \42974 , \42976 );
not \U$42635 ( \42978 , \454 );
and \U$42636 ( \42979 , \465 , RI9870a38_98);
and \U$42637 ( \42980 , RI9870ee8_108, \463 );
nor \U$42638 ( \42981 , \42979 , \42980 );
not \U$42639 ( \42982 , \42981 );
or \U$42640 ( \42983 , \42978 , \42982 );
or \U$42641 ( \42984 , \42981 , \454 );
nand \U$42642 ( \42985 , \42983 , \42984 );
xor \U$42643 ( \42986 , \42977 , \42985 );
not \U$42644 ( \42987 , \367 );
and \U$42645 ( \42988 , \376 , RI9870b28_100);
and \U$42646 ( \42989 , RI9870df8_106, \374 );
nor \U$42647 ( \42990 , \42988 , \42989 );
not \U$42648 ( \42991 , \42990 );
or \U$42649 ( \42992 , \42987 , \42991 );
or \U$42650 ( \42993 , \42990 , \365 );
nand \U$42651 ( \42994 , \42992 , \42993 );
and \U$42652 ( \42995 , \42986 , \42994 );
and \U$42653 ( \42996 , \42977 , \42985 );
or \U$42654 ( \42997 , \42995 , \42996 );
and \U$42655 ( \42998 , \354 , RI986fef8_74);
and \U$42656 ( \42999 , RI98700d8_78, \352 );
nor \U$42657 ( \43000 , \42998 , \42999 );
not \U$42658 ( \43001 , \43000 );
not \U$42659 ( \43002 , \361 );
and \U$42660 ( \43003 , \43001 , \43002 );
and \U$42661 ( \43004 , \43000 , \345 );
nor \U$42662 ( \43005 , \43003 , \43004 );
and \U$42663 ( \43006 , \416 , RI986fd18_70);
and \U$42664 ( \43007 , RI986ffe8_76, \414 );
nor \U$42665 ( \43008 , \43006 , \43007 );
and \U$42666 ( \43009 , \43008 , \421 );
not \U$42667 ( \43010 , \43008 );
and \U$42668 ( \43011 , \43010 , \422 );
nor \U$42669 ( \43012 , \43009 , \43011 );
or \U$42670 ( \43013 , \43005 , \43012 );
not \U$42671 ( \43014 , \43012 );
not \U$42672 ( \43015 , \43005 );
or \U$42673 ( \43016 , \43014 , \43015 );
not \U$42674 ( \43017 , \386 );
and \U$42675 ( \43018 , \395 , RI98701c8_80);
and \U$42676 ( \43019 , RI9870fd8_110, \393 );
nor \U$42677 ( \43020 , \43018 , \43019 );
not \U$42678 ( \43021 , \43020 );
or \U$42679 ( \43022 , \43017 , \43021 );
or \U$42680 ( \43023 , \43020 , \487 );
nand \U$42681 ( \43024 , \43022 , \43023 );
nand \U$42682 ( \43025 , \43016 , \43024 );
nand \U$42683 ( \43026 , \43013 , \43025 );
xor \U$42684 ( \43027 , \42997 , \43026 );
and \U$42685 ( \43028 , \776 , RI9870d08_104);
and \U$42686 ( \43029 , RI98712a8_116, \774 );
nor \U$42687 ( \43030 , \43028 , \43029 );
and \U$42688 ( \43031 , \43030 , \474 );
not \U$42689 ( \43032 , \43030 );
and \U$42690 ( \43033 , \43032 , \451 );
nor \U$42691 ( \43034 , \43031 , \43033 );
not \U$42692 ( \43035 , \1301 );
and \U$42693 ( \43036 , \1293 , RI98711b8_114);
and \U$42694 ( \43037 , RI9871398_118, \1291 );
nor \U$42695 ( \43038 , \43036 , \43037 );
not \U$42696 ( \43039 , \43038 );
or \U$42697 ( \43040 , \43035 , \43039 );
or \U$42698 ( \43041 , \43038 , \1301 );
nand \U$42699 ( \43042 , \43040 , \43041 );
xor \U$42700 ( \43043 , \43034 , \43042 );
and \U$42701 ( \43044 , \1329 , RI9871488_120);
and \U$42702 ( \43045 , RI9871758_126, \1327 );
nor \U$42703 ( \43046 , \43044 , \43045 );
and \U$42704 ( \43047 , \43046 , \1336 );
not \U$42705 ( \43048 , \43046 );
and \U$42706 ( \43049 , \43048 , \1337 );
nor \U$42707 ( \43050 , \43047 , \43049 );
and \U$42708 ( \43051 , \43043 , \43050 );
and \U$42709 ( \43052 , \43034 , \43042 );
or \U$42710 ( \43053 , \43051 , \43052 );
and \U$42711 ( \43054 , \43027 , \43053 );
and \U$42712 ( \43055 , \42997 , \43026 );
or \U$42713 ( \43056 , \43054 , \43055 );
xor \U$42714 ( \43057 , \42970 , \43056 );
not \U$42715 ( \43058 , \4519 );
and \U$42716 ( \43059 , \4710 , RI986f1d8_46);
and \U$42717 ( \43060 , RI986e5a8_20, \4708 );
nor \U$42718 ( \43061 , \43059 , \43060 );
not \U$42719 ( \43062 , \43061 );
or \U$42720 ( \43063 , \43058 , \43062 );
or \U$42721 ( \43064 , \43061 , \4521 );
nand \U$42722 ( \43065 , \43063 , \43064 );
and \U$42723 ( \43066 , \4203 , RI986eff8_42);
and \U$42724 ( \43067 , RI986f2c8_48, \4201 );
nor \U$42725 ( \43068 , \43066 , \43067 );
and \U$42726 ( \43069 , \43068 , \4207 );
not \U$42727 ( \43070 , \43068 );
and \U$42728 ( \43071 , \43070 , \3923 );
nor \U$42729 ( \43072 , \43069 , \43071 );
xor \U$42730 ( \43073 , \43065 , \43072 );
and \U$42731 ( \43074 , \5318 , RI986e4b8_18);
and \U$42732 ( \43075 , RI986e788_24, \5316 );
nor \U$42733 ( \43076 , \43074 , \43075 );
and \U$42734 ( \43077 , \43076 , \5052 );
not \U$42735 ( \43078 , \43076 );
and \U$42736 ( \43079 , \43078 , \5322 );
nor \U$42737 ( \43080 , \43077 , \43079 );
and \U$42738 ( \43081 , \43073 , \43080 );
and \U$42739 ( \43082 , \43065 , \43072 );
or \U$42740 ( \43083 , \43081 , \43082 );
and \U$42741 ( \43084 , \2274 , RI986ea58_30);
and \U$42742 ( \43085 , RI986e968_28, \2272 );
nor \U$42743 ( \43086 , \43084 , \43085 );
and \U$42744 ( \43087 , \43086 , \2030 );
not \U$42745 ( \43088 , \43086 );
and \U$42746 ( \43089 , \43088 , \2031 );
nor \U$42747 ( \43090 , \43087 , \43089 );
and \U$42748 ( \43091 , \1311 , RI9871848_128);
and \U$42749 ( \43092 , RI9871578_122, \1309 );
nor \U$42750 ( \43093 , \43091 , \43092 );
and \U$42751 ( \43094 , \43093 , \1458 );
not \U$42752 ( \43095 , \43093 );
and \U$42753 ( \43096 , \43095 , \1315 );
nor \U$42754 ( \43097 , \43094 , \43096 );
xor \U$42755 ( \43098 , \43090 , \43097 );
not \U$42756 ( \43099 , \1462 );
and \U$42757 ( \43100 , \2042 , RI9871668_124);
and \U$42758 ( \43101 , RI986eb48_32, \2040 );
nor \U$42759 ( \43102 , \43100 , \43101 );
not \U$42760 ( \43103 , \43102 );
or \U$42761 ( \43104 , \43099 , \43103 );
or \U$42762 ( \43105 , \43102 , \1462 );
nand \U$42763 ( \43106 , \43104 , \43105 );
and \U$42764 ( \43107 , \43098 , \43106 );
and \U$42765 ( \43108 , \43090 , \43097 );
or \U$42766 ( \43109 , \43107 , \43108 );
xor \U$42767 ( \43110 , \43083 , \43109 );
not \U$42768 ( \43111 , \2935 );
and \U$42769 ( \43112 , \3254 , RI986ee18_38);
and \U$42770 ( \43113 , RI986ec38_34, \3252 );
nor \U$42771 ( \43114 , \43112 , \43113 );
not \U$42772 ( \43115 , \43114 );
or \U$42773 ( \43116 , \43111 , \43115 );
or \U$42774 ( \43117 , \43114 , \2935 );
nand \U$42775 ( \43118 , \43116 , \43117 );
and \U$42776 ( \43119 , \2464 , RI986e878_26);
and \U$42777 ( \43120 , RI986ef08_40, \2462 );
nor \U$42778 ( \43121 , \43119 , \43120 );
and \U$42779 ( \43122 , \43121 , \2468 );
not \U$42780 ( \43123 , \43121 );
and \U$42781 ( \43124 , \43123 , \2263 );
nor \U$42782 ( \43125 , \43122 , \43124 );
xor \U$42783 ( \43126 , \43118 , \43125 );
not \U$42784 ( \43127 , \3918 );
and \U$42785 ( \43128 , \3683 , RI986ed28_36);
and \U$42786 ( \43129 , RI986f0e8_44, \3681 );
nor \U$42787 ( \43130 , \43128 , \43129 );
not \U$42788 ( \43131 , \43130 );
or \U$42789 ( \43132 , \43127 , \43131 );
or \U$42790 ( \43133 , \43130 , \3918 );
nand \U$42791 ( \43134 , \43132 , \43133 );
and \U$42792 ( \43135 , \43126 , \43134 );
and \U$42793 ( \43136 , \43118 , \43125 );
or \U$42794 ( \43137 , \43135 , \43136 );
and \U$42795 ( \43138 , \43110 , \43137 );
and \U$42796 ( \43139 , \43083 , \43109 );
or \U$42797 ( \43140 , \43138 , \43139 );
and \U$42798 ( \43141 , \43057 , \43140 );
and \U$42799 ( \43142 , \42970 , \43056 );
or \U$42800 ( \43143 , \43141 , \43142 );
xor \U$42801 ( \43144 , \42893 , \43143 );
xor \U$42802 ( \43145 , \42640 , \42645 );
xor \U$42803 ( \43146 , \43145 , \42653 );
xor \U$42804 ( \43147 , \42260 , \42284 );
xor \U$42805 ( \43148 , \43147 , \42309 );
and \U$42806 ( \43149 , \43146 , \43148 );
xor \U$42807 ( \43150 , \42129 , \42136 );
xor \U$42808 ( \43151 , \43150 , \42144 );
xor \U$42809 ( \43152 , \42122 , \42169 );
xor \U$42810 ( \43153 , \43151 , \43152 );
xor \U$42811 ( \43154 , \42260 , \42284 );
xor \U$42812 ( \43155 , \43154 , \42309 );
and \U$42813 ( \43156 , \43153 , \43155 );
and \U$42814 ( \43157 , \43146 , \43153 );
or \U$42815 ( \43158 , \43149 , \43156 , \43157 );
and \U$42816 ( \43159 , \43144 , \43158 );
and \U$42817 ( \43160 , \42893 , \43143 );
or \U$42818 ( \43161 , \43159 , \43160 );
xor \U$42819 ( \43162 , \42399 , \42471 );
xor \U$42820 ( \43163 , \43162 , \42555 );
xor \U$42821 ( \43164 , \42174 , \42235 );
xor \U$42822 ( \43165 , \43164 , \42312 );
and \U$42823 ( \43166 , \43163 , \43165 );
xor \U$42824 ( \43167 , \43161 , \43166 );
or \U$42825 ( \43168 , \42200 , \42234 );
nand \U$42826 ( \43169 , \43168 , \42235 );
xor \U$42827 ( \43170 , \42342 , \42369 );
xor \U$42828 ( \43171 , \43170 , \42396 );
and \U$42829 ( \43172 , \43169 , \43171 );
xor \U$42830 ( \43173 , \42498 , \42525 );
xor \U$42831 ( \43174 , \43173 , \42552 );
xor \U$42832 ( \43175 , \42342 , \42369 );
xor \U$42833 ( \43176 , \43175 , \42396 );
and \U$42834 ( \43177 , \43174 , \43176 );
and \U$42835 ( \43178 , \43169 , \43174 );
or \U$42836 ( \43179 , \43172 , \43177 , \43178 );
xor \U$42837 ( \43180 , \42691 , \42693 );
xor \U$42838 ( \43181 , \43180 , \42696 );
and \U$42839 ( \43182 , \43179 , \43181 );
xor \U$42840 ( \43183 , \42569 , \42571 );
xor \U$42841 ( \43184 , \43183 , \42574 );
xor \U$42842 ( \43185 , \42567 , \42584 );
xor \U$42843 ( \43186 , \43184 , \43185 );
xor \U$42844 ( \43187 , \42691 , \42693 );
xor \U$42845 ( \43188 , \43187 , \42696 );
and \U$42846 ( \43189 , \43186 , \43188 );
and \U$42847 ( \43190 , \43179 , \43186 );
or \U$42848 ( \43191 , \43182 , \43189 , \43190 );
and \U$42849 ( \43192 , \43167 , \43191 );
and \U$42850 ( \43193 , \43161 , \43166 );
or \U$42851 ( \43194 , \43192 , \43193 );
xor \U$42852 ( \43195 , \42855 , \43194 );
xor \U$42853 ( \43196 , \42737 , \42741 );
xor \U$42854 ( \43197 , \43196 , \42750 );
xor \U$42855 ( \43198 , \42733 , \42764 );
xor \U$42856 ( \43199 , \43197 , \43198 );
xor \U$42857 ( \43200 , \43195 , \43199 );
and \U$42858 ( \43201 , \42842 , \43200 );
xor \U$42859 ( \43202 , \43083 , \43109 );
xor \U$42860 ( \43203 , \43202 , \43137 );
xor \U$42861 ( \43204 , \42997 , \43026 );
xor \U$42862 ( \43205 , \43204 , \43053 );
and \U$42863 ( \43206 , \43203 , \43205 );
xor \U$42864 ( \43207 , \42349 , \42357 );
xor \U$42865 ( \43208 , \43207 , \42366 );
xor \U$42866 ( \43209 , \42869 , \42874 );
xor \U$42867 ( \43210 , \43208 , \43209 );
xor \U$42868 ( \43211 , \42997 , \43026 );
xor \U$42869 ( \43212 , \43211 , \43053 );
and \U$42870 ( \43213 , \43210 , \43212 );
and \U$42871 ( \43214 , \43203 , \43210 );
or \U$42872 ( \43215 , \43206 , \43213 , \43214 );
xor \U$42873 ( \43216 , \42424 , \42442 );
xor \U$42874 ( \43217 , \43216 , \42468 );
xor \U$42875 ( \43218 , \43215 , \43217 );
xor \U$42876 ( \43219 , \42342 , \42369 );
xor \U$42877 ( \43220 , \43219 , \42396 );
xor \U$42878 ( \43221 , \43169 , \43174 );
xor \U$42879 ( \43222 , \43220 , \43221 );
and \U$42880 ( \43223 , \43218 , \43222 );
and \U$42881 ( \43224 , \43215 , \43217 );
or \U$42882 ( \43225 , \43223 , \43224 );
xor \U$42883 ( \43226 , \43118 , \43125 );
xor \U$42884 ( \43227 , \43226 , \43134 );
xor \U$42885 ( \43228 , \42949 , \42956 );
xor \U$42886 ( \43229 , \43228 , \42964 );
and \U$42887 ( \43230 , \43227 , \43229 );
xor \U$42888 ( \43231 , \43065 , \43072 );
xor \U$42889 ( \43232 , \43231 , \43080 );
xor \U$42890 ( \43233 , \42949 , \42956 );
xor \U$42891 ( \43234 , \43233 , \42964 );
and \U$42892 ( \43235 , \43232 , \43234 );
and \U$42893 ( \43236 , \43227 , \43232 );
or \U$42894 ( \43237 , \43230 , \43235 , \43236 );
nand \U$42895 ( \43238 , RI986fe08_72, RI9871fc8_144);
not \U$42896 ( \43239 , \43005 );
not \U$42897 ( \43240 , \43024 );
or \U$42898 ( \43241 , \43239 , \43240 );
or \U$42899 ( \43242 , \43005 , \43024 );
nand \U$42900 ( \43243 , \43241 , \43242 );
not \U$42901 ( \43244 , \43243 );
not \U$42902 ( \43245 , \43012 );
and \U$42903 ( \43246 , \43244 , \43245 );
and \U$42904 ( \43247 , \43243 , \43012 );
nor \U$42905 ( \43248 , \43246 , \43247 );
nand \U$42906 ( \43249 , \43238 , \43248 );
xor \U$42907 ( \43250 , \43237 , \43249 );
xor \U$42908 ( \43251 , \43090 , \43097 );
xor \U$42909 ( \43252 , \43251 , \43106 );
xor \U$42910 ( \43253 , \42977 , \42985 );
xor \U$42911 ( \43254 , \43253 , \42994 );
xor \U$42912 ( \43255 , \43252 , \43254 );
xor \U$42913 ( \43256 , \43034 , \43042 );
xor \U$42914 ( \43257 , \43256 , \43050 );
and \U$42915 ( \43258 , \43255 , \43257 );
and \U$42916 ( \43259 , \43252 , \43254 );
or \U$42917 ( \43260 , \43258 , \43259 );
and \U$42918 ( \43261 , \43250 , \43260 );
and \U$42919 ( \43262 , \43237 , \43249 );
or \U$42920 ( \43263 , \43261 , \43262 );
and \U$42921 ( \43264 , \6453 , RI986f868_60);
and \U$42922 ( \43265 , RI986f778_58, \6451 );
nor \U$42923 ( \43266 , \43264 , \43265 );
and \U$42924 ( \43267 , \43266 , \6190 );
not \U$42925 ( \43268 , \43266 );
and \U$42926 ( \43269 , \43268 , \6180 );
nor \U$42927 ( \43270 , \43267 , \43269 );
and \U$42928 ( \43271 , \7079 , RI986fa48_64);
and \U$42929 ( \43272 , RI986f958_62, \7077 );
nor \U$42930 ( \43273 , \43271 , \43272 );
and \U$42931 ( \43274 , \43273 , \6710 );
not \U$42932 ( \43275 , \43273 );
and \U$42933 ( \43276 , \43275 , \6709 );
nor \U$42934 ( \43277 , \43274 , \43276 );
xor \U$42935 ( \43278 , \43270 , \43277 );
and \U$42936 ( \43279 , \7729 , RI986f4a8_52);
and \U$42937 ( \43280 , RI986f3b8_50, \7727 );
nor \U$42938 ( \43281 , \43279 , \43280 );
and \U$42939 ( \43282 , \43281 , \7480 );
not \U$42940 ( \43283 , \43281 );
and \U$42941 ( \43284 , \43283 , \7733 );
nor \U$42942 ( \43285 , \43282 , \43284 );
and \U$42943 ( \43286 , \43278 , \43285 );
and \U$42944 ( \43287 , \43270 , \43277 );
or \U$42945 ( \43288 , \43286 , \43287 );
and \U$42946 ( \43289 , \10424 , RI986e1e8_12);
and \U$42947 ( \43290 , RI986e0f8_10, \10422 );
nor \U$42948 ( \43291 , \43289 , \43290 );
and \U$42949 ( \43292 , \43291 , \9840 );
not \U$42950 ( \43293 , \43291 );
and \U$42951 ( \43294 , \43293 , \10428 );
nor \U$42952 ( \43295 , \43292 , \43294 );
xor \U$42953 ( \43296 , \43295 , \11687 );
and \U$42954 ( \43297 , \11696 , RI986e2d8_14);
and \U$42955 ( \43298 , RI986e3c8_16, \11694 );
nor \U$42956 ( \43299 , \43297 , \43298 );
and \U$42957 ( \43300 , \43299 , \10965 );
not \U$42958 ( \43301 , \43299 );
and \U$42959 ( \43302 , \43301 , \11702 );
nor \U$42960 ( \43303 , \43300 , \43302 );
and \U$42961 ( \43304 , \43296 , \43303 );
and \U$42962 ( \43305 , \43295 , \11687 );
or \U$42963 ( \43306 , \43304 , \43305 );
xor \U$42964 ( \43307 , \43288 , \43306 );
and \U$42965 ( \43308 , \8486 , RI986f598_54);
and \U$42966 ( \43309 , RI986f688_56, \8484 );
nor \U$42967 ( \43310 , \43308 , \43309 );
and \U$42968 ( \43311 , \43310 , \8050 );
not \U$42969 ( \43312 , \43310 );
and \U$42970 ( \43313 , \43312 , \8051 );
nor \U$42971 ( \43314 , \43311 , \43313 );
and \U$42972 ( \43315 , \9237 , RI986e008_8);
and \U$42973 ( \43316 , RI986df18_6, \9235 );
nor \U$42974 ( \43317 , \43315 , \43316 );
and \U$42975 ( \43318 , \43317 , \9241 );
not \U$42976 ( \43319 , \43317 );
and \U$42977 ( \43320 , \43319 , \8836 );
nor \U$42978 ( \43321 , \43318 , \43320 );
xor \U$42979 ( \43322 , \43314 , \43321 );
and \U$42980 ( \43323 , \9505 , RI986de28_4);
and \U$42981 ( \43324 , RI986dd38_2, \9503 );
nor \U$42982 ( \43325 , \43323 , \43324 );
and \U$42983 ( \43326 , \43325 , \9510 );
not \U$42984 ( \43327 , \43325 );
and \U$42985 ( \43328 , \43327 , \9513 );
nor \U$42986 ( \43329 , \43326 , \43328 );
and \U$42987 ( \43330 , \43322 , \43329 );
and \U$42988 ( \43331 , \43314 , \43321 );
or \U$42989 ( \43332 , \43330 , \43331 );
and \U$42990 ( \43333 , \43307 , \43332 );
and \U$42991 ( \43334 , \43288 , \43306 );
or \U$42992 ( \43335 , \43333 , \43334 );
not \U$42993 ( \43336 , \456 );
and \U$42994 ( \43337 , \465 , RI9870df8_106);
and \U$42995 ( \43338 , RI9870a38_98, \463 );
nor \U$42996 ( \43339 , \43337 , \43338 );
not \U$42997 ( \43340 , \43339 );
or \U$42998 ( \43341 , \43336 , \43340 );
or \U$42999 ( \43342 , \43339 , \456 );
nand \U$43000 ( \43343 , \43341 , \43342 );
and \U$43001 ( \43344 , \776 , RI98710c8_112);
and \U$43002 ( \43345 , RI9870d08_104, \774 );
nor \U$43003 ( \43346 , \43344 , \43345 );
and \U$43004 ( \43347 , \43346 , \474 );
not \U$43005 ( \43348 , \43346 );
and \U$43006 ( \43349 , \43348 , \451 );
nor \U$43007 ( \43350 , \43347 , \43349 );
xor \U$43008 ( \43351 , \43343 , \43350 );
and \U$43009 ( \43352 , \438 , RI9870ee8_108);
and \U$43010 ( \43353 , RI9870c18_102, \436 );
nor \U$43011 ( \43354 , \43352 , \43353 );
and \U$43012 ( \43355 , \43354 , \444 );
not \U$43013 ( \43356 , \43354 );
and \U$43014 ( \43357 , \43356 , \443 );
nor \U$43015 ( \43358 , \43355 , \43357 );
and \U$43016 ( \43359 , \43351 , \43358 );
and \U$43017 ( \43360 , \43343 , \43350 );
or \U$43018 ( \43361 , \43359 , \43360 );
not \U$43019 ( \43362 , \365 );
and \U$43020 ( \43363 , \376 , RI9870fd8_110);
and \U$43021 ( \43364 , RI9870b28_100, \374 );
nor \U$43022 ( \43365 , \43363 , \43364 );
not \U$43023 ( \43366 , \43365 );
or \U$43024 ( \43367 , \43362 , \43366 );
or \U$43025 ( \43368 , \43365 , \367 );
nand \U$43026 ( \43369 , \43367 , \43368 );
not \U$43027 ( \43370 , \386 );
and \U$43028 ( \43371 , \395 , RI98700d8_78);
and \U$43029 ( \43372 , RI98701c8_80, \393 );
nor \U$43030 ( \43373 , \43371 , \43372 );
not \U$43031 ( \43374 , \43373 );
or \U$43032 ( \43375 , \43370 , \43374 );
or \U$43033 ( \43376 , \43373 , \386 );
nand \U$43034 ( \43377 , \43375 , \43376 );
xor \U$43035 ( \43378 , \43369 , \43377 );
not \U$43036 ( \43379 , \361 );
and \U$43037 ( \43380 , \354 , RI986ffe8_76);
and \U$43038 ( \43381 , RI986fef8_74, \352 );
nor \U$43039 ( \43382 , \43380 , \43381 );
not \U$43040 ( \43383 , \43382 );
or \U$43041 ( \43384 , \43379 , \43383 );
or \U$43042 ( \43385 , \43382 , \345 );
nand \U$43043 ( \43386 , \43384 , \43385 );
and \U$43044 ( \43387 , \43378 , \43386 );
and \U$43045 ( \43388 , \43369 , \43377 );
or \U$43046 ( \43389 , \43387 , \43388 );
xor \U$43047 ( \43390 , \43361 , \43389 );
and \U$43048 ( \43391 , \1311 , RI9871758_126);
and \U$43049 ( \43392 , RI9871848_128, \1309 );
nor \U$43050 ( \43393 , \43391 , \43392 );
and \U$43051 ( \43394 , \43393 , \1458 );
not \U$43052 ( \43395 , \43393 );
and \U$43053 ( \43396 , \43395 , \1318 );
nor \U$43054 ( \43397 , \43394 , \43396 );
not \U$43055 ( \43398 , \1301 );
and \U$43056 ( \43399 , \1293 , RI98712a8_116);
and \U$43057 ( \43400 , RI98711b8_114, \1291 );
nor \U$43058 ( \43401 , \43399 , \43400 );
not \U$43059 ( \43402 , \43401 );
or \U$43060 ( \43403 , \43398 , \43402 );
or \U$43061 ( \43404 , \43401 , \1128 );
nand \U$43062 ( \43405 , \43403 , \43404 );
xor \U$43063 ( \43406 , \43397 , \43405 );
and \U$43064 ( \43407 , \1329 , RI9871398_118);
and \U$43065 ( \43408 , RI9871488_120, \1327 );
nor \U$43066 ( \43409 , \43407 , \43408 );
and \U$43067 ( \43410 , \43409 , \1336 );
not \U$43068 ( \43411 , \43409 );
and \U$43069 ( \43412 , \43411 , \1337 );
nor \U$43070 ( \43413 , \43410 , \43412 );
and \U$43071 ( \43414 , \43406 , \43413 );
and \U$43072 ( \43415 , \43397 , \43405 );
or \U$43073 ( \43416 , \43414 , \43415 );
and \U$43074 ( \43417 , \43390 , \43416 );
and \U$43075 ( \43418 , \43361 , \43389 );
or \U$43076 ( \43419 , \43417 , \43418 );
xor \U$43077 ( \43420 , \43335 , \43419 );
not \U$43078 ( \43421 , \4521 );
and \U$43079 ( \43422 , \4710 , RI986f2c8_48);
and \U$43080 ( \43423 , RI986f1d8_46, \4708 );
nor \U$43081 ( \43424 , \43422 , \43423 );
not \U$43082 ( \43425 , \43424 );
or \U$43083 ( \43426 , \43421 , \43425 );
or \U$43084 ( \43427 , \43424 , \4519 );
nand \U$43085 ( \43428 , \43426 , \43427 );
and \U$43086 ( \43429 , \5318 , RI986e5a8_20);
and \U$43087 ( \43430 , RI986e4b8_18, \5316 );
nor \U$43088 ( \43431 , \43429 , \43430 );
and \U$43089 ( \43432 , \43431 , \5052 );
not \U$43090 ( \43433 , \43431 );
and \U$43091 ( \43434 , \43433 , \5322 );
nor \U$43092 ( \43435 , \43432 , \43434 );
xor \U$43093 ( \43436 , \43428 , \43435 );
and \U$43094 ( \43437 , \5881 , RI986e788_24);
and \U$43095 ( \43438 , RI986e698_22, \5879 );
nor \U$43096 ( \43439 , \43437 , \43438 );
and \U$43097 ( \43440 , \43439 , \5594 );
not \U$43098 ( \43441 , \43439 );
and \U$43099 ( \43442 , \43441 , \5885 );
nor \U$43100 ( \43443 , \43440 , \43442 );
and \U$43101 ( \43444 , \43436 , \43443 );
and \U$43102 ( \43445 , \43428 , \43435 );
or \U$43103 ( \43446 , \43444 , \43445 );
not \U$43104 ( \43447 , \2034 );
and \U$43105 ( \43448 , \2042 , RI9871578_122);
and \U$43106 ( \43449 , RI9871668_124, \2040 );
nor \U$43107 ( \43450 , \43448 , \43449 );
not \U$43108 ( \43451 , \43450 );
or \U$43109 ( \43452 , \43447 , \43451 );
or \U$43110 ( \43453 , \43450 , \2034 );
nand \U$43111 ( \43454 , \43452 , \43453 );
and \U$43112 ( \43455 , \2274 , RI986eb48_32);
and \U$43113 ( \43456 , RI986ea58_30, \2272 );
nor \U$43114 ( \43457 , \43455 , \43456 );
and \U$43115 ( \43458 , \43457 , \2030 );
not \U$43116 ( \43459 , \43457 );
and \U$43117 ( \43460 , \43459 , \2031 );
nor \U$43118 ( \43461 , \43458 , \43460 );
xor \U$43119 ( \43462 , \43454 , \43461 );
and \U$43120 ( \43463 , \2464 , RI986e968_28);
and \U$43121 ( \43464 , RI986e878_26, \2462 );
nor \U$43122 ( \43465 , \43463 , \43464 );
and \U$43123 ( \43466 , \43465 , \2468 );
not \U$43124 ( \43467 , \43465 );
and \U$43125 ( \43468 , \43467 , \2263 );
nor \U$43126 ( \43469 , \43466 , \43468 );
and \U$43127 ( \43470 , \43462 , \43469 );
and \U$43128 ( \43471 , \43454 , \43461 );
or \U$43129 ( \43472 , \43470 , \43471 );
xor \U$43130 ( \43473 , \43446 , \43472 );
not \U$43131 ( \43474 , \3406 );
and \U$43132 ( \43475 , \3254 , RI986ef08_40);
and \U$43133 ( \43476 , RI986ee18_38, \3252 );
nor \U$43134 ( \43477 , \43475 , \43476 );
not \U$43135 ( \43478 , \43477 );
or \U$43136 ( \43479 , \43474 , \43478 );
or \U$43137 ( \43480 , \43477 , \3406 );
nand \U$43138 ( \43481 , \43479 , \43480 );
not \U$43139 ( \43482 , \3918 );
and \U$43140 ( \43483 , \3683 , RI986ec38_34);
and \U$43141 ( \43484 , RI986ed28_36, \3681 );
nor \U$43142 ( \43485 , \43483 , \43484 );
not \U$43143 ( \43486 , \43485 );
or \U$43144 ( \43487 , \43482 , \43486 );
or \U$43145 ( \43488 , \43485 , \3918 );
nand \U$43146 ( \43489 , \43487 , \43488 );
xor \U$43147 ( \43490 , \43481 , \43489 );
and \U$43148 ( \43491 , \4203 , RI986f0e8_44);
and \U$43149 ( \43492 , RI986eff8_42, \4201 );
nor \U$43150 ( \43493 , \43491 , \43492 );
and \U$43151 ( \43494 , \43493 , \4207 );
not \U$43152 ( \43495 , \43493 );
and \U$43153 ( \43496 , \43495 , \3923 );
nor \U$43154 ( \43497 , \43494 , \43496 );
and \U$43155 ( \43498 , \43490 , \43497 );
and \U$43156 ( \43499 , \43481 , \43489 );
or \U$43157 ( \43500 , \43498 , \43499 );
and \U$43158 ( \43501 , \43473 , \43500 );
and \U$43159 ( \43502 , \43446 , \43472 );
or \U$43160 ( \43503 , \43501 , \43502 );
and \U$43161 ( \43504 , \43420 , \43503 );
and \U$43162 ( \43505 , \43335 , \43419 );
or \U$43163 ( \43506 , \43504 , \43505 );
xor \U$43164 ( \43507 , \43263 , \43506 );
xor \U$43165 ( \43508 , \42431 , \10965 );
xor \U$43166 ( \43509 , \43508 , \42439 );
xor \U$43167 ( \43510 , \42882 , \42884 );
xor \U$43168 ( \43511 , \43510 , \42887 );
and \U$43169 ( \43512 , \43509 , \43511 );
xor \U$43170 ( \43513 , \42533 , \42540 );
xor \U$43171 ( \43514 , \43513 , \42549 );
xor \U$43172 ( \43515 , \42857 , \42862 );
xor \U$43173 ( \43516 , \43514 , \43515 );
xor \U$43174 ( \43517 , \42882 , \42884 );
xor \U$43175 ( \43518 , \43517 , \42887 );
and \U$43176 ( \43519 , \43516 , \43518 );
and \U$43177 ( \43520 , \43509 , \43516 );
or \U$43178 ( \43521 , \43512 , \43519 , \43520 );
and \U$43179 ( \43522 , \43507 , \43521 );
and \U$43180 ( \43523 , \43263 , \43506 );
or \U$43181 ( \43524 , \43522 , \43523 );
xor \U$43182 ( \43525 , \43225 , \43524 );
xor \U$43183 ( \43526 , \42970 , \43056 );
xor \U$43184 ( \43527 , \43526 , \43140 );
xor \U$43185 ( \43528 , \42867 , \42879 );
xor \U$43186 ( \43529 , \43528 , \42890 );
and \U$43187 ( \43530 , \43527 , \43529 );
xor \U$43188 ( \43531 , \42260 , \42284 );
xor \U$43189 ( \43532 , \43531 , \42309 );
xor \U$43190 ( \43533 , \43146 , \43153 );
xor \U$43191 ( \43534 , \43532 , \43533 );
xor \U$43192 ( \43535 , \42867 , \42879 );
xor \U$43193 ( \43536 , \43535 , \42890 );
and \U$43194 ( \43537 , \43534 , \43536 );
and \U$43195 ( \43538 , \43527 , \43534 );
or \U$43196 ( \43539 , \43530 , \43537 , \43538 );
and \U$43197 ( \43540 , \43525 , \43539 );
and \U$43198 ( \43541 , \43225 , \43524 );
or \U$43199 ( \43542 , \43540 , \43541 );
xor \U$43200 ( \43543 , \43163 , \43165 );
xor \U$43201 ( \43544 , \42893 , \43143 );
xor \U$43202 ( \43545 , \43544 , \43158 );
and \U$43203 ( \43546 , \43543 , \43545 );
xor \U$43204 ( \43547 , \42691 , \42693 );
xor \U$43205 ( \43548 , \43547 , \42696 );
xor \U$43206 ( \43549 , \43179 , \43186 );
xor \U$43207 ( \43550 , \43548 , \43549 );
xor \U$43208 ( \43551 , \42893 , \43143 );
xor \U$43209 ( \43552 , \43551 , \43158 );
and \U$43210 ( \43553 , \43550 , \43552 );
and \U$43211 ( \43554 , \43543 , \43550 );
or \U$43212 ( \43555 , \43546 , \43553 , \43554 );
xor \U$43213 ( \43556 , \43542 , \43555 );
xor \U$43214 ( \43557 , \42315 , \42558 );
xor \U$43215 ( \43558 , \43557 , \42589 );
xor \U$43216 ( \43559 , \42843 , \42850 );
xor \U$43217 ( \43560 , \43558 , \43559 );
and \U$43218 ( \43561 , \43556 , \43560 );
and \U$43219 ( \43562 , \43542 , \43555 );
or \U$43220 ( \43563 , \43561 , \43562 );
xor \U$43221 ( \43564 , \42855 , \43194 );
xor \U$43222 ( \43565 , \43564 , \43199 );
and \U$43223 ( \43566 , \43563 , \43565 );
and \U$43224 ( \43567 , \42842 , \43563 );
or \U$43225 ( \43568 , \43201 , \43566 , \43567 );
xor \U$43226 ( \43569 , \42855 , \43194 );
and \U$43227 ( \43570 , \43569 , \43199 );
and \U$43228 ( \43571 , \42855 , \43194 );
or \U$43229 ( \43572 , \43570 , \43571 );
xor \U$43230 ( \43573 , \42789 , \42790 );
xor \U$43231 ( \43574 , \43573 , \42799 );
xor \U$43232 ( \43575 , \43572 , \43574 );
xor \U$43233 ( \43576 , \42728 , \42769 );
xor \U$43234 ( \43577 , \43576 , \42779 );
xor \U$43235 ( \43578 , \43575 , \43577 );
and \U$43236 ( \43579 , \43568 , \43578 );
not \U$43237 ( \43580 , \43579 );
xor \U$43238 ( \43581 , \43572 , \43574 );
and \U$43239 ( \43582 , \43581 , \43577 );
and \U$43240 ( \43583 , \43572 , \43574 );
or \U$43241 ( \43584 , \43582 , \43583 );
xor \U$43242 ( \43585 , \42782 , \42784 );
xor \U$43243 ( \43586 , \43585 , \42816 );
xor \U$43244 ( \43587 , \43584 , \43586 );
not \U$43245 ( \43588 , \43587 );
or \U$43246 ( \43589 , \43580 , \43588 );
xor \U$43247 ( \43590 , \43263 , \43506 );
xor \U$43248 ( \43591 , \43590 , \43521 );
xor \U$43249 ( \43592 , \43215 , \43217 );
xor \U$43250 ( \43593 , \43592 , \43222 );
and \U$43251 ( \43594 , \43591 , \43593 );
xor \U$43252 ( \43595 , \42867 , \42879 );
xor \U$43253 ( \43596 , \43595 , \42890 );
xor \U$43254 ( \43597 , \43527 , \43534 );
xor \U$43255 ( \43598 , \43596 , \43597 );
xor \U$43256 ( \43599 , \43215 , \43217 );
xor \U$43257 ( \43600 , \43599 , \43222 );
and \U$43258 ( \43601 , \43598 , \43600 );
and \U$43259 ( \43602 , \43591 , \43598 );
or \U$43260 ( \43603 , \43594 , \43601 , \43602 );
xor \U$43261 ( \43604 , \43446 , \43472 );
xor \U$43262 ( \43605 , \43604 , \43500 );
xor \U$43263 ( \43606 , \43361 , \43389 );
xor \U$43264 ( \43607 , \43606 , \43416 );
xor \U$43265 ( \43608 , \43605 , \43607 );
xor \U$43266 ( \43609 , \43288 , \43306 );
xor \U$43267 ( \43610 , \43609 , \43332 );
and \U$43268 ( \43611 , \43608 , \43610 );
and \U$43269 ( \43612 , \43605 , \43607 );
or \U$43270 ( \43613 , \43611 , \43612 );
xor \U$43271 ( \43614 , \42918 , \42941 );
xor \U$43272 ( \43615 , \43614 , \42967 );
xor \U$43273 ( \43616 , \43613 , \43615 );
or \U$43274 ( \43617 , \43248 , \43238 );
nand \U$43275 ( \43618 , \43617 , \43249 );
xor \U$43276 ( \43619 , \43252 , \43254 );
xor \U$43277 ( \43620 , \43619 , \43257 );
and \U$43278 ( \43621 , \43618 , \43620 );
xor \U$43279 ( \43622 , \42949 , \42956 );
xor \U$43280 ( \43623 , \43622 , \42964 );
xor \U$43281 ( \43624 , \43227 , \43232 );
xor \U$43282 ( \43625 , \43623 , \43624 );
xor \U$43283 ( \43626 , \43252 , \43254 );
xor \U$43284 ( \43627 , \43626 , \43257 );
and \U$43285 ( \43628 , \43625 , \43627 );
and \U$43286 ( \43629 , \43618 , \43625 );
or \U$43287 ( \43630 , \43621 , \43628 , \43629 );
and \U$43288 ( \43631 , \43616 , \43630 );
and \U$43289 ( \43632 , \43613 , \43615 );
or \U$43290 ( \43633 , \43631 , \43632 );
not \U$43291 ( \43634 , \454 );
and \U$43292 ( \43635 , \465 , RI9870b28_100);
and \U$43293 ( \43636 , RI9870df8_106, \463 );
nor \U$43294 ( \43637 , \43635 , \43636 );
not \U$43295 ( \43638 , \43637 );
or \U$43296 ( \43639 , \43634 , \43638 );
or \U$43297 ( \43640 , \43637 , \454 );
nand \U$43298 ( \43641 , \43639 , \43640 );
and \U$43299 ( \43642 , \776 , RI9870c18_102);
and \U$43300 ( \43643 , RI98710c8_112, \774 );
nor \U$43301 ( \43644 , \43642 , \43643 );
and \U$43302 ( \43645 , \43644 , \474 );
not \U$43303 ( \43646 , \43644 );
and \U$43304 ( \43647 , \43646 , \451 );
nor \U$43305 ( \43648 , \43645 , \43647 );
xor \U$43306 ( \43649 , \43641 , \43648 );
and \U$43307 ( \43650 , \438 , RI9870a38_98);
and \U$43308 ( \43651 , RI9870ee8_108, \436 );
nor \U$43309 ( \43652 , \43650 , \43651 );
and \U$43310 ( \43653 , \43652 , \444 );
not \U$43311 ( \43654 , \43652 );
and \U$43312 ( \43655 , \43654 , \443 );
nor \U$43313 ( \43656 , \43653 , \43655 );
and \U$43314 ( \43657 , \43649 , \43656 );
and \U$43315 ( \43658 , \43641 , \43648 );
or \U$43316 ( \43659 , \43657 , \43658 );
not \U$43317 ( \43660 , \345 );
and \U$43318 ( \43661 , \354 , RI986fd18_70);
and \U$43319 ( \43662 , RI986ffe8_76, \352 );
nor \U$43320 ( \43663 , \43661 , \43662 );
not \U$43321 ( \43664 , \43663 );
or \U$43322 ( \43665 , \43660 , \43664 );
or \U$43323 ( \43666 , \43663 , \361 );
nand \U$43324 ( \43667 , \43665 , \43666 );
not \U$43325 ( \43668 , \365 );
and \U$43326 ( \43669 , \376 , RI98701c8_80);
and \U$43327 ( \43670 , RI9870fd8_110, \374 );
nor \U$43328 ( \43671 , \43669 , \43670 );
not \U$43329 ( \43672 , \43671 );
or \U$43330 ( \43673 , \43668 , \43672 );
or \U$43331 ( \43674 , \43671 , \367 );
nand \U$43332 ( \43675 , \43673 , \43674 );
xor \U$43333 ( \43676 , \43667 , \43675 );
not \U$43334 ( \43677 , \487 );
and \U$43335 ( \43678 , \395 , RI986fef8_74);
and \U$43336 ( \43679 , RI98700d8_78, \393 );
nor \U$43337 ( \43680 , \43678 , \43679 );
not \U$43338 ( \43681 , \43680 );
or \U$43339 ( \43682 , \43677 , \43681 );
or \U$43340 ( \43683 , \43680 , \487 );
nand \U$43341 ( \43684 , \43682 , \43683 );
and \U$43342 ( \43685 , \43676 , \43684 );
and \U$43343 ( \43686 , \43667 , \43675 );
or \U$43344 ( \43687 , \43685 , \43686 );
xor \U$43345 ( \43688 , \43659 , \43687 );
and \U$43346 ( \43689 , \1311 , RI9871488_120);
and \U$43347 ( \43690 , RI9871758_126, \1309 );
nor \U$43348 ( \43691 , \43689 , \43690 );
and \U$43349 ( \43692 , \43691 , \1458 );
not \U$43350 ( \43693 , \43691 );
and \U$43351 ( \43694 , \43693 , \1318 );
nor \U$43352 ( \43695 , \43692 , \43694 );
not \U$43353 ( \43696 , \1301 );
and \U$43354 ( \43697 , \1293 , RI9870d08_104);
and \U$43355 ( \43698 , RI98712a8_116, \1291 );
nor \U$43356 ( \43699 , \43697 , \43698 );
not \U$43357 ( \43700 , \43699 );
or \U$43358 ( \43701 , \43696 , \43700 );
or \U$43359 ( \43702 , \43699 , \1128 );
nand \U$43360 ( \43703 , \43701 , \43702 );
xor \U$43361 ( \43704 , \43695 , \43703 );
and \U$43362 ( \43705 , \1329 , RI98711b8_114);
and \U$43363 ( \43706 , RI9871398_118, \1327 );
nor \U$43364 ( \43707 , \43705 , \43706 );
and \U$43365 ( \43708 , \43707 , \1336 );
not \U$43366 ( \43709 , \43707 );
and \U$43367 ( \43710 , \43709 , \1337 );
nor \U$43368 ( \43711 , \43708 , \43710 );
and \U$43369 ( \43712 , \43704 , \43711 );
and \U$43370 ( \43713 , \43695 , \43703 );
or \U$43371 ( \43714 , \43712 , \43713 );
and \U$43372 ( \43715 , \43688 , \43714 );
and \U$43373 ( \43716 , \43659 , \43687 );
or \U$43374 ( \43717 , \43715 , \43716 );
and \U$43375 ( \43718 , \8486 , RI986f3b8_50);
and \U$43376 ( \43719 , RI986f598_54, \8484 );
nor \U$43377 ( \43720 , \43718 , \43719 );
and \U$43378 ( \43721 , \43720 , \8050 );
not \U$43379 ( \43722 , \43720 );
and \U$43380 ( \43723 , \43722 , \8051 );
nor \U$43381 ( \43724 , \43721 , \43723 );
and \U$43382 ( \43725 , \9237 , RI986f688_56);
and \U$43383 ( \43726 , RI986e008_8, \9235 );
nor \U$43384 ( \43727 , \43725 , \43726 );
and \U$43385 ( \43728 , \43727 , \9241 );
not \U$43386 ( \43729 , \43727 );
and \U$43387 ( \43730 , \43729 , \8836 );
nor \U$43388 ( \43731 , \43728 , \43730 );
xor \U$43389 ( \43732 , \43724 , \43731 );
and \U$43390 ( \43733 , \9505 , RI986df18_6);
and \U$43391 ( \43734 , RI986de28_4, \9503 );
nor \U$43392 ( \43735 , \43733 , \43734 );
and \U$43393 ( \43736 , \43735 , \9510 );
not \U$43394 ( \43737 , \43735 );
and \U$43395 ( \43738 , \43737 , \9513 );
nor \U$43396 ( \43739 , \43736 , \43738 );
and \U$43397 ( \43740 , \43732 , \43739 );
and \U$43398 ( \43741 , \43724 , \43731 );
or \U$43399 ( \43742 , \43740 , \43741 );
and \U$43400 ( \43743 , \10424 , RI986dd38_2);
and \U$43401 ( \43744 , RI986e1e8_12, \10422 );
nor \U$43402 ( \43745 , \43743 , \43744 );
and \U$43403 ( \43746 , \43745 , \9840 );
not \U$43404 ( \43747 , \43745 );
and \U$43405 ( \43748 , \43747 , \10428 );
nor \U$43406 ( \43749 , \43746 , \43748 );
nand \U$43407 ( \43750 , RI986e3c8_16, \12293 );
and \U$43408 ( \43751 , \43750 , \11687 );
not \U$43409 ( \43752 , \43750 );
and \U$43410 ( \43753 , \43752 , \11686 );
nor \U$43411 ( \43754 , \43751 , \43753 );
xor \U$43412 ( \43755 , \43749 , \43754 );
and \U$43413 ( \43756 , \11696 , RI986e0f8_10);
and \U$43414 ( \43757 , RI986e2d8_14, \11694 );
nor \U$43415 ( \43758 , \43756 , \43757 );
and \U$43416 ( \43759 , \43758 , \10965 );
not \U$43417 ( \43760 , \43758 );
and \U$43418 ( \43761 , \43760 , \11702 );
nor \U$43419 ( \43762 , \43759 , \43761 );
and \U$43420 ( \43763 , \43755 , \43762 );
and \U$43421 ( \43764 , \43749 , \43754 );
or \U$43422 ( \43765 , \43763 , \43764 );
xor \U$43423 ( \43766 , \43742 , \43765 );
and \U$43424 ( \43767 , \6453 , RI986e698_22);
and \U$43425 ( \43768 , RI986f868_60, \6451 );
nor \U$43426 ( \43769 , \43767 , \43768 );
and \U$43427 ( \43770 , \43769 , \6190 );
not \U$43428 ( \43771 , \43769 );
and \U$43429 ( \43772 , \43771 , \6705 );
nor \U$43430 ( \43773 , \43770 , \43772 );
and \U$43431 ( \43774 , \7079 , RI986f778_58);
and \U$43432 ( \43775 , RI986fa48_64, \7077 );
nor \U$43433 ( \43776 , \43774 , \43775 );
and \U$43434 ( \43777 , \43776 , \6710 );
not \U$43435 ( \43778 , \43776 );
and \U$43436 ( \43779 , \43778 , \6709 );
nor \U$43437 ( \43780 , \43777 , \43779 );
xor \U$43438 ( \43781 , \43773 , \43780 );
and \U$43439 ( \43782 , \7729 , RI986f958_62);
and \U$43440 ( \43783 , RI986f4a8_52, \7727 );
nor \U$43441 ( \43784 , \43782 , \43783 );
and \U$43442 ( \43785 , \43784 , \7480 );
not \U$43443 ( \43786 , \43784 );
and \U$43444 ( \43787 , \43786 , \7733 );
nor \U$43445 ( \43788 , \43785 , \43787 );
and \U$43446 ( \43789 , \43781 , \43788 );
and \U$43447 ( \43790 , \43773 , \43780 );
or \U$43448 ( \43791 , \43789 , \43790 );
and \U$43449 ( \43792 , \43766 , \43791 );
and \U$43450 ( \43793 , \43742 , \43765 );
or \U$43451 ( \43794 , \43792 , \43793 );
xor \U$43452 ( \43795 , \43717 , \43794 );
and \U$43453 ( \43796 , \4203 , RI986ed28_36);
and \U$43454 ( \43797 , RI986f0e8_44, \4201 );
nor \U$43455 ( \43798 , \43796 , \43797 );
and \U$43456 ( \43799 , \43798 , \4207 );
not \U$43457 ( \43800 , \43798 );
and \U$43458 ( \43801 , \43800 , \3923 );
nor \U$43459 ( \43802 , \43799 , \43801 );
not \U$43460 ( \43803 , \2935 );
and \U$43461 ( \43804 , \3254 , RI986e878_26);
and \U$43462 ( \43805 , RI986ef08_40, \3252 );
nor \U$43463 ( \43806 , \43804 , \43805 );
not \U$43464 ( \43807 , \43806 );
or \U$43465 ( \43808 , \43803 , \43807 );
or \U$43466 ( \43809 , \43806 , \2935 );
nand \U$43467 ( \43810 , \43808 , \43809 );
xor \U$43468 ( \43811 , \43802 , \43810 );
not \U$43469 ( \43812 , \3918 );
and \U$43470 ( \43813 , \3683 , RI986ee18_38);
and \U$43471 ( \43814 , RI986ec38_34, \3681 );
nor \U$43472 ( \43815 , \43813 , \43814 );
not \U$43473 ( \43816 , \43815 );
or \U$43474 ( \43817 , \43812 , \43816 );
or \U$43475 ( \43818 , \43815 , \3918 );
nand \U$43476 ( \43819 , \43817 , \43818 );
and \U$43477 ( \43820 , \43811 , \43819 );
and \U$43478 ( \43821 , \43802 , \43810 );
or \U$43479 ( \43822 , \43820 , \43821 );
and \U$43480 ( \43823 , \2464 , RI986ea58_30);
and \U$43481 ( \43824 , RI986e968_28, \2462 );
nor \U$43482 ( \43825 , \43823 , \43824 );
and \U$43483 ( \43826 , \43825 , \2468 );
not \U$43484 ( \43827 , \43825 );
and \U$43485 ( \43828 , \43827 , \2263 );
nor \U$43486 ( \43829 , \43826 , \43828 );
not \U$43487 ( \43830 , \1462 );
and \U$43488 ( \43831 , \2042 , RI9871848_128);
and \U$43489 ( \43832 , RI9871578_122, \2040 );
nor \U$43490 ( \43833 , \43831 , \43832 );
not \U$43491 ( \43834 , \43833 );
or \U$43492 ( \43835 , \43830 , \43834 );
or \U$43493 ( \43836 , \43833 , \1462 );
nand \U$43494 ( \43837 , \43835 , \43836 );
xor \U$43495 ( \43838 , \43829 , \43837 );
and \U$43496 ( \43839 , \2274 , RI9871668_124);
and \U$43497 ( \43840 , RI986eb48_32, \2272 );
nor \U$43498 ( \43841 , \43839 , \43840 );
and \U$43499 ( \43842 , \43841 , \2030 );
not \U$43500 ( \43843 , \43841 );
and \U$43501 ( \43844 , \43843 , \2031 );
nor \U$43502 ( \43845 , \43842 , \43844 );
and \U$43503 ( \43846 , \43838 , \43845 );
and \U$43504 ( \43847 , \43829 , \43837 );
or \U$43505 ( \43848 , \43846 , \43847 );
xor \U$43506 ( \43849 , \43822 , \43848 );
not \U$43507 ( \43850 , \4521 );
and \U$43508 ( \43851 , \4710 , RI986eff8_42);
and \U$43509 ( \43852 , RI986f2c8_48, \4708 );
nor \U$43510 ( \43853 , \43851 , \43852 );
not \U$43511 ( \43854 , \43853 );
or \U$43512 ( \43855 , \43850 , \43854 );
or \U$43513 ( \43856 , \43853 , \4521 );
nand \U$43514 ( \43857 , \43855 , \43856 );
and \U$43515 ( \43858 , \5318 , RI986f1d8_46);
and \U$43516 ( \43859 , RI986e5a8_20, \5316 );
nor \U$43517 ( \43860 , \43858 , \43859 );
and \U$43518 ( \43861 , \43860 , \5052 );
not \U$43519 ( \43862 , \43860 );
and \U$43520 ( \43863 , \43862 , \5322 );
nor \U$43521 ( \43864 , \43861 , \43863 );
xor \U$43522 ( \43865 , \43857 , \43864 );
and \U$43523 ( \43866 , \5881 , RI986e4b8_18);
and \U$43524 ( \43867 , RI986e788_24, \5879 );
nor \U$43525 ( \43868 , \43866 , \43867 );
and \U$43526 ( \43869 , \43868 , \5594 );
not \U$43527 ( \43870 , \43868 );
and \U$43528 ( \43871 , \43870 , \5885 );
nor \U$43529 ( \43872 , \43869 , \43871 );
and \U$43530 ( \43873 , \43865 , \43872 );
and \U$43531 ( \43874 , \43857 , \43864 );
or \U$43532 ( \43875 , \43873 , \43874 );
and \U$43533 ( \43876 , \43849 , \43875 );
and \U$43534 ( \43877 , \43822 , \43848 );
or \U$43535 ( \43878 , \43876 , \43877 );
and \U$43536 ( \43879 , \43795 , \43878 );
and \U$43537 ( \43880 , \43717 , \43794 );
or \U$43538 ( \43881 , \43879 , \43880 );
xor \U$43539 ( \43882 , \42925 , \42930 );
xor \U$43540 ( \43883 , \43882 , \42938 );
xor \U$43541 ( \43884 , \42900 , \42907 );
xor \U$43542 ( \43885 , \43884 , \42915 );
and \U$43543 ( \43886 , \43883 , \43885 );
xor \U$43544 ( \43887 , \43295 , \11687 );
xor \U$43545 ( \43888 , \43887 , \43303 );
xor \U$43546 ( \43889 , \43314 , \43321 );
xor \U$43547 ( \43890 , \43889 , \43329 );
and \U$43548 ( \43891 , \43888 , \43890 );
xor \U$43549 ( \43892 , \43270 , \43277 );
xor \U$43550 ( \43893 , \43892 , \43285 );
xor \U$43551 ( \43894 , \43314 , \43321 );
xor \U$43552 ( \43895 , \43894 , \43329 );
and \U$43553 ( \43896 , \43893 , \43895 );
and \U$43554 ( \43897 , \43888 , \43893 );
or \U$43555 ( \43898 , \43891 , \43896 , \43897 );
xor \U$43556 ( \43899 , \42900 , \42907 );
xor \U$43557 ( \43900 , \43899 , \42915 );
and \U$43558 ( \43901 , \43898 , \43900 );
and \U$43559 ( \43902 , \43883 , \43898 );
or \U$43560 ( \43903 , \43886 , \43901 , \43902 );
xor \U$43561 ( \43904 , \43881 , \43903 );
xor \U$43562 ( \43905 , \43369 , \43377 );
xor \U$43563 ( \43906 , \43905 , \43386 );
xor \U$43564 ( \43907 , \43343 , \43350 );
xor \U$43565 ( \43908 , \43907 , \43358 );
xor \U$43566 ( \43909 , \43906 , \43908 );
xor \U$43567 ( \43910 , \43397 , \43405 );
xor \U$43568 ( \43911 , \43910 , \43413 );
and \U$43569 ( \43912 , \43909 , \43911 );
and \U$43570 ( \43913 , \43906 , \43908 );
or \U$43571 ( \43914 , \43912 , \43913 );
and \U$43572 ( \43915 , \416 , RI986fe08_72);
and \U$43573 ( \43916 , RI986fd18_70, \414 );
nor \U$43574 ( \43917 , \43915 , \43916 );
and \U$43575 ( \43918 , \43917 , \422 );
not \U$43576 ( \43919 , \43917 );
and \U$43577 ( \43920 , \43919 , \421 );
nor \U$43578 ( \43921 , \43918 , \43920 );
not \U$43579 ( \43922 , RI986fc28_68);
nor \U$43580 ( \43923 , \43922 , \407 );
xor \U$43581 ( \43924 , \43921 , \43923 );
nand \U$43582 ( \43925 , RI986fb38_66, RI9871fc8_144);
and \U$43583 ( \43926 , \416 , RI986fc28_68);
and \U$43584 ( \43927 , RI986fe08_72, \414 );
nor \U$43585 ( \43928 , \43926 , \43927 );
and \U$43586 ( \43929 , \43928 , \421 );
not \U$43587 ( \43930 , \43928 );
and \U$43588 ( \43931 , \43930 , \422 );
nor \U$43589 ( \43932 , \43929 , \43931 );
nand \U$43590 ( \43933 , \43925 , \43932 );
and \U$43591 ( \43934 , \43924 , \43933 );
and \U$43592 ( \43935 , \43921 , \43923 );
or \U$43593 ( \43936 , \43934 , \43935 );
xor \U$43594 ( \43937 , \43914 , \43936 );
xor \U$43595 ( \43938 , \43454 , \43461 );
xor \U$43596 ( \43939 , \43938 , \43469 );
xor \U$43597 ( \43940 , \43481 , \43489 );
xor \U$43598 ( \43941 , \43940 , \43497 );
and \U$43599 ( \43942 , \43939 , \43941 );
xor \U$43600 ( \43943 , \43428 , \43435 );
xor \U$43601 ( \43944 , \43943 , \43443 );
xor \U$43602 ( \43945 , \43481 , \43489 );
xor \U$43603 ( \43946 , \43945 , \43497 );
and \U$43604 ( \43947 , \43944 , \43946 );
and \U$43605 ( \43948 , \43939 , \43944 );
or \U$43606 ( \43949 , \43942 , \43947 , \43948 );
and \U$43607 ( \43950 , \43937 , \43949 );
and \U$43608 ( \43951 , \43914 , \43936 );
or \U$43609 ( \43952 , \43950 , \43951 );
and \U$43610 ( \43953 , \43904 , \43952 );
and \U$43611 ( \43954 , \43881 , \43903 );
or \U$43612 ( \43955 , \43953 , \43954 );
xor \U$43613 ( \43956 , \43633 , \43955 );
xor \U$43614 ( \43957 , \42997 , \43026 );
xor \U$43615 ( \43958 , \43957 , \43053 );
xor \U$43616 ( \43959 , \43203 , \43210 );
xor \U$43617 ( \43960 , \43958 , \43959 );
xor \U$43618 ( \43961 , \43237 , \43249 );
xor \U$43619 ( \43962 , \43961 , \43260 );
and \U$43620 ( \43963 , \43960 , \43962 );
xor \U$43621 ( \43964 , \42882 , \42884 );
xor \U$43622 ( \43965 , \43964 , \42887 );
xor \U$43623 ( \43966 , \43509 , \43516 );
xor \U$43624 ( \43967 , \43965 , \43966 );
xor \U$43625 ( \43968 , \43237 , \43249 );
xor \U$43626 ( \43969 , \43968 , \43260 );
and \U$43627 ( \43970 , \43967 , \43969 );
and \U$43628 ( \43971 , \43960 , \43967 );
or \U$43629 ( \43972 , \43963 , \43970 , \43971 );
and \U$43630 ( \43973 , \43956 , \43972 );
and \U$43631 ( \43974 , \43633 , \43955 );
or \U$43632 ( \43975 , \43973 , \43974 );
xor \U$43633 ( \43976 , \43603 , \43975 );
xor \U$43634 ( \43977 , \42893 , \43143 );
xor \U$43635 ( \43978 , \43977 , \43158 );
xor \U$43636 ( \43979 , \43543 , \43550 );
xor \U$43637 ( \43980 , \43978 , \43979 );
and \U$43638 ( \43981 , \43976 , \43980 );
and \U$43639 ( \43982 , \43603 , \43975 );
or \U$43640 ( \43983 , \43981 , \43982 );
xor \U$43641 ( \43984 , \43161 , \43166 );
xor \U$43642 ( \43985 , \43984 , \43191 );
xor \U$43643 ( \43986 , \43983 , \43985 );
xor \U$43644 ( \43987 , \43542 , \43555 );
xor \U$43645 ( \43988 , \43987 , \43560 );
and \U$43646 ( \43989 , \43986 , \43988 );
and \U$43647 ( \43990 , \43983 , \43985 );
or \U$43648 ( \43991 , \43989 , \43990 );
xor \U$43649 ( \43992 , \42855 , \43194 );
xor \U$43650 ( \43993 , \43992 , \43199 );
xor \U$43651 ( \43994 , \42842 , \43563 );
xor \U$43652 ( \43995 , \43993 , \43994 );
and \U$43653 ( \43996 , \43991 , \43995 );
xor \U$43654 ( \43997 , \43568 , \43578 );
and \U$43655 ( \43998 , \43996 , \43997 );
xor \U$43656 ( \43999 , \43996 , \43997 );
xor \U$43657 ( \44000 , \43225 , \43524 );
xor \U$43658 ( \44001 , \44000 , \43539 );
xor \U$43659 ( \44002 , \43603 , \43975 );
xor \U$43660 ( \44003 , \44002 , \43980 );
and \U$43661 ( \44004 , \44001 , \44003 );
xor \U$43662 ( \44005 , \43335 , \43419 );
xor \U$43663 ( \44006 , \44005 , \43503 );
xor \U$43664 ( \44007 , \43613 , \43615 );
xor \U$43665 ( \44008 , \44007 , \43630 );
and \U$43666 ( \44009 , \44006 , \44008 );
xor \U$43667 ( \44010 , \43237 , \43249 );
xor \U$43668 ( \44011 , \44010 , \43260 );
xor \U$43669 ( \44012 , \43960 , \43967 );
xor \U$43670 ( \44013 , \44011 , \44012 );
xor \U$43671 ( \44014 , \43613 , \43615 );
xor \U$43672 ( \44015 , \44014 , \43630 );
and \U$43673 ( \44016 , \44013 , \44015 );
and \U$43674 ( \44017 , \44006 , \44013 );
or \U$43675 ( \44018 , \44009 , \44016 , \44017 );
xor \U$43676 ( \44019 , \43914 , \43936 );
xor \U$43677 ( \44020 , \44019 , \43949 );
xor \U$43678 ( \44021 , \43717 , \43794 );
xor \U$43679 ( \44022 , \44021 , \43878 );
xor \U$43680 ( \44023 , \44020 , \44022 );
xor \U$43681 ( \44024 , \42900 , \42907 );
xor \U$43682 ( \44025 , \44024 , \42915 );
xor \U$43683 ( \44026 , \43883 , \43898 );
xor \U$43684 ( \44027 , \44025 , \44026 );
and \U$43685 ( \44028 , \44023 , \44027 );
and \U$43686 ( \44029 , \44020 , \44022 );
or \U$43687 ( \44030 , \44028 , \44029 );
xor \U$43688 ( \44031 , \43641 , \43648 );
xor \U$43689 ( \44032 , \44031 , \43656 );
xor \U$43690 ( \44033 , \43695 , \43703 );
xor \U$43691 ( \44034 , \44033 , \43711 );
xor \U$43692 ( \44035 , \44032 , \44034 );
xor \U$43693 ( \44036 , \43829 , \43837 );
xor \U$43694 ( \44037 , \44036 , \43845 );
and \U$43695 ( \44038 , \44035 , \44037 );
and \U$43696 ( \44039 , \44032 , \44034 );
or \U$43697 ( \44040 , \44038 , \44039 );
not \U$43698 ( \44041 , \361 );
and \U$43699 ( \44042 , \354 , RI986fe08_72);
and \U$43700 ( \44043 , RI986fd18_70, \352 );
nor \U$43701 ( \44044 , \44042 , \44043 );
not \U$43702 ( \44045 , \44044 );
or \U$43703 ( \44046 , \44041 , \44045 );
or \U$43704 ( \44047 , \44044 , \345 );
nand \U$43705 ( \44048 , \44046 , \44047 );
not \U$43706 ( \44049 , RI9870858_94);
nor \U$43707 ( \44050 , \44049 , \407 );
xor \U$43708 ( \44051 , \44048 , \44050 );
and \U$43709 ( \44052 , \416 , RI986fb38_66);
and \U$43710 ( \44053 , RI986fc28_68, \414 );
nor \U$43711 ( \44054 , \44052 , \44053 );
and \U$43712 ( \44055 , \44054 , \422 );
not \U$43713 ( \44056 , \44054 );
and \U$43714 ( \44057 , \44056 , \421 );
nor \U$43715 ( \44058 , \44055 , \44057 );
and \U$43716 ( \44059 , \44051 , \44058 );
and \U$43717 ( \44060 , \44048 , \44050 );
or \U$43718 ( \44061 , \44059 , \44060 );
or \U$43719 ( \44062 , \43932 , \43925 );
nand \U$43720 ( \44063 , \44062 , \43933 );
xor \U$43721 ( \44064 , \44061 , \44063 );
xor \U$43722 ( \44065 , \43667 , \43675 );
xor \U$43723 ( \44066 , \44065 , \43684 );
and \U$43724 ( \44067 , \44064 , \44066 );
and \U$43725 ( \44068 , \44061 , \44063 );
or \U$43726 ( \44069 , \44067 , \44068 );
xor \U$43727 ( \44070 , \44040 , \44069 );
xor \U$43728 ( \44071 , \43857 , \43864 );
xor \U$43729 ( \44072 , \44071 , \43872 );
xor \U$43730 ( \44073 , \43802 , \43810 );
xor \U$43731 ( \44074 , \44073 , \43819 );
and \U$43732 ( \44075 , \44072 , \44074 );
xor \U$43733 ( \44076 , \43773 , \43780 );
xor \U$43734 ( \44077 , \44076 , \43788 );
xor \U$43735 ( \44078 , \43802 , \43810 );
xor \U$43736 ( \44079 , \44078 , \43819 );
and \U$43737 ( \44080 , \44077 , \44079 );
and \U$43738 ( \44081 , \44072 , \44077 );
or \U$43739 ( \44082 , \44075 , \44080 , \44081 );
and \U$43740 ( \44083 , \44070 , \44082 );
and \U$43741 ( \44084 , \44040 , \44069 );
or \U$43742 ( \44085 , \44083 , \44084 );
and \U$43743 ( \44086 , \1329 , RI98712a8_116);
and \U$43744 ( \44087 , RI98711b8_114, \1327 );
nor \U$43745 ( \44088 , \44086 , \44087 );
and \U$43746 ( \44089 , \44088 , \1336 );
not \U$43747 ( \44090 , \44088 );
and \U$43748 ( \44091 , \44090 , \1337 );
nor \U$43749 ( \44092 , \44089 , \44091 );
and \U$43750 ( \44093 , \1311 , RI9871398_118);
and \U$43751 ( \44094 , RI9871488_120, \1309 );
nor \U$43752 ( \44095 , \44093 , \44094 );
and \U$43753 ( \44096 , \44095 , \1458 );
not \U$43754 ( \44097 , \44095 );
and \U$43755 ( \44098 , \44097 , \1318 );
nor \U$43756 ( \44099 , \44096 , \44098 );
xor \U$43757 ( \44100 , \44092 , \44099 );
not \U$43758 ( \44101 , \1462 );
and \U$43759 ( \44102 , \2042 , RI9871758_126);
and \U$43760 ( \44103 , RI9871848_128, \2040 );
nor \U$43761 ( \44104 , \44102 , \44103 );
not \U$43762 ( \44105 , \44104 );
or \U$43763 ( \44106 , \44101 , \44105 );
or \U$43764 ( \44107 , \44104 , \2034 );
nand \U$43765 ( \44108 , \44106 , \44107 );
and \U$43766 ( \44109 , \44100 , \44108 );
and \U$43767 ( \44110 , \44092 , \44099 );
or \U$43768 ( \44111 , \44109 , \44110 );
not \U$43769 ( \44112 , \386 );
and \U$43770 ( \44113 , \395 , RI986ffe8_76);
and \U$43771 ( \44114 , RI986fef8_74, \393 );
nor \U$43772 ( \44115 , \44113 , \44114 );
not \U$43773 ( \44116 , \44115 );
or \U$43774 ( \44117 , \44112 , \44116 );
or \U$43775 ( \44118 , \44115 , \386 );
nand \U$43776 ( \44119 , \44117 , \44118 );
not \U$43777 ( \44120 , \454 );
and \U$43778 ( \44121 , \465 , RI9870fd8_110);
and \U$43779 ( \44122 , RI9870b28_100, \463 );
nor \U$43780 ( \44123 , \44121 , \44122 );
not \U$43781 ( \44124 , \44123 );
or \U$43782 ( \44125 , \44120 , \44124 );
or \U$43783 ( \44126 , \44123 , \454 );
nand \U$43784 ( \44127 , \44125 , \44126 );
xor \U$43785 ( \44128 , \44119 , \44127 );
not \U$43786 ( \44129 , \365 );
and \U$43787 ( \44130 , \376 , RI98700d8_78);
and \U$43788 ( \44131 , RI98701c8_80, \374 );
nor \U$43789 ( \44132 , \44130 , \44131 );
not \U$43790 ( \44133 , \44132 );
or \U$43791 ( \44134 , \44129 , \44133 );
or \U$43792 ( \44135 , \44132 , \365 );
nand \U$43793 ( \44136 , \44134 , \44135 );
and \U$43794 ( \44137 , \44128 , \44136 );
and \U$43795 ( \44138 , \44119 , \44127 );
or \U$43796 ( \44139 , \44137 , \44138 );
xor \U$43797 ( \44140 , \44111 , \44139 );
not \U$43798 ( \44141 , \1128 );
and \U$43799 ( \44142 , \1293 , RI98710c8_112);
and \U$43800 ( \44143 , RI9870d08_104, \1291 );
nor \U$43801 ( \44144 , \44142 , \44143 );
not \U$43802 ( \44145 , \44144 );
or \U$43803 ( \44146 , \44141 , \44145 );
or \U$43804 ( \44147 , \44144 , \1128 );
nand \U$43805 ( \44148 , \44146 , \44147 );
and \U$43806 ( \44149 , \776 , RI9870ee8_108);
and \U$43807 ( \44150 , RI9870c18_102, \774 );
nor \U$43808 ( \44151 , \44149 , \44150 );
and \U$43809 ( \44152 , \44151 , \474 );
not \U$43810 ( \44153 , \44151 );
and \U$43811 ( \44154 , \44153 , \451 );
nor \U$43812 ( \44155 , \44152 , \44154 );
xor \U$43813 ( \44156 , \44148 , \44155 );
and \U$43814 ( \44157 , \438 , RI9870df8_106);
and \U$43815 ( \44158 , RI9870a38_98, \436 );
nor \U$43816 ( \44159 , \44157 , \44158 );
and \U$43817 ( \44160 , \44159 , \444 );
not \U$43818 ( \44161 , \44159 );
and \U$43819 ( \44162 , \44161 , \443 );
nor \U$43820 ( \44163 , \44160 , \44162 );
and \U$43821 ( \44164 , \44156 , \44163 );
and \U$43822 ( \44165 , \44148 , \44155 );
or \U$43823 ( \44166 , \44164 , \44165 );
and \U$43824 ( \44167 , \44140 , \44166 );
and \U$43825 ( \44168 , \44111 , \44139 );
or \U$43826 ( \44169 , \44167 , \44168 );
and \U$43827 ( \44170 , \10424 , RI986de28_4);
and \U$43828 ( \44171 , RI986dd38_2, \10422 );
nor \U$43829 ( \44172 , \44170 , \44171 );
and \U$43830 ( \44173 , \44172 , \9840 );
not \U$43831 ( \44174 , \44172 );
and \U$43832 ( \44175 , \44174 , \10428 );
nor \U$43833 ( \44176 , \44173 , \44175 );
and \U$43834 ( \44177 , \9237 , RI986f598_54);
and \U$43835 ( \44178 , RI986f688_56, \9235 );
nor \U$43836 ( \44179 , \44177 , \44178 );
and \U$43837 ( \44180 , \44179 , \9241 );
not \U$43838 ( \44181 , \44179 );
and \U$43839 ( \44182 , \44181 , \8836 );
nor \U$43840 ( \44183 , \44180 , \44182 );
xor \U$43841 ( \44184 , \44176 , \44183 );
and \U$43842 ( \44185 , \9505 , RI986e008_8);
and \U$43843 ( \44186 , RI986df18_6, \9503 );
nor \U$43844 ( \44187 , \44185 , \44186 );
and \U$43845 ( \44188 , \44187 , \9510 );
not \U$43846 ( \44189 , \44187 );
and \U$43847 ( \44190 , \44189 , \9513 );
nor \U$43848 ( \44191 , \44188 , \44190 );
and \U$43849 ( \44192 , \44184 , \44191 );
and \U$43850 ( \44193 , \44176 , \44183 );
or \U$43851 ( \44194 , \44192 , \44193 );
and \U$43852 ( \44195 , \11696 , RI986e1e8_12);
and \U$43853 ( \44196 , RI986e0f8_10, \11694 );
nor \U$43854 ( \44197 , \44195 , \44196 );
and \U$43855 ( \44198 , \44197 , \10965 );
not \U$43856 ( \44199 , \44197 );
and \U$43857 ( \44200 , \44199 , \11702 );
nor \U$43858 ( \44201 , \44198 , \44200 );
xor \U$43859 ( \44202 , \44201 , \13047 );
and \U$43860 ( \44203 , \12293 , RI986e2d8_14);
and \U$43861 ( \44204 , RI986e3c8_16, \12291 );
nor \U$43862 ( \44205 , \44203 , \44204 );
and \U$43863 ( \44206 , \44205 , \11687 );
not \U$43864 ( \44207 , \44205 );
and \U$43865 ( \44208 , \44207 , \11686 );
nor \U$43866 ( \44209 , \44206 , \44208 );
and \U$43867 ( \44210 , \44202 , \44209 );
and \U$43868 ( \44211 , \44201 , \13047 );
or \U$43869 ( \44212 , \44210 , \44211 );
xor \U$43870 ( \44213 , \44194 , \44212 );
and \U$43871 ( \44214 , \7729 , RI986fa48_64);
and \U$43872 ( \44215 , RI986f958_62, \7727 );
nor \U$43873 ( \44216 , \44214 , \44215 );
and \U$43874 ( \44217 , \44216 , \7480 );
not \U$43875 ( \44218 , \44216 );
and \U$43876 ( \44219 , \44218 , \7733 );
nor \U$43877 ( \44220 , \44217 , \44219 );
and \U$43878 ( \44221 , \7079 , RI986f868_60);
and \U$43879 ( \44222 , RI986f778_58, \7077 );
nor \U$43880 ( \44223 , \44221 , \44222 );
and \U$43881 ( \44224 , \44223 , \6710 );
not \U$43882 ( \44225 , \44223 );
and \U$43883 ( \44226 , \44225 , \6709 );
nor \U$43884 ( \44227 , \44224 , \44226 );
xor \U$43885 ( \44228 , \44220 , \44227 );
and \U$43886 ( \44229 , \8486 , RI986f4a8_52);
and \U$43887 ( \44230 , RI986f3b8_50, \8484 );
nor \U$43888 ( \44231 , \44229 , \44230 );
and \U$43889 ( \44232 , \44231 , \8050 );
not \U$43890 ( \44233 , \44231 );
and \U$43891 ( \44234 , \44233 , \8051 );
nor \U$43892 ( \44235 , \44232 , \44234 );
and \U$43893 ( \44236 , \44228 , \44235 );
and \U$43894 ( \44237 , \44220 , \44227 );
or \U$43895 ( \44238 , \44236 , \44237 );
and \U$43896 ( \44239 , \44213 , \44238 );
and \U$43897 ( \44240 , \44194 , \44212 );
or \U$43898 ( \44241 , \44239 , \44240 );
xor \U$43899 ( \44242 , \44169 , \44241 );
not \U$43900 ( \44243 , \3918 );
and \U$43901 ( \44244 , \3683 , RI986ef08_40);
and \U$43902 ( \44245 , RI986ee18_38, \3681 );
nor \U$43903 ( \44246 , \44244 , \44245 );
not \U$43904 ( \44247 , \44246 );
or \U$43905 ( \44248 , \44243 , \44247 );
or \U$43906 ( \44249 , \44246 , \3412 );
nand \U$43907 ( \44250 , \44248 , \44249 );
and \U$43908 ( \44251 , \4203 , RI986ec38_34);
and \U$43909 ( \44252 , RI986ed28_36, \4201 );
nor \U$43910 ( \44253 , \44251 , \44252 );
and \U$43911 ( \44254 , \44253 , \4207 );
not \U$43912 ( \44255 , \44253 );
and \U$43913 ( \44256 , \44255 , \3923 );
nor \U$43914 ( \44257 , \44254 , \44256 );
xor \U$43915 ( \44258 , \44250 , \44257 );
not \U$43916 ( \44259 , \4521 );
and \U$43917 ( \44260 , \4710 , RI986f0e8_44);
and \U$43918 ( \44261 , RI986eff8_42, \4708 );
nor \U$43919 ( \44262 , \44260 , \44261 );
not \U$43920 ( \44263 , \44262 );
or \U$43921 ( \44264 , \44259 , \44263 );
or \U$43922 ( \44265 , \44262 , \4521 );
nand \U$43923 ( \44266 , \44264 , \44265 );
and \U$43924 ( \44267 , \44258 , \44266 );
and \U$43925 ( \44268 , \44250 , \44257 );
or \U$43926 ( \44269 , \44267 , \44268 );
and \U$43927 ( \44270 , \2274 , RI9871578_122);
and \U$43928 ( \44271 , RI9871668_124, \2272 );
nor \U$43929 ( \44272 , \44270 , \44271 );
and \U$43930 ( \44273 , \44272 , \2030 );
not \U$43931 ( \44274 , \44272 );
and \U$43932 ( \44275 , \44274 , \2031 );
nor \U$43933 ( \44276 , \44273 , \44275 );
and \U$43934 ( \44277 , \2464 , RI986eb48_32);
and \U$43935 ( \44278 , RI986ea58_30, \2462 );
nor \U$43936 ( \44279 , \44277 , \44278 );
and \U$43937 ( \44280 , \44279 , \2468 );
not \U$43938 ( \44281 , \44279 );
and \U$43939 ( \44282 , \44281 , \2263 );
nor \U$43940 ( \44283 , \44280 , \44282 );
xor \U$43941 ( \44284 , \44276 , \44283 );
not \U$43942 ( \44285 , \3406 );
and \U$43943 ( \44286 , \3254 , RI986e968_28);
and \U$43944 ( \44287 , RI986e878_26, \3252 );
nor \U$43945 ( \44288 , \44286 , \44287 );
not \U$43946 ( \44289 , \44288 );
or \U$43947 ( \44290 , \44285 , \44289 );
or \U$43948 ( \44291 , \44288 , \3406 );
nand \U$43949 ( \44292 , \44290 , \44291 );
and \U$43950 ( \44293 , \44284 , \44292 );
and \U$43951 ( \44294 , \44276 , \44283 );
or \U$43952 ( \44295 , \44293 , \44294 );
xor \U$43953 ( \44296 , \44269 , \44295 );
and \U$43954 ( \44297 , \5318 , RI986f2c8_48);
and \U$43955 ( \44298 , RI986f1d8_46, \5316 );
nor \U$43956 ( \44299 , \44297 , \44298 );
and \U$43957 ( \44300 , \44299 , \5052 );
not \U$43958 ( \44301 , \44299 );
and \U$43959 ( \44302 , \44301 , \5322 );
nor \U$43960 ( \44303 , \44300 , \44302 );
and \U$43961 ( \44304 , \5881 , RI986e5a8_20);
and \U$43962 ( \44305 , RI986e4b8_18, \5879 );
nor \U$43963 ( \44306 , \44304 , \44305 );
and \U$43964 ( \44307 , \44306 , \5594 );
not \U$43965 ( \44308 , \44306 );
and \U$43966 ( \44309 , \44308 , \5885 );
nor \U$43967 ( \44310 , \44307 , \44309 );
xor \U$43968 ( \44311 , \44303 , \44310 );
and \U$43969 ( \44312 , \6453 , RI986e788_24);
and \U$43970 ( \44313 , RI986e698_22, \6451 );
nor \U$43971 ( \44314 , \44312 , \44313 );
and \U$43972 ( \44315 , \44314 , \6190 );
not \U$43973 ( \44316 , \44314 );
and \U$43974 ( \44317 , \44316 , \6705 );
nor \U$43975 ( \44318 , \44315 , \44317 );
and \U$43976 ( \44319 , \44311 , \44318 );
and \U$43977 ( \44320 , \44303 , \44310 );
or \U$43978 ( \44321 , \44319 , \44320 );
and \U$43979 ( \44322 , \44296 , \44321 );
and \U$43980 ( \44323 , \44269 , \44295 );
or \U$43981 ( \44324 , \44322 , \44323 );
and \U$43982 ( \44325 , \44242 , \44324 );
and \U$43983 ( \44326 , \44169 , \44241 );
or \U$43984 ( \44327 , \44325 , \44326 );
xor \U$43985 ( \44328 , \44085 , \44327 );
xor \U$43986 ( \44329 , \43314 , \43321 );
xor \U$43987 ( \44330 , \44329 , \43329 );
xor \U$43988 ( \44331 , \43888 , \43893 );
xor \U$43989 ( \44332 , \44330 , \44331 );
xor \U$43990 ( \44333 , \43906 , \43908 );
xor \U$43991 ( \44334 , \44333 , \43911 );
and \U$43992 ( \44335 , \44332 , \44334 );
xor \U$43993 ( \44336 , \43481 , \43489 );
xor \U$43994 ( \44337 , \44336 , \43497 );
xor \U$43995 ( \44338 , \43939 , \43944 );
xor \U$43996 ( \44339 , \44337 , \44338 );
xor \U$43997 ( \44340 , \43906 , \43908 );
xor \U$43998 ( \44341 , \44340 , \43911 );
and \U$43999 ( \44342 , \44339 , \44341 );
and \U$44000 ( \44343 , \44332 , \44339 );
or \U$44001 ( \44344 , \44335 , \44342 , \44343 );
and \U$44002 ( \44345 , \44328 , \44344 );
and \U$44003 ( \44346 , \44085 , \44327 );
or \U$44004 ( \44347 , \44345 , \44346 );
xor \U$44005 ( \44348 , \44030 , \44347 );
xor \U$44006 ( \44349 , \43921 , \43923 );
xor \U$44007 ( \44350 , \44349 , \43933 );
xor \U$44008 ( \44351 , \43659 , \43687 );
xor \U$44009 ( \44352 , \44351 , \43714 );
and \U$44010 ( \44353 , \44350 , \44352 );
xor \U$44011 ( \44354 , \43822 , \43848 );
xor \U$44012 ( \44355 , \44354 , \43875 );
xor \U$44013 ( \44356 , \43659 , \43687 );
xor \U$44014 ( \44357 , \44356 , \43714 );
and \U$44015 ( \44358 , \44355 , \44357 );
and \U$44016 ( \44359 , \44350 , \44355 );
or \U$44017 ( \44360 , \44353 , \44358 , \44359 );
xor \U$44018 ( \44361 , \43605 , \43607 );
xor \U$44019 ( \44362 , \44361 , \43610 );
and \U$44020 ( \44363 , \44360 , \44362 );
xor \U$44021 ( \44364 , \43252 , \43254 );
xor \U$44022 ( \44365 , \44364 , \43257 );
xor \U$44023 ( \44366 , \43618 , \43625 );
xor \U$44024 ( \44367 , \44365 , \44366 );
xor \U$44025 ( \44368 , \43605 , \43607 );
xor \U$44026 ( \44369 , \44368 , \43610 );
and \U$44027 ( \44370 , \44367 , \44369 );
and \U$44028 ( \44371 , \44360 , \44367 );
or \U$44029 ( \44372 , \44363 , \44370 , \44371 );
and \U$44030 ( \44373 , \44348 , \44372 );
and \U$44031 ( \44374 , \44030 , \44347 );
or \U$44032 ( \44375 , \44373 , \44374 );
xor \U$44033 ( \44376 , \44018 , \44375 );
xor \U$44034 ( \44377 , \43215 , \43217 );
xor \U$44035 ( \44378 , \44377 , \43222 );
xor \U$44036 ( \44379 , \43591 , \43598 );
xor \U$44037 ( \44380 , \44378 , \44379 );
and \U$44038 ( \44381 , \44376 , \44380 );
and \U$44039 ( \44382 , \44018 , \44375 );
or \U$44040 ( \44383 , \44381 , \44382 );
xor \U$44041 ( \44384 , \43603 , \43975 );
xor \U$44042 ( \44385 , \44384 , \43980 );
and \U$44043 ( \44386 , \44383 , \44385 );
and \U$44044 ( \44387 , \44001 , \44383 );
or \U$44045 ( \44388 , \44004 , \44386 , \44387 );
xor \U$44046 ( \44389 , \43983 , \43985 );
xor \U$44047 ( \44390 , \44389 , \43988 );
and \U$44048 ( \44391 , \44388 , \44390 );
not \U$44049 ( \44392 , \44391 );
xor \U$44050 ( \44393 , \43991 , \43995 );
not \U$44051 ( \44394 , \44393 );
or \U$44052 ( \44395 , \44392 , \44394 );
xor \U$44053 ( \44396 , \44018 , \44375 );
xor \U$44054 ( \44397 , \44396 , \44380 );
xor \U$44055 ( \44398 , \44169 , \44241 );
xor \U$44056 ( \44399 , \44398 , \44324 );
xor \U$44057 ( \44400 , \44040 , \44069 );
xor \U$44058 ( \44401 , \44400 , \44082 );
and \U$44059 ( \44402 , \44399 , \44401 );
xor \U$44060 ( \44403 , \43906 , \43908 );
xor \U$44061 ( \44404 , \44403 , \43911 );
xor \U$44062 ( \44405 , \44332 , \44339 );
xor \U$44063 ( \44406 , \44404 , \44405 );
xor \U$44064 ( \44407 , \44040 , \44069 );
xor \U$44065 ( \44408 , \44407 , \44082 );
and \U$44066 ( \44409 , \44406 , \44408 );
and \U$44067 ( \44410 , \44399 , \44406 );
or \U$44068 ( \44411 , \44402 , \44409 , \44410 );
xor \U$44069 ( \44412 , \43724 , \43731 );
xor \U$44070 ( \44413 , \44412 , \43739 );
xor \U$44071 ( \44414 , \43749 , \43754 );
xor \U$44072 ( \44415 , \44414 , \43762 );
xor \U$44073 ( \44416 , \44413 , \44415 );
xor \U$44074 ( \44417 , \43802 , \43810 );
xor \U$44075 ( \44418 , \44417 , \43819 );
xor \U$44076 ( \44419 , \44072 , \44077 );
xor \U$44077 ( \44420 , \44418 , \44419 );
and \U$44078 ( \44421 , \44416 , \44420 );
and \U$44079 ( \44422 , \44413 , \44415 );
or \U$44080 ( \44423 , \44421 , \44422 );
not \U$44081 ( \44424 , \1301 );
and \U$44082 ( \44425 , \1293 , RI9870c18_102);
and \U$44083 ( \44426 , RI98710c8_112, \1291 );
nor \U$44084 ( \44427 , \44425 , \44426 );
not \U$44085 ( \44428 , \44427 );
or \U$44086 ( \44429 , \44424 , \44428 );
or \U$44087 ( \44430 , \44427 , \1301 );
nand \U$44088 ( \44431 , \44429 , \44430 );
and \U$44089 ( \44432 , \776 , RI9870a38_98);
and \U$44090 ( \44433 , RI9870ee8_108, \774 );
nor \U$44091 ( \44434 , \44432 , \44433 );
and \U$44092 ( \44435 , \44434 , \474 );
not \U$44093 ( \44436 , \44434 );
and \U$44094 ( \44437 , \44436 , \451 );
nor \U$44095 ( \44438 , \44435 , \44437 );
xor \U$44096 ( \44439 , \44431 , \44438 );
and \U$44097 ( \44440 , \438 , RI9870b28_100);
and \U$44098 ( \44441 , RI9870df8_106, \436 );
nor \U$44099 ( \44442 , \44440 , \44441 );
and \U$44100 ( \44443 , \44442 , \444 );
not \U$44101 ( \44444 , \44442 );
and \U$44102 ( \44445 , \44444 , \443 );
nor \U$44103 ( \44446 , \44443 , \44445 );
and \U$44104 ( \44447 , \44439 , \44446 );
and \U$44105 ( \44448 , \44431 , \44438 );
or \U$44106 ( \44449 , \44447 , \44448 );
not \U$44107 ( \44450 , \367 );
and \U$44108 ( \44451 , \376 , RI986fef8_74);
and \U$44109 ( \44452 , RI98700d8_78, \374 );
nor \U$44110 ( \44453 , \44451 , \44452 );
not \U$44111 ( \44454 , \44453 );
or \U$44112 ( \44455 , \44450 , \44454 );
or \U$44113 ( \44456 , \44453 , \367 );
nand \U$44114 ( \44457 , \44455 , \44456 );
not \U$44115 ( \44458 , \454 );
and \U$44116 ( \44459 , \465 , RI98701c8_80);
and \U$44117 ( \44460 , RI9870fd8_110, \463 );
nor \U$44118 ( \44461 , \44459 , \44460 );
not \U$44119 ( \44462 , \44461 );
or \U$44120 ( \44463 , \44458 , \44462 );
or \U$44121 ( \44464 , \44461 , \454 );
nand \U$44122 ( \44465 , \44463 , \44464 );
xor \U$44123 ( \44466 , \44457 , \44465 );
not \U$44124 ( \44467 , \386 );
and \U$44125 ( \44468 , \395 , RI986fd18_70);
and \U$44126 ( \44469 , RI986ffe8_76, \393 );
nor \U$44127 ( \44470 , \44468 , \44469 );
not \U$44128 ( \44471 , \44470 );
or \U$44129 ( \44472 , \44467 , \44471 );
or \U$44130 ( \44473 , \44470 , \487 );
nand \U$44131 ( \44474 , \44472 , \44473 );
and \U$44132 ( \44475 , \44466 , \44474 );
and \U$44133 ( \44476 , \44457 , \44465 );
or \U$44134 ( \44477 , \44475 , \44476 );
xor \U$44135 ( \44478 , \44449 , \44477 );
and \U$44136 ( \44479 , \1311 , RI98711b8_114);
and \U$44137 ( \44480 , RI9871398_118, \1309 );
nor \U$44138 ( \44481 , \44479 , \44480 );
and \U$44139 ( \44482 , \44481 , \1458 );
not \U$44140 ( \44483 , \44481 );
and \U$44141 ( \44484 , \44483 , \1318 );
nor \U$44142 ( \44485 , \44482 , \44484 );
and \U$44143 ( \44486 , \1329 , RI9870d08_104);
and \U$44144 ( \44487 , RI98712a8_116, \1327 );
nor \U$44145 ( \44488 , \44486 , \44487 );
and \U$44146 ( \44489 , \44488 , \1336 );
not \U$44147 ( \44490 , \44488 );
and \U$44148 ( \44491 , \44490 , \1337 );
nor \U$44149 ( \44492 , \44489 , \44491 );
xor \U$44150 ( \44493 , \44485 , \44492 );
not \U$44151 ( \44494 , \1462 );
and \U$44152 ( \44495 , \2042 , RI9871488_120);
and \U$44153 ( \44496 , RI9871758_126, \2040 );
nor \U$44154 ( \44497 , \44495 , \44496 );
not \U$44155 ( \44498 , \44497 );
or \U$44156 ( \44499 , \44494 , \44498 );
or \U$44157 ( \44500 , \44497 , \1462 );
nand \U$44158 ( \44501 , \44499 , \44500 );
and \U$44159 ( \44502 , \44493 , \44501 );
and \U$44160 ( \44503 , \44485 , \44492 );
or \U$44161 ( \44504 , \44502 , \44503 );
and \U$44162 ( \44505 , \44478 , \44504 );
and \U$44163 ( \44506 , \44449 , \44477 );
or \U$44164 ( \44507 , \44505 , \44506 );
and \U$44165 ( \44508 , \7079 , RI986e698_22);
and \U$44166 ( \44509 , RI986f868_60, \7077 );
nor \U$44167 ( \44510 , \44508 , \44509 );
and \U$44168 ( \44511 , \44510 , \6710 );
not \U$44169 ( \44512 , \44510 );
and \U$44170 ( \44513 , \44512 , \6709 );
nor \U$44171 ( \44514 , \44511 , \44513 );
and \U$44172 ( \44515 , \7729 , RI986f778_58);
and \U$44173 ( \44516 , RI986fa48_64, \7727 );
nor \U$44174 ( \44517 , \44515 , \44516 );
and \U$44175 ( \44518 , \44517 , \7480 );
not \U$44176 ( \44519 , \44517 );
and \U$44177 ( \44520 , \44519 , \7733 );
nor \U$44178 ( \44521 , \44518 , \44520 );
xor \U$44179 ( \44522 , \44514 , \44521 );
and \U$44180 ( \44523 , \8486 , RI986f958_62);
and \U$44181 ( \44524 , RI986f4a8_52, \8484 );
nor \U$44182 ( \44525 , \44523 , \44524 );
and \U$44183 ( \44526 , \44525 , \8050 );
not \U$44184 ( \44527 , \44525 );
and \U$44185 ( \44528 , \44527 , \8051 );
nor \U$44186 ( \44529 , \44526 , \44528 );
and \U$44187 ( \44530 , \44522 , \44529 );
and \U$44188 ( \44531 , \44514 , \44521 );
or \U$44189 ( \44532 , \44530 , \44531 );
and \U$44190 ( \44533 , \11696 , RI986dd38_2);
and \U$44191 ( \44534 , RI986e1e8_12, \11694 );
nor \U$44192 ( \44535 , \44533 , \44534 );
and \U$44193 ( \44536 , \44535 , \10965 );
not \U$44194 ( \44537 , \44535 );
and \U$44195 ( \44538 , \44537 , \11702 );
nor \U$44196 ( \44539 , \44536 , \44538 );
nand \U$44197 ( \44540 , RI986e3c8_16, \13045 );
and \U$44198 ( \44541 , \44540 , \13047 );
not \U$44199 ( \44542 , \44540 );
and \U$44200 ( \44543 , \44542 , \12619 );
nor \U$44201 ( \44544 , \44541 , \44543 );
xor \U$44202 ( \44545 , \44539 , \44544 );
and \U$44203 ( \44546 , \12293 , RI986e0f8_10);
and \U$44204 ( \44547 , RI986e2d8_14, \12291 );
nor \U$44205 ( \44548 , \44546 , \44547 );
and \U$44206 ( \44549 , \44548 , \11687 );
not \U$44207 ( \44550 , \44548 );
and \U$44208 ( \44551 , \44550 , \11686 );
nor \U$44209 ( \44552 , \44549 , \44551 );
and \U$44210 ( \44553 , \44545 , \44552 );
and \U$44211 ( \44554 , \44539 , \44544 );
or \U$44212 ( \44555 , \44553 , \44554 );
xor \U$44213 ( \44556 , \44532 , \44555 );
and \U$44214 ( \44557 , \10424 , RI986df18_6);
and \U$44215 ( \44558 , RI986de28_4, \10422 );
nor \U$44216 ( \44559 , \44557 , \44558 );
and \U$44217 ( \44560 , \44559 , \9840 );
not \U$44218 ( \44561 , \44559 );
and \U$44219 ( \44562 , \44561 , \10428 );
nor \U$44220 ( \44563 , \44560 , \44562 );
and \U$44221 ( \44564 , \9237 , RI986f3b8_50);
and \U$44222 ( \44565 , RI986f598_54, \9235 );
nor \U$44223 ( \44566 , \44564 , \44565 );
and \U$44224 ( \44567 , \44566 , \9241 );
not \U$44225 ( \44568 , \44566 );
and \U$44226 ( \44569 , \44568 , \8836 );
nor \U$44227 ( \44570 , \44567 , \44569 );
xor \U$44228 ( \44571 , \44563 , \44570 );
and \U$44229 ( \44572 , \9505 , RI986f688_56);
and \U$44230 ( \44573 , RI986e008_8, \9503 );
nor \U$44231 ( \44574 , \44572 , \44573 );
and \U$44232 ( \44575 , \44574 , \9510 );
not \U$44233 ( \44576 , \44574 );
and \U$44234 ( \44577 , \44576 , \9513 );
nor \U$44235 ( \44578 , \44575 , \44577 );
and \U$44236 ( \44579 , \44571 , \44578 );
and \U$44237 ( \44580 , \44563 , \44570 );
or \U$44238 ( \44581 , \44579 , \44580 );
and \U$44239 ( \44582 , \44556 , \44581 );
and \U$44240 ( \44583 , \44532 , \44555 );
or \U$44241 ( \44584 , \44582 , \44583 );
xor \U$44242 ( \44585 , \44507 , \44584 );
and \U$44243 ( \44586 , \6453 , RI986e4b8_18);
and \U$44244 ( \44587 , RI986e788_24, \6451 );
nor \U$44245 ( \44588 , \44586 , \44587 );
and \U$44246 ( \44589 , \44588 , \6190 );
not \U$44247 ( \44590 , \44588 );
and \U$44248 ( \44591 , \44590 , \6705 );
nor \U$44249 ( \44592 , \44589 , \44591 );
and \U$44250 ( \44593 , \5318 , RI986eff8_42);
and \U$44251 ( \44594 , RI986f2c8_48, \5316 );
nor \U$44252 ( \44595 , \44593 , \44594 );
and \U$44253 ( \44596 , \44595 , \5052 );
not \U$44254 ( \44597 , \44595 );
and \U$44255 ( \44598 , \44597 , \5322 );
nor \U$44256 ( \44599 , \44596 , \44598 );
xor \U$44257 ( \44600 , \44592 , \44599 );
and \U$44258 ( \44601 , \5881 , RI986f1d8_46);
and \U$44259 ( \44602 , RI986e5a8_20, \5879 );
nor \U$44260 ( \44603 , \44601 , \44602 );
and \U$44261 ( \44604 , \44603 , \5594 );
not \U$44262 ( \44605 , \44603 );
and \U$44263 ( \44606 , \44605 , \5885 );
nor \U$44264 ( \44607 , \44604 , \44606 );
and \U$44265 ( \44608 , \44600 , \44607 );
and \U$44266 ( \44609 , \44592 , \44599 );
or \U$44267 ( \44610 , \44608 , \44609 );
and \U$44268 ( \44611 , \2464 , RI9871668_124);
and \U$44269 ( \44612 , RI986eb48_32, \2462 );
nor \U$44270 ( \44613 , \44611 , \44612 );
and \U$44271 ( \44614 , \44613 , \2468 );
not \U$44272 ( \44615 , \44613 );
and \U$44273 ( \44616 , \44615 , \2263 );
nor \U$44274 ( \44617 , \44614 , \44616 );
and \U$44275 ( \44618 , \2274 , RI9871848_128);
and \U$44276 ( \44619 , RI9871578_122, \2272 );
nor \U$44277 ( \44620 , \44618 , \44619 );
and \U$44278 ( \44621 , \44620 , \2030 );
not \U$44279 ( \44622 , \44620 );
and \U$44280 ( \44623 , \44622 , \2031 );
nor \U$44281 ( \44624 , \44621 , \44623 );
xor \U$44282 ( \44625 , \44617 , \44624 );
not \U$44283 ( \44626 , \3406 );
and \U$44284 ( \44627 , \3254 , RI986ea58_30);
and \U$44285 ( \44628 , RI986e968_28, \3252 );
nor \U$44286 ( \44629 , \44627 , \44628 );
not \U$44287 ( \44630 , \44629 );
or \U$44288 ( \44631 , \44626 , \44630 );
or \U$44289 ( \44632 , \44629 , \3406 );
nand \U$44290 ( \44633 , \44631 , \44632 );
and \U$44291 ( \44634 , \44625 , \44633 );
and \U$44292 ( \44635 , \44617 , \44624 );
or \U$44293 ( \44636 , \44634 , \44635 );
xor \U$44294 ( \44637 , \44610 , \44636 );
not \U$44295 ( \44638 , \3412 );
and \U$44296 ( \44639 , \3683 , RI986e878_26);
and \U$44297 ( \44640 , RI986ef08_40, \3681 );
nor \U$44298 ( \44641 , \44639 , \44640 );
not \U$44299 ( \44642 , \44641 );
or \U$44300 ( \44643 , \44638 , \44642 );
or \U$44301 ( \44644 , \44641 , \3412 );
nand \U$44302 ( \44645 , \44643 , \44644 );
and \U$44303 ( \44646 , \4203 , RI986ee18_38);
and \U$44304 ( \44647 , RI986ec38_34, \4201 );
nor \U$44305 ( \44648 , \44646 , \44647 );
and \U$44306 ( \44649 , \44648 , \4207 );
not \U$44307 ( \44650 , \44648 );
and \U$44308 ( \44651 , \44650 , \3922 );
nor \U$44309 ( \44652 , \44649 , \44651 );
xor \U$44310 ( \44653 , \44645 , \44652 );
not \U$44311 ( \44654 , \4521 );
and \U$44312 ( \44655 , \4710 , RI986ed28_36);
and \U$44313 ( \44656 , RI986f0e8_44, \4708 );
nor \U$44314 ( \44657 , \44655 , \44656 );
not \U$44315 ( \44658 , \44657 );
or \U$44316 ( \44659 , \44654 , \44658 );
or \U$44317 ( \44660 , \44657 , \4521 );
nand \U$44318 ( \44661 , \44659 , \44660 );
and \U$44319 ( \44662 , \44653 , \44661 );
and \U$44320 ( \44663 , \44645 , \44652 );
or \U$44321 ( \44664 , \44662 , \44663 );
and \U$44322 ( \44665 , \44637 , \44664 );
and \U$44323 ( \44666 , \44610 , \44636 );
or \U$44324 ( \44667 , \44665 , \44666 );
and \U$44325 ( \44668 , \44585 , \44667 );
and \U$44326 ( \44669 , \44507 , \44584 );
or \U$44327 ( \44670 , \44668 , \44669 );
xor \U$44328 ( \44671 , \44423 , \44670 );
xor \U$44329 ( \44672 , \44276 , \44283 );
xor \U$44330 ( \44673 , \44672 , \44292 );
xor \U$44331 ( \44674 , \44148 , \44155 );
xor \U$44332 ( \44675 , \44674 , \44163 );
xor \U$44333 ( \44676 , \44673 , \44675 );
xor \U$44334 ( \44677 , \44092 , \44099 );
xor \U$44335 ( \44678 , \44677 , \44108 );
and \U$44336 ( \44679 , \44676 , \44678 );
and \U$44337 ( \44680 , \44673 , \44675 );
or \U$44338 ( \44681 , \44679 , \44680 );
and \U$44339 ( \44682 , \416 , RI9870858_94);
and \U$44340 ( \44683 , RI986fb38_66, \414 );
nor \U$44341 ( \44684 , \44682 , \44683 );
and \U$44342 ( \44685 , \44684 , \421 );
not \U$44343 ( \44686 , \44684 );
and \U$44344 ( \44687 , \44686 , \422 );
nor \U$44345 ( \44688 , \44685 , \44687 );
nand \U$44346 ( \44689 , RI9870948_96, RI9871fc8_144);
or \U$44347 ( \44690 , \44688 , \44689 );
not \U$44348 ( \44691 , \44689 );
not \U$44349 ( \44692 , \44688 );
or \U$44350 ( \44693 , \44691 , \44692 );
not \U$44351 ( \44694 , \361 );
and \U$44352 ( \44695 , \354 , RI986fc28_68);
and \U$44353 ( \44696 , RI986fe08_72, \352 );
nor \U$44354 ( \44697 , \44695 , \44696 );
not \U$44355 ( \44698 , \44697 );
or \U$44356 ( \44699 , \44694 , \44698 );
or \U$44357 ( \44700 , \44697 , \345 );
nand \U$44358 ( \44701 , \44699 , \44700 );
nand \U$44359 ( \44702 , \44693 , \44701 );
nand \U$44360 ( \44703 , \44690 , \44702 );
xor \U$44361 ( \44704 , \44119 , \44127 );
xor \U$44362 ( \44705 , \44704 , \44136 );
and \U$44363 ( \44706 , \44703 , \44705 );
xor \U$44364 ( \44707 , \44048 , \44050 );
xor \U$44365 ( \44708 , \44707 , \44058 );
xor \U$44366 ( \44709 , \44119 , \44127 );
xor \U$44367 ( \44710 , \44709 , \44136 );
and \U$44368 ( \44711 , \44708 , \44710 );
and \U$44369 ( \44712 , \44703 , \44708 );
or \U$44370 ( \44713 , \44706 , \44711 , \44712 );
xor \U$44371 ( \44714 , \44681 , \44713 );
xor \U$44372 ( \44715 , \44250 , \44257 );
xor \U$44373 ( \44716 , \44715 , \44266 );
xor \U$44374 ( \44717 , \44220 , \44227 );
xor \U$44375 ( \44718 , \44717 , \44235 );
and \U$44376 ( \44719 , \44716 , \44718 );
xor \U$44377 ( \44720 , \44303 , \44310 );
xor \U$44378 ( \44721 , \44720 , \44318 );
xor \U$44379 ( \44722 , \44220 , \44227 );
xor \U$44380 ( \44723 , \44722 , \44235 );
and \U$44381 ( \44724 , \44721 , \44723 );
and \U$44382 ( \44725 , \44716 , \44721 );
or \U$44383 ( \44726 , \44719 , \44724 , \44725 );
and \U$44384 ( \44727 , \44714 , \44726 );
and \U$44385 ( \44728 , \44681 , \44713 );
or \U$44386 ( \44729 , \44727 , \44728 );
and \U$44387 ( \44730 , \44671 , \44729 );
and \U$44388 ( \44731 , \44423 , \44670 );
or \U$44389 ( \44732 , \44730 , \44731 );
xor \U$44390 ( \44733 , \44411 , \44732 );
xor \U$44391 ( \44734 , \44111 , \44139 );
xor \U$44392 ( \44735 , \44734 , \44166 );
xor \U$44393 ( \44736 , \44032 , \44034 );
xor \U$44394 ( \44737 , \44736 , \44037 );
and \U$44395 ( \44738 , \44735 , \44737 );
xor \U$44396 ( \44739 , \44061 , \44063 );
xor \U$44397 ( \44740 , \44739 , \44066 );
xor \U$44398 ( \44741 , \44032 , \44034 );
xor \U$44399 ( \44742 , \44741 , \44037 );
and \U$44400 ( \44743 , \44740 , \44742 );
and \U$44401 ( \44744 , \44735 , \44740 );
or \U$44402 ( \44745 , \44738 , \44743 , \44744 );
xor \U$44403 ( \44746 , \43742 , \43765 );
xor \U$44404 ( \44747 , \44746 , \43791 );
xor \U$44405 ( \44748 , \44745 , \44747 );
xor \U$44406 ( \44749 , \43659 , \43687 );
xor \U$44407 ( \44750 , \44749 , \43714 );
xor \U$44408 ( \44751 , \44350 , \44355 );
xor \U$44409 ( \44752 , \44750 , \44751 );
and \U$44410 ( \44753 , \44748 , \44752 );
and \U$44411 ( \44754 , \44745 , \44747 );
or \U$44412 ( \44755 , \44753 , \44754 );
and \U$44413 ( \44756 , \44733 , \44755 );
and \U$44414 ( \44757 , \44411 , \44732 );
or \U$44415 ( \44758 , \44756 , \44757 );
xor \U$44416 ( \44759 , \43881 , \43903 );
xor \U$44417 ( \44760 , \44759 , \43952 );
xor \U$44418 ( \44761 , \44758 , \44760 );
xor \U$44419 ( \44762 , \44085 , \44327 );
xor \U$44420 ( \44763 , \44762 , \44344 );
xor \U$44421 ( \44764 , \44020 , \44022 );
xor \U$44422 ( \44765 , \44764 , \44027 );
and \U$44423 ( \44766 , \44763 , \44765 );
xor \U$44424 ( \44767 , \43605 , \43607 );
xor \U$44425 ( \44768 , \44767 , \43610 );
xor \U$44426 ( \44769 , \44360 , \44367 );
xor \U$44427 ( \44770 , \44768 , \44769 );
xor \U$44428 ( \44771 , \44020 , \44022 );
xor \U$44429 ( \44772 , \44771 , \44027 );
and \U$44430 ( \44773 , \44770 , \44772 );
and \U$44431 ( \44774 , \44763 , \44770 );
or \U$44432 ( \44775 , \44766 , \44773 , \44774 );
and \U$44433 ( \44776 , \44761 , \44775 );
and \U$44434 ( \44777 , \44758 , \44760 );
or \U$44435 ( \44778 , \44776 , \44777 );
xor \U$44436 ( \44779 , \43633 , \43955 );
xor \U$44437 ( \44780 , \44779 , \43972 );
xor \U$44438 ( \44781 , \44778 , \44780 );
xor \U$44439 ( \44782 , \44030 , \44347 );
xor \U$44440 ( \44783 , \44782 , \44372 );
xor \U$44441 ( \44784 , \43613 , \43615 );
xor \U$44442 ( \44785 , \44784 , \43630 );
xor \U$44443 ( \44786 , \44006 , \44013 );
xor \U$44444 ( \44787 , \44785 , \44786 );
and \U$44445 ( \44788 , \44783 , \44787 );
xor \U$44446 ( \44789 , \44781 , \44788 );
and \U$44447 ( \44790 , \44397 , \44789 );
xor \U$44448 ( \44791 , \44423 , \44670 );
xor \U$44449 ( \44792 , \44791 , \44729 );
xor \U$44450 ( \44793 , \44745 , \44747 );
xor \U$44451 ( \44794 , \44793 , \44752 );
and \U$44452 ( \44795 , \44792 , \44794 );
xor \U$44453 ( \44796 , \44040 , \44069 );
xor \U$44454 ( \44797 , \44796 , \44082 );
xor \U$44455 ( \44798 , \44399 , \44406 );
xor \U$44456 ( \44799 , \44797 , \44798 );
xor \U$44457 ( \44800 , \44745 , \44747 );
xor \U$44458 ( \44801 , \44800 , \44752 );
and \U$44459 ( \44802 , \44799 , \44801 );
and \U$44460 ( \44803 , \44792 , \44799 );
or \U$44461 ( \44804 , \44795 , \44802 , \44803 );
xor \U$44462 ( \44805 , \44194 , \44212 );
xor \U$44463 ( \44806 , \44805 , \44238 );
xor \U$44464 ( \44807 , \44413 , \44415 );
xor \U$44465 ( \44808 , \44807 , \44420 );
and \U$44466 ( \44809 , \44806 , \44808 );
xor \U$44467 ( \44810 , \44032 , \44034 );
xor \U$44468 ( \44811 , \44810 , \44037 );
xor \U$44469 ( \44812 , \44735 , \44740 );
xor \U$44470 ( \44813 , \44811 , \44812 );
xor \U$44471 ( \44814 , \44413 , \44415 );
xor \U$44472 ( \44815 , \44814 , \44420 );
and \U$44473 ( \44816 , \44813 , \44815 );
and \U$44474 ( \44817 , \44806 , \44813 );
or \U$44475 ( \44818 , \44809 , \44816 , \44817 );
and \U$44476 ( \44819 , \1329 , RI98710c8_112);
and \U$44477 ( \44820 , RI9870d08_104, \1327 );
nor \U$44478 ( \44821 , \44819 , \44820 );
and \U$44479 ( \44822 , \44821 , \1336 );
not \U$44480 ( \44823 , \44821 );
and \U$44481 ( \44824 , \44823 , \1337 );
nor \U$44482 ( \44825 , \44822 , \44824 );
and \U$44483 ( \44826 , \776 , RI9870df8_106);
and \U$44484 ( \44827 , RI9870a38_98, \774 );
nor \U$44485 ( \44828 , \44826 , \44827 );
and \U$44486 ( \44829 , \44828 , \474 );
not \U$44487 ( \44830 , \44828 );
and \U$44488 ( \44831 , \44830 , \451 );
nor \U$44489 ( \44832 , \44829 , \44831 );
xor \U$44490 ( \44833 , \44825 , \44832 );
not \U$44491 ( \44834 , \1301 );
and \U$44492 ( \44835 , \1293 , RI9870ee8_108);
and \U$44493 ( \44836 , RI9870c18_102, \1291 );
nor \U$44494 ( \44837 , \44835 , \44836 );
not \U$44495 ( \44838 , \44837 );
or \U$44496 ( \44839 , \44834 , \44838 );
or \U$44497 ( \44840 , \44837 , \1128 );
nand \U$44498 ( \44841 , \44839 , \44840 );
and \U$44499 ( \44842 , \44833 , \44841 );
and \U$44500 ( \44843 , \44825 , \44832 );
or \U$44501 ( \44844 , \44842 , \44843 );
and \U$44502 ( \44845 , \438 , RI9870fd8_110);
and \U$44503 ( \44846 , RI9870b28_100, \436 );
nor \U$44504 ( \44847 , \44845 , \44846 );
and \U$44505 ( \44848 , \44847 , \444 );
not \U$44506 ( \44849 , \44847 );
and \U$44507 ( \44850 , \44849 , \443 );
nor \U$44508 ( \44851 , \44848 , \44850 );
not \U$44509 ( \44852 , \456 );
and \U$44510 ( \44853 , \465 , RI98700d8_78);
and \U$44511 ( \44854 , RI98701c8_80, \463 );
nor \U$44512 ( \44855 , \44853 , \44854 );
not \U$44513 ( \44856 , \44855 );
or \U$44514 ( \44857 , \44852 , \44856 );
or \U$44515 ( \44858 , \44855 , \454 );
nand \U$44516 ( \44859 , \44857 , \44858 );
xor \U$44517 ( \44860 , \44851 , \44859 );
not \U$44518 ( \44861 , \365 );
and \U$44519 ( \44862 , \376 , RI986ffe8_76);
and \U$44520 ( \44863 , RI986fef8_74, \374 );
nor \U$44521 ( \44864 , \44862 , \44863 );
not \U$44522 ( \44865 , \44864 );
or \U$44523 ( \44866 , \44861 , \44865 );
or \U$44524 ( \44867 , \44864 , \365 );
nand \U$44525 ( \44868 , \44866 , \44867 );
and \U$44526 ( \44869 , \44860 , \44868 );
and \U$44527 ( \44870 , \44851 , \44859 );
or \U$44528 ( \44871 , \44869 , \44870 );
xor \U$44529 ( \44872 , \44844 , \44871 );
and \U$44530 ( \44873 , \2274 , RI9871758_126);
and \U$44531 ( \44874 , RI9871848_128, \2272 );
nor \U$44532 ( \44875 , \44873 , \44874 );
and \U$44533 ( \44876 , \44875 , \2030 );
not \U$44534 ( \44877 , \44875 );
and \U$44535 ( \44878 , \44877 , \2031 );
nor \U$44536 ( \44879 , \44876 , \44878 );
and \U$44537 ( \44880 , \1311 , RI98712a8_116);
and \U$44538 ( \44881 , RI98711b8_114, \1309 );
nor \U$44539 ( \44882 , \44880 , \44881 );
and \U$44540 ( \44883 , \44882 , \1458 );
not \U$44541 ( \44884 , \44882 );
and \U$44542 ( \44885 , \44884 , \1318 );
nor \U$44543 ( \44886 , \44883 , \44885 );
xor \U$44544 ( \44887 , \44879 , \44886 );
not \U$44545 ( \44888 , \1462 );
and \U$44546 ( \44889 , \2042 , RI9871398_118);
and \U$44547 ( \44890 , RI9871488_120, \2040 );
nor \U$44548 ( \44891 , \44889 , \44890 );
not \U$44549 ( \44892 , \44891 );
or \U$44550 ( \44893 , \44888 , \44892 );
or \U$44551 ( \44894 , \44891 , \1462 );
nand \U$44552 ( \44895 , \44893 , \44894 );
and \U$44553 ( \44896 , \44887 , \44895 );
and \U$44554 ( \44897 , \44879 , \44886 );
or \U$44555 ( \44898 , \44896 , \44897 );
and \U$44556 ( \44899 , \44872 , \44898 );
and \U$44557 ( \44900 , \44844 , \44871 );
or \U$44558 ( \44901 , \44899 , \44900 );
and \U$44559 ( \44902 , \8486 , RI986fa48_64);
and \U$44560 ( \44903 , RI986f958_62, \8484 );
nor \U$44561 ( \44904 , \44902 , \44903 );
and \U$44562 ( \44905 , \44904 , \8050 );
not \U$44563 ( \44906 , \44904 );
and \U$44564 ( \44907 , \44906 , \8051 );
nor \U$44565 ( \44908 , \44905 , \44907 );
and \U$44566 ( \44909 , \7729 , RI986f868_60);
and \U$44567 ( \44910 , RI986f778_58, \7727 );
nor \U$44568 ( \44911 , \44909 , \44910 );
and \U$44569 ( \44912 , \44911 , \7480 );
not \U$44570 ( \44913 , \44911 );
and \U$44571 ( \44914 , \44913 , \7733 );
nor \U$44572 ( \44915 , \44912 , \44914 );
xor \U$44573 ( \44916 , \44908 , \44915 );
and \U$44574 ( \44917 , \9237 , RI986f4a8_52);
and \U$44575 ( \44918 , RI986f3b8_50, \9235 );
nor \U$44576 ( \44919 , \44917 , \44918 );
and \U$44577 ( \44920 , \44919 , \9241 );
not \U$44578 ( \44921 , \44919 );
and \U$44579 ( \44922 , \44921 , \8836 );
nor \U$44580 ( \44923 , \44920 , \44922 );
and \U$44581 ( \44924 , \44916 , \44923 );
and \U$44582 ( \44925 , \44908 , \44915 );
or \U$44583 ( \44926 , \44924 , \44925 );
and \U$44584 ( \44927 , \12293 , RI986e1e8_12);
and \U$44585 ( \44928 , RI986e0f8_10, \12291 );
nor \U$44586 ( \44929 , \44927 , \44928 );
and \U$44587 ( \44930 , \44929 , \11687 );
not \U$44588 ( \44931 , \44929 );
and \U$44589 ( \44932 , \44931 , \11686 );
nor \U$44590 ( \44933 , \44930 , \44932 );
xor \U$44591 ( \44934 , \44933 , \13358 );
and \U$44592 ( \44935 , \13045 , RI986e2d8_14);
and \U$44593 ( \44936 , RI986e3c8_16, \13043 );
nor \U$44594 ( \44937 , \44935 , \44936 );
and \U$44595 ( \44938 , \44937 , \13047 );
not \U$44596 ( \44939 , \44937 );
and \U$44597 ( \44940 , \44939 , \12619 );
nor \U$44598 ( \44941 , \44938 , \44940 );
and \U$44599 ( \44942 , \44934 , \44941 );
and \U$44600 ( \44943 , \44933 , \13358 );
or \U$44601 ( \44944 , \44942 , \44943 );
xor \U$44602 ( \44945 , \44926 , \44944 );
and \U$44603 ( \44946 , \11696 , RI986de28_4);
and \U$44604 ( \44947 , RI986dd38_2, \11694 );
nor \U$44605 ( \44948 , \44946 , \44947 );
and \U$44606 ( \44949 , \44948 , \10965 );
not \U$44607 ( \44950 , \44948 );
and \U$44608 ( \44951 , \44950 , \11702 );
nor \U$44609 ( \44952 , \44949 , \44951 );
and \U$44610 ( \44953 , \9505 , RI986f598_54);
and \U$44611 ( \44954 , RI986f688_56, \9503 );
nor \U$44612 ( \44955 , \44953 , \44954 );
and \U$44613 ( \44956 , \44955 , \9510 );
not \U$44614 ( \44957 , \44955 );
and \U$44615 ( \44958 , \44957 , \9513 );
nor \U$44616 ( \44959 , \44956 , \44958 );
xor \U$44617 ( \44960 , \44952 , \44959 );
and \U$44618 ( \44961 , \10424 , RI986e008_8);
and \U$44619 ( \44962 , RI986df18_6, \10422 );
nor \U$44620 ( \44963 , \44961 , \44962 );
and \U$44621 ( \44964 , \44963 , \9840 );
not \U$44622 ( \44965 , \44963 );
and \U$44623 ( \44966 , \44965 , \10428 );
nor \U$44624 ( \44967 , \44964 , \44966 );
and \U$44625 ( \44968 , \44960 , \44967 );
and \U$44626 ( \44969 , \44952 , \44959 );
or \U$44627 ( \44970 , \44968 , \44969 );
and \U$44628 ( \44971 , \44945 , \44970 );
and \U$44629 ( \44972 , \44926 , \44944 );
or \U$44630 ( \44973 , \44971 , \44972 );
xor \U$44631 ( \44974 , \44901 , \44973 );
and \U$44632 ( \44975 , \5318 , RI986f0e8_44);
and \U$44633 ( \44976 , RI986eff8_42, \5316 );
nor \U$44634 ( \44977 , \44975 , \44976 );
and \U$44635 ( \44978 , \44977 , \5052 );
not \U$44636 ( \44979 , \44977 );
and \U$44637 ( \44980 , \44979 , \5322 );
nor \U$44638 ( \44981 , \44978 , \44980 );
and \U$44639 ( \44982 , \4203 , RI986ef08_40);
and \U$44640 ( \44983 , RI986ee18_38, \4201 );
nor \U$44641 ( \44984 , \44982 , \44983 );
and \U$44642 ( \44985 , \44984 , \4207 );
not \U$44643 ( \44986 , \44984 );
and \U$44644 ( \44987 , \44986 , \3922 );
nor \U$44645 ( \44988 , \44985 , \44987 );
xor \U$44646 ( \44989 , \44981 , \44988 );
not \U$44647 ( \44990 , \4521 );
and \U$44648 ( \44991 , \4710 , RI986ec38_34);
and \U$44649 ( \44992 , RI986ed28_36, \4708 );
nor \U$44650 ( \44993 , \44991 , \44992 );
not \U$44651 ( \44994 , \44993 );
or \U$44652 ( \44995 , \44990 , \44994 );
or \U$44653 ( \44996 , \44993 , \4519 );
nand \U$44654 ( \44997 , \44995 , \44996 );
and \U$44655 ( \44998 , \44989 , \44997 );
and \U$44656 ( \44999 , \44981 , \44988 );
or \U$44657 ( \45000 , \44998 , \44999 );
not \U$44658 ( \45001 , \3918 );
and \U$44659 ( \45002 , \3683 , RI986e968_28);
and \U$44660 ( \45003 , RI986e878_26, \3681 );
nor \U$44661 ( \45004 , \45002 , \45003 );
not \U$44662 ( \45005 , \45004 );
or \U$44663 ( \45006 , \45001 , \45005 );
or \U$44664 ( \45007 , \45004 , \3918 );
nand \U$44665 ( \45008 , \45006 , \45007 );
and \U$44666 ( \45009 , \2464 , RI9871578_122);
and \U$44667 ( \45010 , RI9871668_124, \2462 );
nor \U$44668 ( \45011 , \45009 , \45010 );
and \U$44669 ( \45012 , \45011 , \2468 );
not \U$44670 ( \45013 , \45011 );
and \U$44671 ( \45014 , \45013 , \2263 );
nor \U$44672 ( \45015 , \45012 , \45014 );
xor \U$44673 ( \45016 , \45008 , \45015 );
not \U$44674 ( \45017 , \2935 );
and \U$44675 ( \45018 , \3254 , RI986eb48_32);
and \U$44676 ( \45019 , RI986ea58_30, \3252 );
nor \U$44677 ( \45020 , \45018 , \45019 );
not \U$44678 ( \45021 , \45020 );
or \U$44679 ( \45022 , \45017 , \45021 );
or \U$44680 ( \45023 , \45020 , \3406 );
nand \U$44681 ( \45024 , \45022 , \45023 );
and \U$44682 ( \45025 , \45016 , \45024 );
and \U$44683 ( \45026 , \45008 , \45015 );
or \U$44684 ( \45027 , \45025 , \45026 );
xor \U$44685 ( \45028 , \45000 , \45027 );
and \U$44686 ( \45029 , \7079 , RI986e788_24);
and \U$44687 ( \45030 , RI986e698_22, \7077 );
nor \U$44688 ( \45031 , \45029 , \45030 );
and \U$44689 ( \45032 , \45031 , \6710 );
not \U$44690 ( \45033 , \45031 );
and \U$44691 ( \45034 , \45033 , \6709 );
nor \U$44692 ( \45035 , \45032 , \45034 );
and \U$44693 ( \45036 , \5881 , RI986f2c8_48);
and \U$44694 ( \45037 , RI986f1d8_46, \5879 );
nor \U$44695 ( \45038 , \45036 , \45037 );
and \U$44696 ( \45039 , \45038 , \5594 );
not \U$44697 ( \45040 , \45038 );
and \U$44698 ( \45041 , \45040 , \5885 );
nor \U$44699 ( \45042 , \45039 , \45041 );
xor \U$44700 ( \45043 , \45035 , \45042 );
and \U$44701 ( \45044 , \6453 , RI986e5a8_20);
and \U$44702 ( \45045 , RI986e4b8_18, \6451 );
nor \U$44703 ( \45046 , \45044 , \45045 );
and \U$44704 ( \45047 , \45046 , \6190 );
not \U$44705 ( \45048 , \45046 );
and \U$44706 ( \45049 , \45048 , \6705 );
nor \U$44707 ( \45050 , \45047 , \45049 );
and \U$44708 ( \45051 , \45043 , \45050 );
and \U$44709 ( \45052 , \45035 , \45042 );
or \U$44710 ( \45053 , \45051 , \45052 );
and \U$44711 ( \45054 , \45028 , \45053 );
and \U$44712 ( \45055 , \45000 , \45027 );
or \U$44713 ( \45056 , \45054 , \45055 );
and \U$44714 ( \45057 , \44974 , \45056 );
and \U$44715 ( \45058 , \44901 , \44973 );
or \U$44716 ( \45059 , \45057 , \45058 );
xor \U$44717 ( \45060 , \44201 , \13047 );
xor \U$44718 ( \45061 , \45060 , \44209 );
xor \U$44719 ( \45062 , \44176 , \44183 );
xor \U$44720 ( \45063 , \45062 , \44191 );
and \U$44721 ( \45064 , \45061 , \45063 );
xor \U$44722 ( \45065 , \44563 , \44570 );
xor \U$44723 ( \45066 , \45065 , \44578 );
xor \U$44724 ( \45067 , \44539 , \44544 );
xor \U$44725 ( \45068 , \45067 , \44552 );
xor \U$44726 ( \45069 , \45066 , \45068 );
xor \U$44727 ( \45070 , \44514 , \44521 );
xor \U$44728 ( \45071 , \45070 , \44529 );
and \U$44729 ( \45072 , \45069 , \45071 );
and \U$44730 ( \45073 , \45066 , \45068 );
or \U$44731 ( \45074 , \45072 , \45073 );
xor \U$44732 ( \45075 , \44176 , \44183 );
xor \U$44733 ( \45076 , \45075 , \44191 );
and \U$44734 ( \45077 , \45074 , \45076 );
and \U$44735 ( \45078 , \45061 , \45074 );
or \U$44736 ( \45079 , \45064 , \45077 , \45078 );
xor \U$44737 ( \45080 , \45059 , \45079 );
xor \U$44738 ( \45081 , \44457 , \44465 );
xor \U$44739 ( \45082 , \45081 , \44474 );
xor \U$44740 ( \45083 , \44485 , \44492 );
xor \U$44741 ( \45084 , \45083 , \44501 );
and \U$44742 ( \45085 , \45082 , \45084 );
xor \U$44743 ( \45086 , \44431 , \44438 );
xor \U$44744 ( \45087 , \45086 , \44446 );
xor \U$44745 ( \45088 , \44485 , \44492 );
xor \U$44746 ( \45089 , \45088 , \44501 );
and \U$44747 ( \45090 , \45087 , \45089 );
and \U$44748 ( \45091 , \45082 , \45087 );
or \U$44749 ( \45092 , \45085 , \45090 , \45091 );
not \U$44750 ( \45093 , \487 );
and \U$44751 ( \45094 , \395 , RI986fe08_72);
and \U$44752 ( \45095 , RI986fd18_70, \393 );
nor \U$44753 ( \45096 , \45094 , \45095 );
not \U$44754 ( \45097 , \45096 );
or \U$44755 ( \45098 , \45093 , \45097 );
or \U$44756 ( \45099 , \45096 , \386 );
nand \U$44757 ( \45100 , \45098 , \45099 );
not \U$44758 ( \45101 , \361 );
and \U$44759 ( \45102 , \354 , RI986fb38_66);
and \U$44760 ( \45103 , RI986fc28_68, \352 );
nor \U$44761 ( \45104 , \45102 , \45103 );
not \U$44762 ( \45105 , \45104 );
or \U$44763 ( \45106 , \45101 , \45105 );
or \U$44764 ( \45107 , \45104 , \345 );
nand \U$44765 ( \45108 , \45106 , \45107 );
xor \U$44766 ( \45109 , \45100 , \45108 );
and \U$44767 ( \45110 , \416 , RI9870948_96);
and \U$44768 ( \45111 , RI9870858_94, \414 );
nor \U$44769 ( \45112 , \45110 , \45111 );
and \U$44770 ( \45113 , \45112 , \422 );
not \U$44771 ( \45114 , \45112 );
and \U$44772 ( \45115 , \45114 , \421 );
nor \U$44773 ( \45116 , \45113 , \45115 );
and \U$44774 ( \45117 , \45109 , \45116 );
and \U$44775 ( \45118 , \45100 , \45108 );
nor \U$44776 ( \45119 , \45117 , \45118 );
not \U$44777 ( \45120 , \44688 );
not \U$44778 ( \45121 , \44701 );
or \U$44779 ( \45122 , \45120 , \45121 );
or \U$44780 ( \45123 , \44688 , \44701 );
nand \U$44781 ( \45124 , \45122 , \45123 );
not \U$44782 ( \45125 , \45124 );
not \U$44783 ( \45126 , \44689 );
and \U$44784 ( \45127 , \45125 , \45126 );
and \U$44785 ( \45128 , \45124 , \44689 );
nor \U$44786 ( \45129 , \45127 , \45128 );
nand \U$44787 ( \45130 , \45119 , \45129 );
xor \U$44788 ( \45131 , \45092 , \45130 );
xor \U$44789 ( \45132 , \44645 , \44652 );
xor \U$44790 ( \45133 , \45132 , \44661 );
xor \U$44791 ( \45134 , \44617 , \44624 );
xor \U$44792 ( \45135 , \45134 , \44633 );
and \U$44793 ( \45136 , \45133 , \45135 );
xor \U$44794 ( \45137 , \44592 , \44599 );
xor \U$44795 ( \45138 , \45137 , \44607 );
xor \U$44796 ( \45139 , \44617 , \44624 );
xor \U$44797 ( \45140 , \45139 , \44633 );
and \U$44798 ( \45141 , \45138 , \45140 );
and \U$44799 ( \45142 , \45133 , \45138 );
or \U$44800 ( \45143 , \45136 , \45141 , \45142 );
and \U$44801 ( \45144 , \45131 , \45143 );
and \U$44802 ( \45145 , \45092 , \45130 );
or \U$44803 ( \45146 , \45144 , \45145 );
and \U$44804 ( \45147 , \45080 , \45146 );
and \U$44805 ( \45148 , \45059 , \45079 );
or \U$44806 ( \45149 , \45147 , \45148 );
xor \U$44807 ( \45150 , \44818 , \45149 );
xor \U$44808 ( \45151 , \44449 , \44477 );
xor \U$44809 ( \45152 , \45151 , \44504 );
xor \U$44810 ( \45153 , \44532 , \44555 );
xor \U$44811 ( \45154 , \45153 , \44581 );
xor \U$44812 ( \45155 , \45152 , \45154 );
xor \U$44813 ( \45156 , \44610 , \44636 );
xor \U$44814 ( \45157 , \45156 , \44664 );
and \U$44815 ( \45158 , \45155 , \45157 );
and \U$44816 ( \45159 , \45152 , \45154 );
or \U$44817 ( \45160 , \45158 , \45159 );
xor \U$44818 ( \45161 , \44269 , \44295 );
xor \U$44819 ( \45162 , \45161 , \44321 );
xor \U$44820 ( \45163 , \45160 , \45162 );
xor \U$44821 ( \45164 , \44119 , \44127 );
xor \U$44822 ( \45165 , \45164 , \44136 );
xor \U$44823 ( \45166 , \44703 , \44708 );
xor \U$44824 ( \45167 , \45165 , \45166 );
xor \U$44825 ( \45168 , \44673 , \44675 );
xor \U$44826 ( \45169 , \45168 , \44678 );
and \U$44827 ( \45170 , \45167 , \45169 );
xor \U$44828 ( \45171 , \44220 , \44227 );
xor \U$44829 ( \45172 , \45171 , \44235 );
xor \U$44830 ( \45173 , \44716 , \44721 );
xor \U$44831 ( \45174 , \45172 , \45173 );
xor \U$44832 ( \45175 , \44673 , \44675 );
xor \U$44833 ( \45176 , \45175 , \44678 );
and \U$44834 ( \45177 , \45174 , \45176 );
and \U$44835 ( \45178 , \45167 , \45174 );
or \U$44836 ( \45179 , \45170 , \45177 , \45178 );
and \U$44837 ( \45180 , \45163 , \45179 );
and \U$44838 ( \45181 , \45160 , \45162 );
or \U$44839 ( \45182 , \45180 , \45181 );
and \U$44840 ( \45183 , \45150 , \45182 );
and \U$44841 ( \45184 , \44818 , \45149 );
or \U$44842 ( \45185 , \45183 , \45184 );
xor \U$44843 ( \45186 , \44804 , \45185 );
xor \U$44844 ( \45187 , \44020 , \44022 );
xor \U$44845 ( \45188 , \45187 , \44027 );
xor \U$44846 ( \45189 , \44763 , \44770 );
xor \U$44847 ( \45190 , \45188 , \45189 );
and \U$44848 ( \45191 , \45186 , \45190 );
and \U$44849 ( \45192 , \44804 , \45185 );
or \U$44850 ( \45193 , \45191 , \45192 );
xor \U$44851 ( \45194 , \44783 , \44787 );
xor \U$44852 ( \45195 , \45193 , \45194 );
xor \U$44853 ( \45196 , \44758 , \44760 );
xor \U$44854 ( \45197 , \45196 , \44775 );
and \U$44855 ( \45198 , \45195 , \45197 );
and \U$44856 ( \45199 , \45193 , \45194 );
or \U$44857 ( \45200 , \45198 , \45199 );
xor \U$44858 ( \45201 , \44778 , \44780 );
xor \U$44859 ( \45202 , \45201 , \44788 );
and \U$44860 ( \45203 , \45200 , \45202 );
and \U$44861 ( \45204 , \44397 , \45200 );
or \U$44862 ( \45205 , \44790 , \45203 , \45204 );
not \U$44863 ( \45206 , \45205 );
xor \U$44864 ( \45207 , \44778 , \44780 );
and \U$44865 ( \45208 , \45207 , \44788 );
and \U$44866 ( \45209 , \44778 , \44780 );
or \U$44867 ( \45210 , \45208 , \45209 );
xor \U$44868 ( \45211 , \43603 , \43975 );
xor \U$44869 ( \45212 , \45211 , \43980 );
xor \U$44870 ( \45213 , \44001 , \44383 );
xor \U$44871 ( \45214 , \45212 , \45213 );
xor \U$44872 ( \45215 , \45210 , \45214 );
not \U$44873 ( \45216 , \45215 );
or \U$44874 ( \45217 , \45206 , \45216 );
xor \U$44875 ( \45218 , \44778 , \44780 );
xor \U$44876 ( \45219 , \45218 , \44788 );
xor \U$44877 ( \45220 , \44397 , \45200 );
xor \U$44878 ( \45221 , \45219 , \45220 );
xor \U$44879 ( \45222 , \44176 , \44183 );
xor \U$44880 ( \45223 , \45222 , \44191 );
xor \U$44881 ( \45224 , \45061 , \45074 );
xor \U$44882 ( \45225 , \45223 , \45224 );
xor \U$44883 ( \45226 , \44901 , \44973 );
xor \U$44884 ( \45227 , \45226 , \45056 );
xor \U$44885 ( \45228 , \45225 , \45227 );
xor \U$44886 ( \45229 , \45092 , \45130 );
xor \U$44887 ( \45230 , \45229 , \45143 );
and \U$44888 ( \45231 , \45228 , \45230 );
and \U$44889 ( \45232 , \45225 , \45227 );
or \U$44890 ( \45233 , \45231 , \45232 );
xor \U$44891 ( \45234 , \45100 , \45108 );
xor \U$44892 ( \45235 , \45234 , \45116 );
xor \U$44893 ( \45236 , \44851 , \44859 );
xor \U$44894 ( \45237 , \45236 , \44868 );
and \U$44895 ( \45238 , \45235 , \45237 );
xor \U$44896 ( \45239 , \44825 , \44832 );
xor \U$44897 ( \45240 , \45239 , \44841 );
xor \U$44898 ( \45241 , \44851 , \44859 );
xor \U$44899 ( \45242 , \45241 , \44868 );
and \U$44900 ( \45243 , \45240 , \45242 );
and \U$44901 ( \45244 , \45235 , \45240 );
or \U$44902 ( \45245 , \45238 , \45243 , \45244 );
nand \U$44903 ( \45246 , RI9870768_92, RI9871fc8_144);
not \U$44904 ( \45247 , \45246 );
not \U$44905 ( \45248 , RI9870678_90);
nor \U$44906 ( \45249 , \45248 , \407 );
xor \U$44907 ( \45250 , \45247 , \45249 );
not \U$44908 ( \45251 , \386 );
and \U$44909 ( \45252 , \395 , RI986fc28_68);
and \U$44910 ( \45253 , RI986fe08_72, \393 );
nor \U$44911 ( \45254 , \45252 , \45253 );
not \U$44912 ( \45255 , \45254 );
or \U$44913 ( \45256 , \45251 , \45255 );
or \U$44914 ( \45257 , \45254 , \386 );
nand \U$44915 ( \45258 , \45256 , \45257 );
not \U$44916 ( \45259 , \361 );
and \U$44917 ( \45260 , \354 , RI9870858_94);
and \U$44918 ( \45261 , RI986fb38_66, \352 );
nor \U$44919 ( \45262 , \45260 , \45261 );
not \U$44920 ( \45263 , \45262 );
or \U$44921 ( \45264 , \45259 , \45263 );
or \U$44922 ( \45265 , \45262 , \345 );
nand \U$44923 ( \45266 , \45264 , \45265 );
xor \U$44924 ( \45267 , \45258 , \45266 );
and \U$44925 ( \45268 , \416 , RI9870678_90);
and \U$44926 ( \45269 , RI9870948_96, \414 );
nor \U$44927 ( \45270 , \45268 , \45269 );
and \U$44928 ( \45271 , \45270 , \422 );
not \U$44929 ( \45272 , \45270 );
and \U$44930 ( \45273 , \45272 , \421 );
nor \U$44931 ( \45274 , \45271 , \45273 );
and \U$44932 ( \45275 , \45267 , \45274 );
and \U$44933 ( \45276 , \45258 , \45266 );
or \U$44934 ( \45277 , \45275 , \45276 );
and \U$44935 ( \45278 , \45250 , \45277 );
and \U$44936 ( \45279 , \45247 , \45249 );
or \U$44937 ( \45280 , \45278 , \45279 );
xor \U$44938 ( \45281 , \45245 , \45280 );
xor \U$44939 ( \45282 , \44981 , \44988 );
xor \U$44940 ( \45283 , \45282 , \44997 );
xor \U$44941 ( \45284 , \44879 , \44886 );
xor \U$44942 ( \45285 , \45284 , \44895 );
xor \U$44943 ( \45286 , \45283 , \45285 );
xor \U$44944 ( \45287 , \45008 , \45015 );
xor \U$44945 ( \45288 , \45287 , \45024 );
and \U$44946 ( \45289 , \45286 , \45288 );
and \U$44947 ( \45290 , \45283 , \45285 );
or \U$44948 ( \45291 , \45289 , \45290 );
and \U$44949 ( \45292 , \45281 , \45291 );
and \U$44950 ( \45293 , \45245 , \45280 );
or \U$44951 ( \45294 , \45292 , \45293 );
and \U$44952 ( \45295 , \7079 , RI986e4b8_18);
and \U$44953 ( \45296 , RI986e788_24, \7077 );
nor \U$44954 ( \45297 , \45295 , \45296 );
and \U$44955 ( \45298 , \45297 , \6710 );
not \U$44956 ( \45299 , \45297 );
and \U$44957 ( \45300 , \45299 , \6709 );
nor \U$44958 ( \45301 , \45298 , \45300 );
and \U$44959 ( \45302 , \5881 , RI986eff8_42);
and \U$44960 ( \45303 , RI986f2c8_48, \5879 );
nor \U$44961 ( \45304 , \45302 , \45303 );
and \U$44962 ( \45305 , \45304 , \5594 );
not \U$44963 ( \45306 , \45304 );
and \U$44964 ( \45307 , \45306 , \5885 );
nor \U$44965 ( \45308 , \45305 , \45307 );
xor \U$44966 ( \45309 , \45301 , \45308 );
and \U$44967 ( \45310 , \6453 , RI986f1d8_46);
and \U$44968 ( \45311 , RI986e5a8_20, \6451 );
nor \U$44969 ( \45312 , \45310 , \45311 );
and \U$44970 ( \45313 , \45312 , \6190 );
not \U$44971 ( \45314 , \45312 );
and \U$44972 ( \45315 , \45314 , \6180 );
nor \U$44973 ( \45316 , \45313 , \45315 );
and \U$44974 ( \45317 , \45309 , \45316 );
and \U$44975 ( \45318 , \45301 , \45308 );
or \U$44976 ( \45319 , \45317 , \45318 );
not \U$44977 ( \45320 , \2935 );
and \U$44978 ( \45321 , \3254 , RI9871668_124);
and \U$44979 ( \45322 , RI986eb48_32, \3252 );
nor \U$44980 ( \45323 , \45321 , \45322 );
not \U$44981 ( \45324 , \45323 );
or \U$44982 ( \45325 , \45320 , \45324 );
or \U$44983 ( \45326 , \45323 , \3406 );
nand \U$44984 ( \45327 , \45325 , \45326 );
and \U$44985 ( \45328 , \2464 , RI9871848_128);
and \U$44986 ( \45329 , RI9871578_122, \2462 );
nor \U$44987 ( \45330 , \45328 , \45329 );
and \U$44988 ( \45331 , \45330 , \2468 );
not \U$44989 ( \45332 , \45330 );
and \U$44990 ( \45333 , \45332 , \2263 );
nor \U$44991 ( \45334 , \45331 , \45333 );
xor \U$44992 ( \45335 , \45327 , \45334 );
not \U$44993 ( \45336 , \3918 );
and \U$44994 ( \45337 , \3683 , RI986ea58_30);
and \U$44995 ( \45338 , RI986e968_28, \3681 );
nor \U$44996 ( \45339 , \45337 , \45338 );
not \U$44997 ( \45340 , \45339 );
or \U$44998 ( \45341 , \45336 , \45340 );
or \U$44999 ( \45342 , \45339 , \3918 );
nand \U$45000 ( \45343 , \45341 , \45342 );
and \U$45001 ( \45344 , \45335 , \45343 );
and \U$45002 ( \45345 , \45327 , \45334 );
or \U$45003 ( \45346 , \45344 , \45345 );
xor \U$45004 ( \45347 , \45319 , \45346 );
not \U$45005 ( \45348 , \4519 );
and \U$45006 ( \45349 , \4710 , RI986ee18_38);
and \U$45007 ( \45350 , RI986ec38_34, \4708 );
nor \U$45008 ( \45351 , \45349 , \45350 );
not \U$45009 ( \45352 , \45351 );
or \U$45010 ( \45353 , \45348 , \45352 );
or \U$45011 ( \45354 , \45351 , \4519 );
nand \U$45012 ( \45355 , \45353 , \45354 );
and \U$45013 ( \45356 , \4203 , RI986e878_26);
and \U$45014 ( \45357 , RI986ef08_40, \4201 );
nor \U$45015 ( \45358 , \45356 , \45357 );
and \U$45016 ( \45359 , \45358 , \4207 );
not \U$45017 ( \45360 , \45358 );
and \U$45018 ( \45361 , \45360 , \3923 );
nor \U$45019 ( \45362 , \45359 , \45361 );
xor \U$45020 ( \45363 , \45355 , \45362 );
and \U$45021 ( \45364 , \5318 , RI986ed28_36);
and \U$45022 ( \45365 , RI986f0e8_44, \5316 );
nor \U$45023 ( \45366 , \45364 , \45365 );
and \U$45024 ( \45367 , \45366 , \5052 );
not \U$45025 ( \45368 , \45366 );
and \U$45026 ( \45369 , \45368 , \5322 );
nor \U$45027 ( \45370 , \45367 , \45369 );
and \U$45028 ( \45371 , \45363 , \45370 );
and \U$45029 ( \45372 , \45355 , \45362 );
or \U$45030 ( \45373 , \45371 , \45372 );
and \U$45031 ( \45374 , \45347 , \45373 );
and \U$45032 ( \45375 , \45319 , \45346 );
or \U$45033 ( \45376 , \45374 , \45375 );
and \U$45034 ( \45377 , \2274 , RI9871488_120);
and \U$45035 ( \45378 , RI9871758_126, \2272 );
nor \U$45036 ( \45379 , \45377 , \45378 );
and \U$45037 ( \45380 , \45379 , \2030 );
not \U$45038 ( \45381 , \45379 );
and \U$45039 ( \45382 , \45381 , \2031 );
nor \U$45040 ( \45383 , \45380 , \45382 );
and \U$45041 ( \45384 , \1311 , RI9870d08_104);
and \U$45042 ( \45385 , RI98712a8_116, \1309 );
nor \U$45043 ( \45386 , \45384 , \45385 );
and \U$45044 ( \45387 , \45386 , \1458 );
not \U$45045 ( \45388 , \45386 );
and \U$45046 ( \45389 , \45388 , \1315 );
nor \U$45047 ( \45390 , \45387 , \45389 );
xor \U$45048 ( \45391 , \45383 , \45390 );
not \U$45049 ( \45392 , \2034 );
and \U$45050 ( \45393 , \2042 , RI98711b8_114);
and \U$45051 ( \45394 , RI9871398_118, \2040 );
nor \U$45052 ( \45395 , \45393 , \45394 );
not \U$45053 ( \45396 , \45395 );
or \U$45054 ( \45397 , \45392 , \45396 );
or \U$45055 ( \45398 , \45395 , \1462 );
nand \U$45056 ( \45399 , \45397 , \45398 );
and \U$45057 ( \45400 , \45391 , \45399 );
and \U$45058 ( \45401 , \45383 , \45390 );
or \U$45059 ( \45402 , \45400 , \45401 );
and \U$45060 ( \45403 , \1329 , RI9870c18_102);
and \U$45061 ( \45404 , RI98710c8_112, \1327 );
nor \U$45062 ( \45405 , \45403 , \45404 );
and \U$45063 ( \45406 , \45405 , \1336 );
not \U$45064 ( \45407 , \45405 );
and \U$45065 ( \45408 , \45407 , \1337 );
nor \U$45066 ( \45409 , \45406 , \45408 );
and \U$45067 ( \45410 , \776 , RI9870b28_100);
and \U$45068 ( \45411 , RI9870df8_106, \774 );
nor \U$45069 ( \45412 , \45410 , \45411 );
and \U$45070 ( \45413 , \45412 , \474 );
not \U$45071 ( \45414 , \45412 );
and \U$45072 ( \45415 , \45414 , \451 );
nor \U$45073 ( \45416 , \45413 , \45415 );
xor \U$45074 ( \45417 , \45409 , \45416 );
not \U$45075 ( \45418 , \1301 );
and \U$45076 ( \45419 , \1293 , RI9870a38_98);
and \U$45077 ( \45420 , RI9870ee8_108, \1291 );
nor \U$45078 ( \45421 , \45419 , \45420 );
not \U$45079 ( \45422 , \45421 );
or \U$45080 ( \45423 , \45418 , \45422 );
or \U$45081 ( \45424 , \45421 , \1301 );
nand \U$45082 ( \45425 , \45423 , \45424 );
and \U$45083 ( \45426 , \45417 , \45425 );
and \U$45084 ( \45427 , \45409 , \45416 );
or \U$45085 ( \45428 , \45426 , \45427 );
xor \U$45086 ( \45429 , \45402 , \45428 );
not \U$45087 ( \45430 , \367 );
and \U$45088 ( \45431 , \376 , RI986fd18_70);
and \U$45089 ( \45432 , RI986ffe8_76, \374 );
nor \U$45090 ( \45433 , \45431 , \45432 );
not \U$45091 ( \45434 , \45433 );
or \U$45092 ( \45435 , \45430 , \45434 );
or \U$45093 ( \45436 , \45433 , \365 );
nand \U$45094 ( \45437 , \45435 , \45436 );
and \U$45095 ( \45438 , \438 , RI98701c8_80);
and \U$45096 ( \45439 , RI9870fd8_110, \436 );
nor \U$45097 ( \45440 , \45438 , \45439 );
and \U$45098 ( \45441 , \45440 , \444 );
not \U$45099 ( \45442 , \45440 );
and \U$45100 ( \45443 , \45442 , \443 );
nor \U$45101 ( \45444 , \45441 , \45443 );
xor \U$45102 ( \45445 , \45437 , \45444 );
not \U$45103 ( \45446 , \456 );
and \U$45104 ( \45447 , \465 , RI986fef8_74);
and \U$45105 ( \45448 , RI98700d8_78, \463 );
nor \U$45106 ( \45449 , \45447 , \45448 );
not \U$45107 ( \45450 , \45449 );
or \U$45108 ( \45451 , \45446 , \45450 );
or \U$45109 ( \45452 , \45449 , \456 );
nand \U$45110 ( \45453 , \45451 , \45452 );
and \U$45111 ( \45454 , \45445 , \45453 );
and \U$45112 ( \45455 , \45437 , \45444 );
or \U$45113 ( \45456 , \45454 , \45455 );
and \U$45114 ( \45457 , \45429 , \45456 );
and \U$45115 ( \45458 , \45402 , \45428 );
or \U$45116 ( \45459 , \45457 , \45458 );
xor \U$45117 ( \45460 , \45376 , \45459 );
and \U$45118 ( \45461 , \9237 , RI986f958_62);
and \U$45119 ( \45462 , RI986f4a8_52, \9235 );
nor \U$45120 ( \45463 , \45461 , \45462 );
and \U$45121 ( \45464 , \45463 , \9241 );
not \U$45122 ( \45465 , \45463 );
and \U$45123 ( \45466 , \45465 , \8836 );
nor \U$45124 ( \45467 , \45464 , \45466 );
and \U$45125 ( \45468 , \7729 , RI986e698_22);
and \U$45126 ( \45469 , RI986f868_60, \7727 );
nor \U$45127 ( \45470 , \45468 , \45469 );
and \U$45128 ( \45471 , \45470 , \7480 );
not \U$45129 ( \45472 , \45470 );
and \U$45130 ( \45473 , \45472 , \7733 );
nor \U$45131 ( \45474 , \45471 , \45473 );
xor \U$45132 ( \45475 , \45467 , \45474 );
and \U$45133 ( \45476 , \8486 , RI986f778_58);
and \U$45134 ( \45477 , RI986fa48_64, \8484 );
nor \U$45135 ( \45478 , \45476 , \45477 );
and \U$45136 ( \45479 , \45478 , \8050 );
not \U$45137 ( \45480 , \45478 );
and \U$45138 ( \45481 , \45480 , \8051 );
nor \U$45139 ( \45482 , \45479 , \45481 );
and \U$45140 ( \45483 , \45475 , \45482 );
and \U$45141 ( \45484 , \45467 , \45474 );
or \U$45142 ( \45485 , \45483 , \45484 );
and \U$45143 ( \45486 , \12293 , RI986dd38_2);
and \U$45144 ( \45487 , RI986e1e8_12, \12291 );
nor \U$45145 ( \45488 , \45486 , \45487 );
and \U$45146 ( \45489 , \45488 , \11687 );
not \U$45147 ( \45490 , \45488 );
and \U$45148 ( \45491 , \45490 , \11686 );
nor \U$45149 ( \45492 , \45489 , \45491 );
nand \U$45150 ( \45493 , RI986e3c8_16, \13882 );
and \U$45151 ( \45494 , \45493 , \13358 );
not \U$45152 ( \45495 , \45493 );
and \U$45153 ( \45496 , \45495 , \13359 );
nor \U$45154 ( \45497 , \45494 , \45496 );
xor \U$45155 ( \45498 , \45492 , \45497 );
and \U$45156 ( \45499 , \13045 , RI986e0f8_10);
and \U$45157 ( \45500 , RI986e2d8_14, \13043 );
nor \U$45158 ( \45501 , \45499 , \45500 );
and \U$45159 ( \45502 , \45501 , \13047 );
not \U$45160 ( \45503 , \45501 );
and \U$45161 ( \45504 , \45503 , \12619 );
nor \U$45162 ( \45505 , \45502 , \45504 );
and \U$45163 ( \45506 , \45498 , \45505 );
and \U$45164 ( \45507 , \45492 , \45497 );
or \U$45165 ( \45508 , \45506 , \45507 );
xor \U$45166 ( \45509 , \45485 , \45508 );
and \U$45167 ( \45510 , \11696 , RI986df18_6);
and \U$45168 ( \45511 , RI986de28_4, \11694 );
nor \U$45169 ( \45512 , \45510 , \45511 );
and \U$45170 ( \45513 , \45512 , \10965 );
not \U$45171 ( \45514 , \45512 );
and \U$45172 ( \45515 , \45514 , \11702 );
nor \U$45173 ( \45516 , \45513 , \45515 );
and \U$45174 ( \45517 , \9505 , RI986f3b8_50);
and \U$45175 ( \45518 , RI986f598_54, \9503 );
nor \U$45176 ( \45519 , \45517 , \45518 );
and \U$45177 ( \45520 , \45519 , \9510 );
not \U$45178 ( \45521 , \45519 );
and \U$45179 ( \45522 , \45521 , \9513 );
nor \U$45180 ( \45523 , \45520 , \45522 );
xor \U$45181 ( \45524 , \45516 , \45523 );
and \U$45182 ( \45525 , \10424 , RI986f688_56);
and \U$45183 ( \45526 , RI986e008_8, \10422 );
nor \U$45184 ( \45527 , \45525 , \45526 );
and \U$45185 ( \45528 , \45527 , \9840 );
not \U$45186 ( \45529 , \45527 );
and \U$45187 ( \45530 , \45529 , \10428 );
nor \U$45188 ( \45531 , \45528 , \45530 );
and \U$45189 ( \45532 , \45524 , \45531 );
and \U$45190 ( \45533 , \45516 , \45523 );
or \U$45191 ( \45534 , \45532 , \45533 );
and \U$45192 ( \45535 , \45509 , \45534 );
and \U$45193 ( \45536 , \45485 , \45508 );
or \U$45194 ( \45537 , \45535 , \45536 );
and \U$45195 ( \45538 , \45460 , \45537 );
and \U$45196 ( \45539 , \45376 , \45459 );
or \U$45197 ( \45540 , \45538 , \45539 );
xor \U$45198 ( \45541 , \45294 , \45540 );
xor \U$45199 ( \45542 , \45035 , \45042 );
xor \U$45200 ( \45543 , \45542 , \45050 );
xor \U$45201 ( \45544 , \44908 , \44915 );
xor \U$45202 ( \45545 , \45544 , \44923 );
and \U$45203 ( \45546 , \45543 , \45545 );
xor \U$45204 ( \45547 , \44952 , \44959 );
xor \U$45205 ( \45548 , \45547 , \44967 );
xor \U$45206 ( \45549 , \44908 , \44915 );
xor \U$45207 ( \45550 , \45549 , \44923 );
and \U$45208 ( \45551 , \45548 , \45550 );
and \U$45209 ( \45552 , \45543 , \45548 );
or \U$45210 ( \45553 , \45546 , \45551 , \45552 );
xor \U$45211 ( \45554 , \45066 , \45068 );
xor \U$45212 ( \45555 , \45554 , \45071 );
and \U$45213 ( \45556 , \45553 , \45555 );
xor \U$45214 ( \45557 , \44617 , \44624 );
xor \U$45215 ( \45558 , \45557 , \44633 );
xor \U$45216 ( \45559 , \45133 , \45138 );
xor \U$45217 ( \45560 , \45558 , \45559 );
xor \U$45218 ( \45561 , \45066 , \45068 );
xor \U$45219 ( \45562 , \45561 , \45071 );
and \U$45220 ( \45563 , \45560 , \45562 );
and \U$45221 ( \45564 , \45553 , \45560 );
or \U$45222 ( \45565 , \45556 , \45563 , \45564 );
and \U$45223 ( \45566 , \45541 , \45565 );
and \U$45224 ( \45567 , \45294 , \45540 );
or \U$45225 ( \45568 , \45566 , \45567 );
xor \U$45226 ( \45569 , \45233 , \45568 );
xor \U$45227 ( \45570 , \44844 , \44871 );
xor \U$45228 ( \45571 , \45570 , \44898 );
or \U$45229 ( \45572 , \45129 , \45119 );
nand \U$45230 ( \45573 , \45572 , \45130 );
xor \U$45231 ( \45574 , \45571 , \45573 );
xor \U$45232 ( \45575 , \44485 , \44492 );
xor \U$45233 ( \45576 , \45575 , \44501 );
xor \U$45234 ( \45577 , \45082 , \45087 );
xor \U$45235 ( \45578 , \45576 , \45577 );
and \U$45236 ( \45579 , \45574 , \45578 );
and \U$45237 ( \45580 , \45571 , \45573 );
or \U$45238 ( \45581 , \45579 , \45580 );
xor \U$45239 ( \45582 , \45152 , \45154 );
xor \U$45240 ( \45583 , \45582 , \45157 );
and \U$45241 ( \45584 , \45581 , \45583 );
xor \U$45242 ( \45585 , \44673 , \44675 );
xor \U$45243 ( \45586 , \45585 , \44678 );
xor \U$45244 ( \45587 , \45167 , \45174 );
xor \U$45245 ( \45588 , \45586 , \45587 );
xor \U$45246 ( \45589 , \45152 , \45154 );
xor \U$45247 ( \45590 , \45589 , \45157 );
and \U$45248 ( \45591 , \45588 , \45590 );
and \U$45249 ( \45592 , \45581 , \45588 );
or \U$45250 ( \45593 , \45584 , \45591 , \45592 );
and \U$45251 ( \45594 , \45569 , \45593 );
and \U$45252 ( \45595 , \45233 , \45568 );
or \U$45253 ( \45596 , \45594 , \45595 );
xor \U$45254 ( \45597 , \44681 , \44713 );
xor \U$45255 ( \45598 , \45597 , \44726 );
xor \U$45256 ( \45599 , \44507 , \44584 );
xor \U$45257 ( \45600 , \45599 , \44667 );
xor \U$45258 ( \45601 , \45598 , \45600 );
xor \U$45259 ( \45602 , \44413 , \44415 );
xor \U$45260 ( \45603 , \45602 , \44420 );
xor \U$45261 ( \45604 , \44806 , \44813 );
xor \U$45262 ( \45605 , \45603 , \45604 );
and \U$45263 ( \45606 , \45601 , \45605 );
and \U$45264 ( \45607 , \45598 , \45600 );
or \U$45265 ( \45608 , \45606 , \45607 );
xor \U$45266 ( \45609 , \45596 , \45608 );
xor \U$45267 ( \45610 , \44745 , \44747 );
xor \U$45268 ( \45611 , \45610 , \44752 );
xor \U$45269 ( \45612 , \44792 , \44799 );
xor \U$45270 ( \45613 , \45611 , \45612 );
and \U$45271 ( \45614 , \45609 , \45613 );
and \U$45272 ( \45615 , \45596 , \45608 );
or \U$45273 ( \45616 , \45614 , \45615 );
xor \U$45274 ( \45617 , \44411 , \44732 );
xor \U$45275 ( \45618 , \45617 , \44755 );
xor \U$45276 ( \45619 , \45616 , \45618 );
xor \U$45277 ( \45620 , \44804 , \45185 );
xor \U$45278 ( \45621 , \45620 , \45190 );
and \U$45279 ( \45622 , \45619 , \45621 );
and \U$45280 ( \45623 , \45616 , \45618 );
or \U$45281 ( \45624 , \45622 , \45623 );
xor \U$45282 ( \45625 , \45193 , \45194 );
xor \U$45283 ( \45626 , \45625 , \45197 );
and \U$45284 ( \45627 , \45624 , \45626 );
and \U$45285 ( \45628 , \45221 , \45627 );
xor \U$45286 ( \45629 , \45627 , \45221 );
xor \U$45287 ( \45630 , \45624 , \45626 );
not \U$45288 ( \45631 , \45630 );
xor \U$45289 ( \45632 , \44818 , \45149 );
xor \U$45290 ( \45633 , \45632 , \45182 );
xor \U$45291 ( \45634 , \45059 , \45079 );
xor \U$45292 ( \45635 , \45634 , \45146 );
xor \U$45293 ( \45636 , \45598 , \45600 );
xor \U$45294 ( \45637 , \45636 , \45605 );
and \U$45295 ( \45638 , \45635 , \45637 );
xor \U$45296 ( \45639 , \45233 , \45568 );
xor \U$45297 ( \45640 , \45639 , \45593 );
xor \U$45298 ( \45641 , \45598 , \45600 );
xor \U$45299 ( \45642 , \45641 , \45605 );
and \U$45300 ( \45643 , \45640 , \45642 );
and \U$45301 ( \45644 , \45635 , \45640 );
or \U$45302 ( \45645 , \45638 , \45643 , \45644 );
xor \U$45303 ( \45646 , \45633 , \45645 );
xor \U$45304 ( \45647 , \45485 , \45508 );
xor \U$45305 ( \45648 , \45647 , \45534 );
xor \U$45306 ( \45649 , \45402 , \45428 );
xor \U$45307 ( \45650 , \45649 , \45456 );
and \U$45308 ( \45651 , \45648 , \45650 );
xor \U$45309 ( \45652 , \45319 , \45346 );
xor \U$45310 ( \45653 , \45652 , \45373 );
xor \U$45311 ( \45654 , \45402 , \45428 );
xor \U$45312 ( \45655 , \45654 , \45456 );
and \U$45313 ( \45656 , \45653 , \45655 );
and \U$45314 ( \45657 , \45648 , \45653 );
or \U$45315 ( \45658 , \45651 , \45656 , \45657 );
xor \U$45316 ( \45659 , \45000 , \45027 );
xor \U$45317 ( \45660 , \45659 , \45053 );
xor \U$45318 ( \45661 , \45658 , \45660 );
xor \U$45319 ( \45662 , \45247 , \45249 );
xor \U$45320 ( \45663 , \45662 , \45277 );
xor \U$45321 ( \45664 , \45283 , \45285 );
xor \U$45322 ( \45665 , \45664 , \45288 );
and \U$45323 ( \45666 , \45663 , \45665 );
xor \U$45324 ( \45667 , \44851 , \44859 );
xor \U$45325 ( \45668 , \45667 , \44868 );
xor \U$45326 ( \45669 , \45235 , \45240 );
xor \U$45327 ( \45670 , \45668 , \45669 );
xor \U$45328 ( \45671 , \45283 , \45285 );
xor \U$45329 ( \45672 , \45671 , \45288 );
and \U$45330 ( \45673 , \45670 , \45672 );
and \U$45331 ( \45674 , \45663 , \45670 );
or \U$45332 ( \45675 , \45666 , \45673 , \45674 );
and \U$45333 ( \45676 , \45661 , \45675 );
and \U$45334 ( \45677 , \45658 , \45660 );
or \U$45335 ( \45678 , \45676 , \45677 );
xor \U$45336 ( \45679 , \45492 , \45497 );
xor \U$45337 ( \45680 , \45679 , \45505 );
xor \U$45338 ( \45681 , \45516 , \45523 );
xor \U$45339 ( \45682 , \45681 , \45531 );
and \U$45340 ( \45683 , \45680 , \45682 );
xor \U$45341 ( \45684 , \45467 , \45474 );
xor \U$45342 ( \45685 , \45684 , \45482 );
xor \U$45343 ( \45686 , \45516 , \45523 );
xor \U$45344 ( \45687 , \45686 , \45531 );
and \U$45345 ( \45688 , \45685 , \45687 );
and \U$45346 ( \45689 , \45680 , \45685 );
or \U$45347 ( \45690 , \45683 , \45688 , \45689 );
xor \U$45348 ( \45691 , \44933 , \13358 );
xor \U$45349 ( \45692 , \45691 , \44941 );
xor \U$45350 ( \45693 , \45690 , \45692 );
xor \U$45351 ( \45694 , \44908 , \44915 );
xor \U$45352 ( \45695 , \45694 , \44923 );
xor \U$45353 ( \45696 , \45543 , \45548 );
xor \U$45354 ( \45697 , \45695 , \45696 );
and \U$45355 ( \45698 , \45693 , \45697 );
and \U$45356 ( \45699 , \45690 , \45692 );
or \U$45357 ( \45700 , \45698 , \45699 );
and \U$45358 ( \45701 , \2464 , RI9871758_126);
and \U$45359 ( \45702 , RI9871848_128, \2462 );
nor \U$45360 ( \45703 , \45701 , \45702 );
and \U$45361 ( \45704 , \45703 , \2468 );
not \U$45362 ( \45705 , \45703 );
and \U$45363 ( \45706 , \45705 , \2263 );
nor \U$45364 ( \45707 , \45704 , \45706 );
not \U$45365 ( \45708 , \1462 );
and \U$45366 ( \45709 , \2042 , RI98712a8_116);
and \U$45367 ( \45710 , RI98711b8_114, \2040 );
nor \U$45368 ( \45711 , \45709 , \45710 );
not \U$45369 ( \45712 , \45711 );
or \U$45370 ( \45713 , \45708 , \45712 );
or \U$45371 ( \45714 , \45711 , \2034 );
nand \U$45372 ( \45715 , \45713 , \45714 );
xor \U$45373 ( \45716 , \45707 , \45715 );
and \U$45374 ( \45717 , \2274 , RI9871398_118);
and \U$45375 ( \45718 , RI9871488_120, \2272 );
nor \U$45376 ( \45719 , \45717 , \45718 );
and \U$45377 ( \45720 , \45719 , \2030 );
not \U$45378 ( \45721 , \45719 );
and \U$45379 ( \45722 , \45721 , \2031 );
nor \U$45380 ( \45723 , \45720 , \45722 );
and \U$45381 ( \45724 , \45716 , \45723 );
and \U$45382 ( \45725 , \45707 , \45715 );
or \U$45383 ( \45726 , \45724 , \45725 );
and \U$45384 ( \45727 , \1311 , RI98710c8_112);
and \U$45385 ( \45728 , RI9870d08_104, \1309 );
nor \U$45386 ( \45729 , \45727 , \45728 );
and \U$45387 ( \45730 , \45729 , \1458 );
not \U$45388 ( \45731 , \45729 );
and \U$45389 ( \45732 , \45731 , \1318 );
nor \U$45390 ( \45733 , \45730 , \45732 );
not \U$45391 ( \45734 , \1128 );
and \U$45392 ( \45735 , \1293 , RI9870df8_106);
and \U$45393 ( \45736 , RI9870a38_98, \1291 );
nor \U$45394 ( \45737 , \45735 , \45736 );
not \U$45395 ( \45738 , \45737 );
or \U$45396 ( \45739 , \45734 , \45738 );
or \U$45397 ( \45740 , \45737 , \1301 );
nand \U$45398 ( \45741 , \45739 , \45740 );
xor \U$45399 ( \45742 , \45733 , \45741 );
and \U$45400 ( \45743 , \1329 , RI9870ee8_108);
and \U$45401 ( \45744 , RI9870c18_102, \1327 );
nor \U$45402 ( \45745 , \45743 , \45744 );
and \U$45403 ( \45746 , \45745 , \1336 );
not \U$45404 ( \45747 , \45745 );
and \U$45405 ( \45748 , \45747 , \1337 );
nor \U$45406 ( \45749 , \45746 , \45748 );
and \U$45407 ( \45750 , \45742 , \45749 );
and \U$45408 ( \45751 , \45733 , \45741 );
or \U$45409 ( \45752 , \45750 , \45751 );
xor \U$45410 ( \45753 , \45726 , \45752 );
and \U$45411 ( \45754 , \776 , RI9870fd8_110);
and \U$45412 ( \45755 , RI9870b28_100, \774 );
nor \U$45413 ( \45756 , \45754 , \45755 );
and \U$45414 ( \45757 , \45756 , \474 );
not \U$45415 ( \45758 , \45756 );
and \U$45416 ( \45759 , \45758 , \451 );
nor \U$45417 ( \45760 , \45757 , \45759 );
and \U$45418 ( \45761 , \438 , RI98700d8_78);
and \U$45419 ( \45762 , RI98701c8_80, \436 );
nor \U$45420 ( \45763 , \45761 , \45762 );
and \U$45421 ( \45764 , \45763 , \444 );
not \U$45422 ( \45765 , \45763 );
and \U$45423 ( \45766 , \45765 , \443 );
nor \U$45424 ( \45767 , \45764 , \45766 );
xor \U$45425 ( \45768 , \45760 , \45767 );
not \U$45426 ( \45769 , \454 );
and \U$45427 ( \45770 , \465 , RI986ffe8_76);
and \U$45428 ( \45771 , RI986fef8_74, \463 );
nor \U$45429 ( \45772 , \45770 , \45771 );
not \U$45430 ( \45773 , \45772 );
or \U$45431 ( \45774 , \45769 , \45773 );
or \U$45432 ( \45775 , \45772 , \454 );
nand \U$45433 ( \45776 , \45774 , \45775 );
and \U$45434 ( \45777 , \45768 , \45776 );
and \U$45435 ( \45778 , \45760 , \45767 );
or \U$45436 ( \45779 , \45777 , \45778 );
and \U$45437 ( \45780 , \45753 , \45779 );
and \U$45438 ( \45781 , \45726 , \45752 );
or \U$45439 ( \45782 , \45780 , \45781 );
and \U$45440 ( \45783 , \12293 , RI986de28_4);
and \U$45441 ( \45784 , RI986dd38_2, \12291 );
nor \U$45442 ( \45785 , \45783 , \45784 );
and \U$45443 ( \45786 , \45785 , \11687 );
not \U$45444 ( \45787 , \45785 );
and \U$45445 ( \45788 , \45787 , \11686 );
nor \U$45446 ( \45789 , \45786 , \45788 );
and \U$45447 ( \45790 , \10424 , RI986f598_54);
and \U$45448 ( \45791 , RI986f688_56, \10422 );
nor \U$45449 ( \45792 , \45790 , \45791 );
and \U$45450 ( \45793 , \45792 , \9840 );
not \U$45451 ( \45794 , \45792 );
and \U$45452 ( \45795 , \45794 , \10428 );
nor \U$45453 ( \45796 , \45793 , \45795 );
xor \U$45454 ( \45797 , \45789 , \45796 );
and \U$45455 ( \45798 , \11696 , RI986e008_8);
and \U$45456 ( \45799 , RI986df18_6, \11694 );
nor \U$45457 ( \45800 , \45798 , \45799 );
and \U$45458 ( \45801 , \45800 , \10965 );
not \U$45459 ( \45802 , \45800 );
and \U$45460 ( \45803 , \45802 , \11702 );
nor \U$45461 ( \45804 , \45801 , \45803 );
and \U$45462 ( \45805 , \45797 , \45804 );
and \U$45463 ( \45806 , \45789 , \45796 );
or \U$45464 ( \45807 , \45805 , \45806 );
and \U$45465 ( \45808 , \13882 , RI986e2d8_14);
and \U$45466 ( \45809 , RI986e3c8_16, \13880 );
nor \U$45467 ( \45810 , \45808 , \45809 );
and \U$45468 ( \45811 , \45810 , \13358 );
not \U$45469 ( \45812 , \45810 );
and \U$45470 ( \45813 , \45812 , \13359 );
nor \U$45471 ( \45814 , \45811 , \45813 );
xor \U$45472 ( \45815 , \45814 , \14539 );
and \U$45473 ( \45816 , \13045 , RI986e1e8_12);
and \U$45474 ( \45817 , RI986e0f8_10, \13043 );
nor \U$45475 ( \45818 , \45816 , \45817 );
and \U$45476 ( \45819 , \45818 , \13047 );
not \U$45477 ( \45820 , \45818 );
and \U$45478 ( \45821 , \45820 , \12619 );
nor \U$45479 ( \45822 , \45819 , \45821 );
and \U$45480 ( \45823 , \45815 , \45822 );
and \U$45481 ( \45824 , \45814 , \14539 );
or \U$45482 ( \45825 , \45823 , \45824 );
xor \U$45483 ( \45826 , \45807 , \45825 );
and \U$45484 ( \45827 , \9237 , RI986fa48_64);
and \U$45485 ( \45828 , RI986f958_62, \9235 );
nor \U$45486 ( \45829 , \45827 , \45828 );
and \U$45487 ( \45830 , \45829 , \9241 );
not \U$45488 ( \45831 , \45829 );
and \U$45489 ( \45832 , \45831 , \8836 );
nor \U$45490 ( \45833 , \45830 , \45832 );
and \U$45491 ( \45834 , \8486 , RI986f868_60);
and \U$45492 ( \45835 , RI986f778_58, \8484 );
nor \U$45493 ( \45836 , \45834 , \45835 );
and \U$45494 ( \45837 , \45836 , \8050 );
not \U$45495 ( \45838 , \45836 );
and \U$45496 ( \45839 , \45838 , \8051 );
nor \U$45497 ( \45840 , \45837 , \45839 );
xor \U$45498 ( \45841 , \45833 , \45840 );
and \U$45499 ( \45842 , \9505 , RI986f4a8_52);
and \U$45500 ( \45843 , RI986f3b8_50, \9503 );
nor \U$45501 ( \45844 , \45842 , \45843 );
and \U$45502 ( \45845 , \45844 , \9510 );
not \U$45503 ( \45846 , \45844 );
and \U$45504 ( \45847 , \45846 , \9513 );
nor \U$45505 ( \45848 , \45845 , \45847 );
and \U$45506 ( \45849 , \45841 , \45848 );
and \U$45507 ( \45850 , \45833 , \45840 );
or \U$45508 ( \45851 , \45849 , \45850 );
and \U$45509 ( \45852 , \45826 , \45851 );
and \U$45510 ( \45853 , \45807 , \45825 );
or \U$45511 ( \45854 , \45852 , \45853 );
xor \U$45512 ( \45855 , \45782 , \45854 );
and \U$45513 ( \45856 , \5881 , RI986f0e8_44);
and \U$45514 ( \45857 , RI986eff8_42, \5879 );
nor \U$45515 ( \45858 , \45856 , \45857 );
and \U$45516 ( \45859 , \45858 , \5594 );
not \U$45517 ( \45860 , \45858 );
and \U$45518 ( \45861 , \45860 , \5885 );
nor \U$45519 ( \45862 , \45859 , \45861 );
not \U$45520 ( \45863 , \4521 );
and \U$45521 ( \45864 , \4710 , RI986ef08_40);
and \U$45522 ( \45865 , RI986ee18_38, \4708 );
nor \U$45523 ( \45866 , \45864 , \45865 );
not \U$45524 ( \45867 , \45866 );
or \U$45525 ( \45868 , \45863 , \45867 );
or \U$45526 ( \45869 , \45866 , \4521 );
nand \U$45527 ( \45870 , \45868 , \45869 );
xor \U$45528 ( \45871 , \45862 , \45870 );
and \U$45529 ( \45872 , \5318 , RI986ec38_34);
and \U$45530 ( \45873 , RI986ed28_36, \5316 );
nor \U$45531 ( \45874 , \45872 , \45873 );
and \U$45532 ( \45875 , \45874 , \5052 );
not \U$45533 ( \45876 , \45874 );
and \U$45534 ( \45877 , \45876 , \5322 );
nor \U$45535 ( \45878 , \45875 , \45877 );
and \U$45536 ( \45879 , \45871 , \45878 );
and \U$45537 ( \45880 , \45862 , \45870 );
or \U$45538 ( \45881 , \45879 , \45880 );
not \U$45539 ( \45882 , \2935 );
and \U$45540 ( \45883 , \3254 , RI9871578_122);
and \U$45541 ( \45884 , RI9871668_124, \3252 );
nor \U$45542 ( \45885 , \45883 , \45884 );
not \U$45543 ( \45886 , \45885 );
or \U$45544 ( \45887 , \45882 , \45886 );
or \U$45545 ( \45888 , \45885 , \2935 );
nand \U$45546 ( \45889 , \45887 , \45888 );
not \U$45547 ( \45890 , \3412 );
and \U$45548 ( \45891 , \3683 , RI986eb48_32);
and \U$45549 ( \45892 , RI986ea58_30, \3681 );
nor \U$45550 ( \45893 , \45891 , \45892 );
not \U$45551 ( \45894 , \45893 );
or \U$45552 ( \45895 , \45890 , \45894 );
or \U$45553 ( \45896 , \45893 , \3412 );
nand \U$45554 ( \45897 , \45895 , \45896 );
xor \U$45555 ( \45898 , \45889 , \45897 );
and \U$45556 ( \45899 , \4203 , RI986e968_28);
and \U$45557 ( \45900 , RI986e878_26, \4201 );
nor \U$45558 ( \45901 , \45899 , \45900 );
and \U$45559 ( \45902 , \45901 , \4207 );
not \U$45560 ( \45903 , \45901 );
and \U$45561 ( \45904 , \45903 , \3922 );
nor \U$45562 ( \45905 , \45902 , \45904 );
and \U$45563 ( \45906 , \45898 , \45905 );
and \U$45564 ( \45907 , \45889 , \45897 );
or \U$45565 ( \45908 , \45906 , \45907 );
xor \U$45566 ( \45909 , \45881 , \45908 );
and \U$45567 ( \45910 , \7079 , RI986e5a8_20);
and \U$45568 ( \45911 , RI986e4b8_18, \7077 );
nor \U$45569 ( \45912 , \45910 , \45911 );
and \U$45570 ( \45913 , \45912 , \6710 );
not \U$45571 ( \45914 , \45912 );
and \U$45572 ( \45915 , \45914 , \6709 );
nor \U$45573 ( \45916 , \45913 , \45915 );
and \U$45574 ( \45917 , \6453 , RI986f2c8_48);
and \U$45575 ( \45918 , RI986f1d8_46, \6451 );
nor \U$45576 ( \45919 , \45917 , \45918 );
and \U$45577 ( \45920 , \45919 , \6190 );
not \U$45578 ( \45921 , \45919 );
and \U$45579 ( \45922 , \45921 , \6180 );
nor \U$45580 ( \45923 , \45920 , \45922 );
xor \U$45581 ( \45924 , \45916 , \45923 );
and \U$45582 ( \45925 , \7729 , RI986e788_24);
and \U$45583 ( \45926 , RI986e698_22, \7727 );
nor \U$45584 ( \45927 , \45925 , \45926 );
and \U$45585 ( \45928 , \45927 , \7480 );
not \U$45586 ( \45929 , \45927 );
and \U$45587 ( \45930 , \45929 , \7733 );
nor \U$45588 ( \45931 , \45928 , \45930 );
and \U$45589 ( \45932 , \45924 , \45931 );
and \U$45590 ( \45933 , \45916 , \45923 );
or \U$45591 ( \45934 , \45932 , \45933 );
and \U$45592 ( \45935 , \45909 , \45934 );
and \U$45593 ( \45936 , \45881 , \45908 );
or \U$45594 ( \45937 , \45935 , \45936 );
and \U$45595 ( \45938 , \45855 , \45937 );
and \U$45596 ( \45939 , \45782 , \45854 );
or \U$45597 ( \45940 , \45938 , \45939 );
xor \U$45598 ( \45941 , \45700 , \45940 );
xor \U$45599 ( \45942 , \45409 , \45416 );
xor \U$45600 ( \45943 , \45942 , \45425 );
xor \U$45601 ( \45944 , \45437 , \45444 );
xor \U$45602 ( \45945 , \45944 , \45453 );
and \U$45603 ( \45946 , \45943 , \45945 );
xor \U$45604 ( \45947 , \45383 , \45390 );
xor \U$45605 ( \45948 , \45947 , \45399 );
xor \U$45606 ( \45949 , \45437 , \45444 );
xor \U$45607 ( \45950 , \45949 , \45453 );
and \U$45608 ( \45951 , \45948 , \45950 );
and \U$45609 ( \45952 , \45943 , \45948 );
or \U$45610 ( \45953 , \45946 , \45951 , \45952 );
not \U$45611 ( \45954 , \367 );
and \U$45612 ( \45955 , \376 , RI986fe08_72);
and \U$45613 ( \45956 , RI986fd18_70, \374 );
nor \U$45614 ( \45957 , \45955 , \45956 );
not \U$45615 ( \45958 , \45957 );
or \U$45616 ( \45959 , \45954 , \45958 );
or \U$45617 ( \45960 , \45957 , \365 );
nand \U$45618 ( \45961 , \45959 , \45960 );
not \U$45619 ( \45962 , \487 );
and \U$45620 ( \45963 , \395 , RI986fb38_66);
and \U$45621 ( \45964 , RI986fc28_68, \393 );
nor \U$45622 ( \45965 , \45963 , \45964 );
not \U$45623 ( \45966 , \45965 );
or \U$45624 ( \45967 , \45962 , \45966 );
or \U$45625 ( \45968 , \45965 , \386 );
nand \U$45626 ( \45969 , \45967 , \45968 );
xor \U$45627 ( \45970 , \45961 , \45969 );
not \U$45628 ( \45971 , \345 );
and \U$45629 ( \45972 , \354 , RI9870948_96);
and \U$45630 ( \45973 , RI9870858_94, \352 );
nor \U$45631 ( \45974 , \45972 , \45973 );
not \U$45632 ( \45975 , \45974 );
or \U$45633 ( \45976 , \45971 , \45975 );
or \U$45634 ( \45977 , \45974 , \361 );
nand \U$45635 ( \45978 , \45976 , \45977 );
and \U$45636 ( \45979 , \45970 , \45978 );
and \U$45637 ( \45980 , \45961 , \45969 );
or \U$45638 ( \45981 , \45979 , \45980 );
xor \U$45639 ( \45982 , \45981 , \45246 );
xor \U$45640 ( \45983 , \45258 , \45266 );
xor \U$45641 ( \45984 , \45983 , \45274 );
and \U$45642 ( \45985 , \45982 , \45984 );
and \U$45643 ( \45986 , \45981 , \45246 );
or \U$45644 ( \45987 , \45985 , \45986 );
xor \U$45645 ( \45988 , \45953 , \45987 );
xor \U$45646 ( \45989 , \45327 , \45334 );
xor \U$45647 ( \45990 , \45989 , \45343 );
xor \U$45648 ( \45991 , \45355 , \45362 );
xor \U$45649 ( \45992 , \45991 , \45370 );
xor \U$45650 ( \45993 , \45990 , \45992 );
xor \U$45651 ( \45994 , \45301 , \45308 );
xor \U$45652 ( \45995 , \45994 , \45316 );
and \U$45653 ( \45996 , \45993 , \45995 );
and \U$45654 ( \45997 , \45990 , \45992 );
or \U$45655 ( \45998 , \45996 , \45997 );
and \U$45656 ( \45999 , \45988 , \45998 );
and \U$45657 ( \46000 , \45953 , \45987 );
or \U$45658 ( \46001 , \45999 , \46000 );
and \U$45659 ( \46002 , \45941 , \46001 );
and \U$45660 ( \46003 , \45700 , \45940 );
or \U$45661 ( \46004 , \46002 , \46003 );
xor \U$45662 ( \46005 , \45678 , \46004 );
xor \U$45663 ( \46006 , \44926 , \44944 );
xor \U$45664 ( \46007 , \46006 , \44970 );
xor \U$45665 ( \46008 , \45571 , \45573 );
xor \U$45666 ( \46009 , \46008 , \45578 );
and \U$45667 ( \46010 , \46007 , \46009 );
xor \U$45668 ( \46011 , \45066 , \45068 );
xor \U$45669 ( \46012 , \46011 , \45071 );
xor \U$45670 ( \46013 , \45553 , \45560 );
xor \U$45671 ( \46014 , \46012 , \46013 );
xor \U$45672 ( \46015 , \45571 , \45573 );
xor \U$45673 ( \46016 , \46015 , \45578 );
and \U$45674 ( \46017 , \46014 , \46016 );
and \U$45675 ( \46018 , \46007 , \46014 );
or \U$45676 ( \46019 , \46010 , \46017 , \46018 );
and \U$45677 ( \46020 , \46005 , \46019 );
and \U$45678 ( \46021 , \45678 , \46004 );
or \U$45679 ( \46022 , \46020 , \46021 );
xor \U$45680 ( \46023 , \45160 , \45162 );
xor \U$45681 ( \46024 , \46023 , \45179 );
xor \U$45682 ( \46025 , \46022 , \46024 );
xor \U$45683 ( \46026 , \45294 , \45540 );
xor \U$45684 ( \46027 , \46026 , \45565 );
xor \U$45685 ( \46028 , \45225 , \45227 );
xor \U$45686 ( \46029 , \46028 , \45230 );
and \U$45687 ( \46030 , \46027 , \46029 );
xor \U$45688 ( \46031 , \45152 , \45154 );
xor \U$45689 ( \46032 , \46031 , \45157 );
xor \U$45690 ( \46033 , \45581 , \45588 );
xor \U$45691 ( \46034 , \46032 , \46033 );
xor \U$45692 ( \46035 , \45225 , \45227 );
xor \U$45693 ( \46036 , \46035 , \45230 );
and \U$45694 ( \46037 , \46034 , \46036 );
and \U$45695 ( \46038 , \46027 , \46034 );
or \U$45696 ( \46039 , \46030 , \46037 , \46038 );
and \U$45697 ( \46040 , \46025 , \46039 );
and \U$45698 ( \46041 , \46022 , \46024 );
or \U$45699 ( \46042 , \46040 , \46041 );
and \U$45700 ( \46043 , \45646 , \46042 );
and \U$45701 ( \46044 , \45633 , \45645 );
nor \U$45702 ( \46045 , \46043 , \46044 );
not \U$45703 ( \46046 , \46045 );
xor \U$45704 ( \46047 , \45616 , \45618 );
xor \U$45705 ( \46048 , \46047 , \45621 );
nand \U$45706 ( \46049 , \46046 , \46048 );
or \U$45707 ( \46050 , \45631 , \46049 );
not \U$45708 ( \46051 , \45630 );
not \U$45709 ( \46052 , \46049 );
and \U$45710 ( \46053 , \46051 , \46052 );
and \U$45711 ( \46054 , \45630 , \46049 );
nor \U$45712 ( \46055 , \46053 , \46054 );
xor \U$45713 ( \46056 , \45760 , \45767 );
xor \U$45714 ( \46057 , \46056 , \45776 );
not \U$45715 ( \46058 , RI98702b8_82);
nor \U$45716 ( \46059 , \46058 , \407 );
xor \U$45717 ( \46060 , \46057 , \46059 );
xor \U$45718 ( \46061 , \45961 , \45969 );
xor \U$45719 ( \46062 , \46061 , \45978 );
and \U$45720 ( \46063 , \46060 , \46062 );
and \U$45721 ( \46064 , \46057 , \46059 );
or \U$45722 ( \46065 , \46063 , \46064 );
nand \U$45723 ( \46066 , RI98703a8_84, RI9871fc8_144);
and \U$45724 ( \46067 , \416 , RI98702b8_82);
and \U$45725 ( \46068 , RI9870768_92, \414 );
nor \U$45726 ( \46069 , \46067 , \46068 );
and \U$45727 ( \46070 , \46069 , \421 );
not \U$45728 ( \46071 , \46069 );
and \U$45729 ( \46072 , \46071 , \422 );
nor \U$45730 ( \46073 , \46070 , \46072 );
nand \U$45731 ( \46074 , \46066 , \46073 );
and \U$45732 ( \46075 , \416 , RI9870768_92);
and \U$45733 ( \46076 , RI9870678_90, \414 );
nor \U$45734 ( \46077 , \46075 , \46076 );
and \U$45735 ( \46078 , \46077 , \422 );
not \U$45736 ( \46079 , \46077 );
and \U$45737 ( \46080 , \46079 , \421 );
nor \U$45738 ( \46081 , \46078 , \46080 );
xor \U$45739 ( \46082 , \46074 , \46081 );
and \U$45740 ( \46083 , \395 , RI9870858_94);
and \U$45741 ( \46084 , RI986fb38_66, \393 );
nor \U$45742 ( \46085 , \46083 , \46084 );
not \U$45743 ( \46086 , \46085 );
not \U$45744 ( \46087 , \386 );
and \U$45745 ( \46088 , \46086 , \46087 );
and \U$45746 ( \46089 , \46085 , \386 );
nor \U$45747 ( \46090 , \46088 , \46089 );
and \U$45748 ( \46091 , \354 , RI9870678_90);
and \U$45749 ( \46092 , RI9870948_96, \352 );
nor \U$45750 ( \46093 , \46091 , \46092 );
not \U$45751 ( \46094 , \46093 );
not \U$45752 ( \46095 , \361 );
and \U$45753 ( \46096 , \46094 , \46095 );
and \U$45754 ( \46097 , \46093 , \345 );
nor \U$45755 ( \46098 , \46096 , \46097 );
or \U$45756 ( \46099 , \46090 , \46098 );
not \U$45757 ( \46100 , \46098 );
not \U$45758 ( \46101 , \46090 );
or \U$45759 ( \46102 , \46100 , \46101 );
not \U$45760 ( \46103 , \365 );
and \U$45761 ( \46104 , \376 , RI986fc28_68);
and \U$45762 ( \46105 , RI986fe08_72, \374 );
nor \U$45763 ( \46106 , \46104 , \46105 );
not \U$45764 ( \46107 , \46106 );
or \U$45765 ( \46108 , \46103 , \46107 );
or \U$45766 ( \46109 , \46106 , \365 );
nand \U$45767 ( \46110 , \46108 , \46109 );
nand \U$45768 ( \46111 , \46102 , \46110 );
nand \U$45769 ( \46112 , \46099 , \46111 );
and \U$45770 ( \46113 , \46082 , \46112 );
and \U$45771 ( \46114 , \46074 , \46081 );
or \U$45772 ( \46115 , \46113 , \46114 );
xor \U$45773 ( \46116 , \46065 , \46115 );
xor \U$45774 ( \46117 , \45707 , \45715 );
xor \U$45775 ( \46118 , \46117 , \45723 );
xor \U$45776 ( \46119 , \45733 , \45741 );
xor \U$45777 ( \46120 , \46119 , \45749 );
and \U$45778 ( \46121 , \46118 , \46120 );
xor \U$45779 ( \46122 , \45889 , \45897 );
xor \U$45780 ( \46123 , \46122 , \45905 );
xor \U$45781 ( \46124 , \45733 , \45741 );
xor \U$45782 ( \46125 , \46124 , \45749 );
and \U$45783 ( \46126 , \46123 , \46125 );
and \U$45784 ( \46127 , \46118 , \46123 );
or \U$45785 ( \46128 , \46121 , \46126 , \46127 );
xor \U$45786 ( \46129 , \46116 , \46128 );
xor \U$45787 ( \46130 , \45862 , \45870 );
xor \U$45788 ( \46131 , \46130 , \45878 );
xor \U$45789 ( \46132 , \45833 , \45840 );
xor \U$45790 ( \46133 , \46132 , \45848 );
and \U$45791 ( \46134 , \46131 , \46133 );
xor \U$45792 ( \46135 , \45916 , \45923 );
xor \U$45793 ( \46136 , \46135 , \45931 );
xor \U$45794 ( \46137 , \45833 , \45840 );
xor \U$45795 ( \46138 , \46137 , \45848 );
and \U$45796 ( \46139 , \46136 , \46138 );
and \U$45797 ( \46140 , \46131 , \46136 );
or \U$45798 ( \46141 , \46134 , \46139 , \46140 );
xor \U$45799 ( \46142 , \45789 , \45796 );
xor \U$45800 ( \46143 , \46142 , \45804 );
xor \U$45801 ( \46144 , \45814 , \14539 );
xor \U$45802 ( \46145 , \46144 , \45822 );
and \U$45803 ( \46146 , \46143 , \46145 );
xor \U$45804 ( \46147 , \46141 , \46146 );
xor \U$45805 ( \46148 , \45516 , \45523 );
xor \U$45806 ( \46149 , \46148 , \45531 );
xor \U$45807 ( \46150 , \45680 , \45685 );
xor \U$45808 ( \46151 , \46149 , \46150 );
xor \U$45809 ( \46152 , \46147 , \46151 );
and \U$45810 ( \46153 , \46129 , \46152 );
xor \U$45811 ( \46154 , \45990 , \45992 );
xor \U$45812 ( \46155 , \46154 , \45995 );
xor \U$45813 ( \46156 , \45981 , \45246 );
xor \U$45814 ( \46157 , \46156 , \45984 );
xor \U$45815 ( \46158 , \45437 , \45444 );
xor \U$45816 ( \46159 , \46158 , \45453 );
xor \U$45817 ( \46160 , \45943 , \45948 );
xor \U$45818 ( \46161 , \46159 , \46160 );
xor \U$45819 ( \46162 , \46157 , \46161 );
xor \U$45820 ( \46163 , \46155 , \46162 );
xor \U$45821 ( \46164 , \46141 , \46146 );
xor \U$45822 ( \46165 , \46164 , \46151 );
and \U$45823 ( \46166 , \46163 , \46165 );
and \U$45824 ( \46167 , \46129 , \46163 );
or \U$45825 ( \46168 , \46153 , \46166 , \46167 );
not \U$45826 ( \46169 , \46168 );
xor \U$45827 ( \46170 , \46074 , \46081 );
xor \U$45828 ( \46171 , \46170 , \46112 );
xor \U$45829 ( \46172 , \46057 , \46059 );
xor \U$45830 ( \46173 , \46172 , \46062 );
and \U$45831 ( \46174 , \46171 , \46173 );
xor \U$45832 ( \46175 , \45733 , \45741 );
xor \U$45833 ( \46176 , \46175 , \45749 );
xor \U$45834 ( \46177 , \46118 , \46123 );
xor \U$45835 ( \46178 , \46176 , \46177 );
xor \U$45836 ( \46179 , \46057 , \46059 );
xor \U$45837 ( \46180 , \46179 , \46062 );
and \U$45838 ( \46181 , \46178 , \46180 );
and \U$45839 ( \46182 , \46171 , \46178 );
or \U$45840 ( \46183 , \46174 , \46181 , \46182 );
and \U$45841 ( \46184 , \13045 , RI986dd38_2);
and \U$45842 ( \46185 , RI986e1e8_12, \13043 );
nor \U$45843 ( \46186 , \46184 , \46185 );
and \U$45844 ( \46187 , \46186 , \12619 );
not \U$45845 ( \46188 , \46186 );
and \U$45846 ( \46189 , \46188 , \13047 );
nor \U$45847 ( \46190 , \46187 , \46189 );
not \U$45848 ( \46191 , \46190 );
and \U$45849 ( \46192 , \13882 , RI986e0f8_10);
and \U$45850 ( \46193 , RI986e2d8_14, \13880 );
nor \U$45851 ( \46194 , \46192 , \46193 );
and \U$45852 ( \46195 , \46194 , \13359 );
not \U$45853 ( \46196 , \46194 );
and \U$45854 ( \46197 , \46196 , \13358 );
nor \U$45855 ( \46198 , \46195 , \46197 );
not \U$45856 ( \46199 , \46198 );
and \U$45857 ( \46200 , \46191 , \46199 );
and \U$45858 ( \46201 , \46198 , \46190 );
nand \U$45859 ( \46202 , RI986e3c8_16, \14937 );
and \U$45860 ( \46203 , \46202 , \14538 );
not \U$45861 ( \46204 , \46202 );
and \U$45862 ( \46205 , \46204 , \14539 );
nor \U$45863 ( \46206 , \46203 , \46205 );
nor \U$45864 ( \46207 , \46201 , \46206 );
nor \U$45865 ( \46208 , \46200 , \46207 );
and \U$45866 ( \46209 , \9505 , RI986f958_62);
and \U$45867 ( \46210 , RI986f4a8_52, \9503 );
nor \U$45868 ( \46211 , \46209 , \46210 );
and \U$45869 ( \46212 , \46211 , \9513 );
not \U$45870 ( \46213 , \46211 );
and \U$45871 ( \46214 , \46213 , \9510 );
nor \U$45872 ( \46215 , \46212 , \46214 );
and \U$45873 ( \46216 , \8486 , RI986e698_22);
and \U$45874 ( \46217 , RI986f868_60, \8484 );
nor \U$45875 ( \46218 , \46216 , \46217 );
and \U$45876 ( \46219 , \46218 , \8051 );
not \U$45877 ( \46220 , \46218 );
and \U$45878 ( \46221 , \46220 , \8050 );
nor \U$45879 ( \46222 , \46219 , \46221 );
xor \U$45880 ( \46223 , \46215 , \46222 );
and \U$45881 ( \46224 , \9237 , RI986f778_58);
and \U$45882 ( \46225 , RI986fa48_64, \9235 );
nor \U$45883 ( \46226 , \46224 , \46225 );
and \U$45884 ( \46227 , \46226 , \8836 );
not \U$45885 ( \46228 , \46226 );
and \U$45886 ( \46229 , \46228 , \9241 );
nor \U$45887 ( \46230 , \46227 , \46229 );
and \U$45888 ( \46231 , \46223 , \46230 );
and \U$45889 ( \46232 , \46215 , \46222 );
or \U$45890 ( \46233 , \46231 , \46232 );
xor \U$45891 ( \46234 , \46208 , \46233 );
and \U$45892 ( \46235 , \12293 , RI986df18_6);
and \U$45893 ( \46236 , RI986de28_4, \12291 );
nor \U$45894 ( \46237 , \46235 , \46236 );
and \U$45895 ( \46238 , \46237 , \11686 );
not \U$45896 ( \46239 , \46237 );
and \U$45897 ( \46240 , \46239 , \11687 );
nor \U$45898 ( \46241 , \46238 , \46240 );
and \U$45899 ( \46242 , \10424 , RI986f3b8_50);
and \U$45900 ( \46243 , RI986f598_54, \10422 );
nor \U$45901 ( \46244 , \46242 , \46243 );
and \U$45902 ( \46245 , \46244 , \10428 );
not \U$45903 ( \46246 , \46244 );
and \U$45904 ( \46247 , \46246 , \9840 );
nor \U$45905 ( \46248 , \46245 , \46247 );
xor \U$45906 ( \46249 , \46241 , \46248 );
and \U$45907 ( \46250 , \11696 , RI986f688_56);
and \U$45908 ( \46251 , RI986e008_8, \11694 );
nor \U$45909 ( \46252 , \46250 , \46251 );
and \U$45910 ( \46253 , \46252 , \11702 );
not \U$45911 ( \46254 , \46252 );
and \U$45912 ( \46255 , \46254 , \10965 );
nor \U$45913 ( \46256 , \46253 , \46255 );
and \U$45914 ( \46257 , \46249 , \46256 );
and \U$45915 ( \46258 , \46241 , \46248 );
or \U$45916 ( \46259 , \46257 , \46258 );
xor \U$45917 ( \46260 , \46234 , \46259 );
and \U$45918 ( \46261 , \438 , RI986fef8_74);
and \U$45919 ( \46262 , RI98700d8_78, \436 );
nor \U$45920 ( \46263 , \46261 , \46262 );
and \U$45921 ( \46264 , \46263 , \443 );
not \U$45922 ( \46265 , \46263 );
and \U$45923 ( \46266 , \46265 , \444 );
nor \U$45924 ( \46267 , \46264 , \46266 );
and \U$45925 ( \46268 , \776 , RI98701c8_80);
and \U$45926 ( \46269 , RI9870fd8_110, \774 );
nor \U$45927 ( \46270 , \46268 , \46269 );
and \U$45928 ( \46271 , \46270 , \451 );
not \U$45929 ( \46272 , \46270 );
and \U$45930 ( \46273 , \46272 , \474 );
nor \U$45931 ( \46274 , \46271 , \46273 );
xor \U$45932 ( \46275 , \46267 , \46274 );
and \U$45933 ( \46276 , \465 , RI986fd18_70);
and \U$45934 ( \46277 , RI986ffe8_76, \463 );
nor \U$45935 ( \46278 , \46276 , \46277 );
not \U$45936 ( \46279 , \46278 );
not \U$45937 ( \46280 , \456 );
and \U$45938 ( \46281 , \46279 , \46280 );
and \U$45939 ( \46282 , \46278 , \456 );
nor \U$45940 ( \46283 , \46281 , \46282 );
and \U$45941 ( \46284 , \46275 , \46283 );
and \U$45942 ( \46285 , \46267 , \46274 );
or \U$45943 ( \46286 , \46284 , \46285 );
and \U$45944 ( \46287 , \2464 , RI9871488_120);
and \U$45945 ( \46288 , RI9871758_126, \2462 );
nor \U$45946 ( \46289 , \46287 , \46288 );
and \U$45947 ( \46290 , \46289 , \2263 );
not \U$45948 ( \46291 , \46289 );
and \U$45949 ( \46292 , \46291 , \2468 );
nor \U$45950 ( \46293 , \46290 , \46292 );
and \U$45951 ( \46294 , \2042 , RI9870d08_104);
and \U$45952 ( \46295 , RI98712a8_116, \2040 );
nor \U$45953 ( \46296 , \46294 , \46295 );
not \U$45954 ( \46297 , \46296 );
not \U$45955 ( \46298 , \1462 );
and \U$45956 ( \46299 , \46297 , \46298 );
and \U$45957 ( \46300 , \46296 , \1462 );
nor \U$45958 ( \46301 , \46299 , \46300 );
xor \U$45959 ( \46302 , \46293 , \46301 );
and \U$45960 ( \46303 , \2274 , RI98711b8_114);
and \U$45961 ( \46304 , RI9871398_118, \2272 );
nor \U$45962 ( \46305 , \46303 , \46304 );
and \U$45963 ( \46306 , \46305 , \2031 );
not \U$45964 ( \46307 , \46305 );
and \U$45965 ( \46308 , \46307 , \2030 );
nor \U$45966 ( \46309 , \46306 , \46308 );
and \U$45967 ( \46310 , \46302 , \46309 );
and \U$45968 ( \46311 , \46293 , \46301 );
or \U$45969 ( \46312 , \46310 , \46311 );
xor \U$45970 ( \46313 , \46286 , \46312 );
and \U$45971 ( \46314 , \1329 , RI9870a38_98);
and \U$45972 ( \46315 , RI9870ee8_108, \1327 );
nor \U$45973 ( \46316 , \46314 , \46315 );
and \U$45974 ( \46317 , \46316 , \1337 );
not \U$45975 ( \46318 , \46316 );
and \U$45976 ( \46319 , \46318 , \1336 );
nor \U$45977 ( \46320 , \46317 , \46319 );
and \U$45978 ( \46321 , \1293 , RI9870b28_100);
and \U$45979 ( \46322 , RI9870df8_106, \1291 );
nor \U$45980 ( \46323 , \46321 , \46322 );
not \U$45981 ( \46324 , \46323 );
not \U$45982 ( \46325 , \1301 );
and \U$45983 ( \46326 , \46324 , \46325 );
and \U$45984 ( \46327 , \46323 , \1128 );
nor \U$45985 ( \46328 , \46326 , \46327 );
xor \U$45986 ( \46329 , \46320 , \46328 );
and \U$45987 ( \46330 , \1311 , RI9870c18_102);
and \U$45988 ( \46331 , RI98710c8_112, \1309 );
nor \U$45989 ( \46332 , \46330 , \46331 );
and \U$45990 ( \46333 , \46332 , \1315 );
not \U$45991 ( \46334 , \46332 );
and \U$45992 ( \46335 , \46334 , \1458 );
nor \U$45993 ( \46336 , \46333 , \46335 );
and \U$45994 ( \46337 , \46329 , \46336 );
and \U$45995 ( \46338 , \46320 , \46328 );
or \U$45996 ( \46339 , \46337 , \46338 );
xor \U$45997 ( \46340 , \46313 , \46339 );
xor \U$45998 ( \46341 , \46260 , \46340 );
and \U$45999 ( \46342 , \3683 , RI9871668_124);
and \U$46000 ( \46343 , RI986eb48_32, \3681 );
nor \U$46001 ( \46344 , \46342 , \46343 );
not \U$46002 ( \46345 , \46344 );
not \U$46003 ( \46346 , \3412 );
and \U$46004 ( \46347 , \46345 , \46346 );
and \U$46005 ( \46348 , \46344 , \3412 );
nor \U$46006 ( \46349 , \46347 , \46348 );
and \U$46007 ( \46350 , \3254 , RI9871848_128);
and \U$46008 ( \46351 , RI9871578_122, \3252 );
nor \U$46009 ( \46352 , \46350 , \46351 );
not \U$46010 ( \46353 , \46352 );
not \U$46011 ( \46354 , \3406 );
and \U$46012 ( \46355 , \46353 , \46354 );
and \U$46013 ( \46356 , \46352 , \3406 );
nor \U$46014 ( \46357 , \46355 , \46356 );
xor \U$46015 ( \46358 , \46349 , \46357 );
and \U$46016 ( \46359 , \4203 , RI986ea58_30);
and \U$46017 ( \46360 , RI986e968_28, \4201 );
nor \U$46018 ( \46361 , \46359 , \46360 );
and \U$46019 ( \46362 , \46361 , \3922 );
not \U$46020 ( \46363 , \46361 );
and \U$46021 ( \46364 , \46363 , \4207 );
nor \U$46022 ( \46365 , \46362 , \46364 );
and \U$46023 ( \46366 , \46358 , \46365 );
and \U$46024 ( \46367 , \46349 , \46357 );
or \U$46025 ( \46368 , \46366 , \46367 );
and \U$46026 ( \46369 , \7729 , RI986e4b8_18);
and \U$46027 ( \46370 , RI986e788_24, \7727 );
nor \U$46028 ( \46371 , \46369 , \46370 );
and \U$46029 ( \46372 , \46371 , \7733 );
not \U$46030 ( \46373 , \46371 );
and \U$46031 ( \46374 , \46373 , \7480 );
nor \U$46032 ( \46375 , \46372 , \46374 );
and \U$46033 ( \46376 , \6453 , RI986eff8_42);
and \U$46034 ( \46377 , RI986f2c8_48, \6451 );
nor \U$46035 ( \46378 , \46376 , \46377 );
and \U$46036 ( \46379 , \46378 , \6180 );
not \U$46037 ( \46380 , \46378 );
and \U$46038 ( \46381 , \46380 , \6190 );
nor \U$46039 ( \46382 , \46379 , \46381 );
xor \U$46040 ( \46383 , \46375 , \46382 );
and \U$46041 ( \46384 , \7079 , RI986f1d8_46);
and \U$46042 ( \46385 , RI986e5a8_20, \7077 );
nor \U$46043 ( \46386 , \46384 , \46385 );
and \U$46044 ( \46387 , \46386 , \6709 );
not \U$46045 ( \46388 , \46386 );
and \U$46046 ( \46389 , \46388 , \6710 );
nor \U$46047 ( \46390 , \46387 , \46389 );
and \U$46048 ( \46391 , \46383 , \46390 );
and \U$46049 ( \46392 , \46375 , \46382 );
or \U$46050 ( \46393 , \46391 , \46392 );
xor \U$46051 ( \46394 , \46368 , \46393 );
and \U$46052 ( \46395 , \5881 , RI986ed28_36);
and \U$46053 ( \46396 , RI986f0e8_44, \5879 );
nor \U$46054 ( \46397 , \46395 , \46396 );
and \U$46055 ( \46398 , \46397 , \5885 );
not \U$46056 ( \46399 , \46397 );
and \U$46057 ( \46400 , \46399 , \5594 );
nor \U$46058 ( \46401 , \46398 , \46400 );
and \U$46059 ( \46402 , \4710 , RI986e878_26);
and \U$46060 ( \46403 , RI986ef08_40, \4708 );
nor \U$46061 ( \46404 , \46402 , \46403 );
not \U$46062 ( \46405 , \46404 );
not \U$46063 ( \46406 , \4519 );
and \U$46064 ( \46407 , \46405 , \46406 );
and \U$46065 ( \46408 , \46404 , \4519 );
nor \U$46066 ( \46409 , \46407 , \46408 );
xor \U$46067 ( \46410 , \46401 , \46409 );
and \U$46068 ( \46411 , \5318 , RI986ee18_38);
and \U$46069 ( \46412 , RI986ec38_34, \5316 );
nor \U$46070 ( \46413 , \46411 , \46412 );
and \U$46071 ( \46414 , \46413 , \5322 );
not \U$46072 ( \46415 , \46413 );
and \U$46073 ( \46416 , \46415 , \5052 );
nor \U$46074 ( \46417 , \46414 , \46416 );
and \U$46075 ( \46418 , \46410 , \46417 );
and \U$46076 ( \46419 , \46401 , \46409 );
or \U$46077 ( \46420 , \46418 , \46419 );
xor \U$46078 ( \46421 , \46394 , \46420 );
and \U$46079 ( \46422 , \46341 , \46421 );
and \U$46080 ( \46423 , \46260 , \46340 );
nor \U$46081 ( \46424 , \46422 , \46423 );
xor \U$46082 ( \46425 , \46183 , \46424 );
xor \U$46083 ( \46426 , \45807 , \45825 );
xor \U$46084 ( \46427 , \46426 , \45851 );
xor \U$46085 ( \46428 , \45726 , \45752 );
xor \U$46086 ( \46429 , \46428 , \45779 );
xor \U$46087 ( \46430 , \45881 , \45908 );
xor \U$46088 ( \46431 , \46430 , \45934 );
xor \U$46089 ( \46432 , \46429 , \46431 );
xor \U$46090 ( \46433 , \46427 , \46432 );
and \U$46091 ( \46434 , \46425 , \46433 );
and \U$46092 ( \46435 , \46183 , \46424 );
or \U$46093 ( \46436 , \46434 , \46435 );
not \U$46094 ( \46437 , \46436 );
or \U$46095 ( \46438 , \46169 , \46437 );
or \U$46096 ( \46439 , \46436 , \46168 );
not \U$46097 ( \46440 , \46090 );
not \U$46098 ( \46441 , \46110 );
or \U$46099 ( \46442 , \46440 , \46441 );
or \U$46100 ( \46443 , \46090 , \46110 );
nand \U$46101 ( \46444 , \46442 , \46443 );
not \U$46102 ( \46445 , \46444 );
not \U$46103 ( \46446 , \46098 );
and \U$46104 ( \46447 , \46445 , \46446 );
and \U$46105 ( \46448 , \46444 , \46098 );
nor \U$46106 ( \46449 , \46447 , \46448 );
xor \U$46107 ( \46450 , \46267 , \46274 );
xor \U$46108 ( \46451 , \46450 , \46283 );
xor \U$46109 ( \46452 , \46449 , \46451 );
xor \U$46110 ( \46453 , \46320 , \46328 );
xor \U$46111 ( \46454 , \46453 , \46336 );
and \U$46112 ( \46455 , \46452 , \46454 );
and \U$46113 ( \46456 , \46449 , \46451 );
nor \U$46114 ( \46457 , \46455 , \46456 );
and \U$46115 ( \46458 , \416 , RI98703a8_84);
and \U$46116 ( \46459 , RI98702b8_82, \414 );
nor \U$46117 ( \46460 , \46458 , \46459 );
and \U$46118 ( \46461 , \46460 , \422 );
not \U$46119 ( \46462 , \46460 );
and \U$46120 ( \46463 , \46462 , \421 );
nor \U$46121 ( \46464 , \46461 , \46463 );
not \U$46122 ( \46465 , RI9870588_88);
nor \U$46123 ( \46466 , \46465 , \407 );
xor \U$46124 ( \46467 , \46464 , \46466 );
not \U$46125 ( \46468 , \345 );
and \U$46126 ( \46469 , \354 , RI9870768_92);
and \U$46127 ( \46470 , RI9870678_90, \352 );
nor \U$46128 ( \46471 , \46469 , \46470 );
not \U$46129 ( \46472 , \46471 );
or \U$46130 ( \46473 , \46468 , \46472 );
or \U$46131 ( \46474 , \46471 , \345 );
nand \U$46132 ( \46475 , \46473 , \46474 );
and \U$46133 ( \46476 , \46467 , \46475 );
and \U$46134 ( \46477 , \46464 , \46466 );
or \U$46135 ( \46478 , \46476 , \46477 );
or \U$46136 ( \46479 , \46073 , \46066 );
nand \U$46137 ( \46480 , \46479 , \46074 );
xor \U$46138 ( \46481 , \46478 , \46480 );
not \U$46139 ( \46482 , \365 );
and \U$46140 ( \46483 , \376 , RI986fb38_66);
and \U$46141 ( \46484 , RI986fc28_68, \374 );
nor \U$46142 ( \46485 , \46483 , \46484 );
not \U$46143 ( \46486 , \46485 );
or \U$46144 ( \46487 , \46482 , \46486 );
or \U$46145 ( \46488 , \46485 , \365 );
nand \U$46146 ( \46489 , \46487 , \46488 );
not \U$46147 ( \46490 , \454 );
and \U$46148 ( \46491 , \465 , RI986fe08_72);
and \U$46149 ( \46492 , RI986fd18_70, \463 );
nor \U$46150 ( \46493 , \46491 , \46492 );
not \U$46151 ( \46494 , \46493 );
or \U$46152 ( \46495 , \46490 , \46494 );
or \U$46153 ( \46496 , \46493 , \454 );
nand \U$46154 ( \46497 , \46495 , \46496 );
xor \U$46155 ( \46498 , \46489 , \46497 );
not \U$46156 ( \46499 , \487 );
and \U$46157 ( \46500 , \395 , RI9870948_96);
and \U$46158 ( \46501 , RI9870858_94, \393 );
nor \U$46159 ( \46502 , \46500 , \46501 );
not \U$46160 ( \46503 , \46502 );
or \U$46161 ( \46504 , \46499 , \46503 );
or \U$46162 ( \46505 , \46502 , \386 );
nand \U$46163 ( \46506 , \46504 , \46505 );
and \U$46164 ( \46507 , \46498 , \46506 );
and \U$46165 ( \46508 , \46489 , \46497 );
or \U$46166 ( \46509 , \46507 , \46508 );
and \U$46167 ( \46510 , \46481 , \46509 );
and \U$46168 ( \46511 , \46478 , \46480 );
or \U$46169 ( \46512 , \46510 , \46511 );
xor \U$46170 ( \46513 , \46457 , \46512 );
xor \U$46171 ( \46514 , \46349 , \46357 );
xor \U$46172 ( \46515 , \46514 , \46365 );
xor \U$46173 ( \46516 , \46401 , \46409 );
xor \U$46174 ( \46517 , \46516 , \46417 );
xor \U$46175 ( \46518 , \46515 , \46517 );
xor \U$46176 ( \46519 , \46293 , \46301 );
xor \U$46177 ( \46520 , \46519 , \46309 );
and \U$46178 ( \46521 , \46518 , \46520 );
and \U$46179 ( \46522 , \46515 , \46517 );
nor \U$46180 ( \46523 , \46521 , \46522 );
and \U$46181 ( \46524 , \46513 , \46523 );
and \U$46182 ( \46525 , \46457 , \46512 );
or \U$46183 ( \46526 , \46524 , \46525 );
and \U$46184 ( \46527 , \7079 , RI986f2c8_48);
and \U$46185 ( \46528 , RI986f1d8_46, \7077 );
nor \U$46186 ( \46529 , \46527 , \46528 );
and \U$46187 ( \46530 , \46529 , \6709 );
not \U$46188 ( \46531 , \46529 );
and \U$46189 ( \46532 , \46531 , \6710 );
nor \U$46190 ( \46533 , \46530 , \46532 );
and \U$46191 ( \46534 , \7729 , RI986e5a8_20);
and \U$46192 ( \46535 , RI986e4b8_18, \7727 );
nor \U$46193 ( \46536 , \46534 , \46535 );
and \U$46194 ( \46537 , \46536 , \7733 );
not \U$46195 ( \46538 , \46536 );
and \U$46196 ( \46539 , \46538 , \7480 );
nor \U$46197 ( \46540 , \46537 , \46539 );
or \U$46198 ( \46541 , \46533 , \46540 );
not \U$46199 ( \46542 , \46540 );
not \U$46200 ( \46543 , \46533 );
or \U$46201 ( \46544 , \46542 , \46543 );
and \U$46202 ( \46545 , \8486 , RI986e788_24);
and \U$46203 ( \46546 , RI986e698_22, \8484 );
nor \U$46204 ( \46547 , \46545 , \46546 );
and \U$46205 ( \46548 , \46547 , \8050 );
not \U$46206 ( \46549 , \46547 );
and \U$46207 ( \46550 , \46549 , \8051 );
nor \U$46208 ( \46551 , \46548 , \46550 );
nand \U$46209 ( \46552 , \46544 , \46551 );
nand \U$46210 ( \46553 , \46541 , \46552 );
and \U$46211 ( \46554 , \4203 , RI986eb48_32);
and \U$46212 ( \46555 , RI986ea58_30, \4201 );
nor \U$46213 ( \46556 , \46554 , \46555 );
and \U$46214 ( \46557 , \46556 , \3923 );
not \U$46215 ( \46558 , \46556 );
and \U$46216 ( \46559 , \46558 , \4207 );
nor \U$46217 ( \46560 , \46557 , \46559 );
and \U$46218 ( \46561 , \4710 , RI986e968_28);
and \U$46219 ( \46562 , RI986e878_26, \4708 );
nor \U$46220 ( \46563 , \46561 , \46562 );
not \U$46221 ( \46564 , \46563 );
not \U$46222 ( \46565 , \4521 );
and \U$46223 ( \46566 , \46564 , \46565 );
and \U$46224 ( \46567 , \46563 , \4521 );
nor \U$46225 ( \46568 , \46566 , \46567 );
xor \U$46226 ( \46569 , \46560 , \46568 );
and \U$46227 ( \46570 , \3683 , RI9871578_122);
and \U$46228 ( \46571 , RI9871668_124, \3681 );
nor \U$46229 ( \46572 , \46570 , \46571 );
not \U$46230 ( \46573 , \46572 );
not \U$46231 ( \46574 , \3918 );
and \U$46232 ( \46575 , \46573 , \46574 );
and \U$46233 ( \46576 , \46572 , \3918 );
nor \U$46234 ( \46577 , \46575 , \46576 );
and \U$46235 ( \46578 , \46569 , \46577 );
and \U$46236 ( \46579 , \46560 , \46568 );
nor \U$46237 ( \46580 , \46578 , \46579 );
xor \U$46238 ( \46581 , \46553 , \46580 );
and \U$46239 ( \46582 , \5318 , RI986ef08_40);
and \U$46240 ( \46583 , RI986ee18_38, \5316 );
nor \U$46241 ( \46584 , \46582 , \46583 );
and \U$46242 ( \46585 , \46584 , \5322 );
not \U$46243 ( \46586 , \46584 );
and \U$46244 ( \46587 , \46586 , \5052 );
nor \U$46245 ( \46588 , \46585 , \46587 );
and \U$46246 ( \46589 , \5881 , RI986ec38_34);
and \U$46247 ( \46590 , RI986ed28_36, \5879 );
nor \U$46248 ( \46591 , \46589 , \46590 );
and \U$46249 ( \46592 , \46591 , \5885 );
not \U$46250 ( \46593 , \46591 );
and \U$46251 ( \46594 , \46593 , \5594 );
nor \U$46252 ( \46595 , \46592 , \46594 );
or \U$46253 ( \46596 , \46588 , \46595 );
not \U$46254 ( \46597 , \46595 );
not \U$46255 ( \46598 , \46588 );
or \U$46256 ( \46599 , \46597 , \46598 );
and \U$46257 ( \46600 , \6453 , RI986f0e8_44);
and \U$46258 ( \46601 , RI986eff8_42, \6451 );
nor \U$46259 ( \46602 , \46600 , \46601 );
and \U$46260 ( \46603 , \46602 , \6190 );
not \U$46261 ( \46604 , \46602 );
and \U$46262 ( \46605 , \46604 , \6180 );
nor \U$46263 ( \46606 , \46603 , \46605 );
nand \U$46264 ( \46607 , \46599 , \46606 );
nand \U$46265 ( \46608 , \46596 , \46607 );
and \U$46266 ( \46609 , \46581 , \46608 );
and \U$46267 ( \46610 , \46553 , \46580 );
or \U$46268 ( \46611 , \46609 , \46610 );
and \U$46269 ( \46612 , \9237 , RI986f868_60);
and \U$46270 ( \46613 , RI986f778_58, \9235 );
nor \U$46271 ( \46614 , \46612 , \46613 );
and \U$46272 ( \46615 , \46614 , \8836 );
not \U$46273 ( \46616 , \46614 );
and \U$46274 ( \46617 , \46616 , \9241 );
nor \U$46275 ( \46618 , \46615 , \46617 );
and \U$46276 ( \46619 , \9505 , RI986fa48_64);
and \U$46277 ( \46620 , RI986f958_62, \9503 );
nor \U$46278 ( \46621 , \46619 , \46620 );
and \U$46279 ( \46622 , \46621 , \9513 );
not \U$46280 ( \46623 , \46621 );
and \U$46281 ( \46624 , \46623 , \9510 );
nor \U$46282 ( \46625 , \46622 , \46624 );
xor \U$46283 ( \46626 , \46618 , \46625 );
and \U$46284 ( \46627 , \10424 , RI986f4a8_52);
and \U$46285 ( \46628 , RI986f3b8_50, \10422 );
nor \U$46286 ( \46629 , \46627 , \46628 );
and \U$46287 ( \46630 , \46629 , \10428 );
not \U$46288 ( \46631 , \46629 );
and \U$46289 ( \46632 , \46631 , \9840 );
nor \U$46290 ( \46633 , \46630 , \46632 );
and \U$46291 ( \46634 , \46626 , \46633 );
and \U$46292 ( \46635 , \46618 , \46625 );
or \U$46293 ( \46636 , \46634 , \46635 );
and \U$46294 ( \46637 , \14937 , RI986e2d8_14);
and \U$46295 ( \46638 , RI986e3c8_16, \14935 );
nor \U$46296 ( \46639 , \46637 , \46638 );
and \U$46297 ( \46640 , \46639 , \14538 );
not \U$46298 ( \46641 , \46639 );
and \U$46299 ( \46642 , \46641 , \14539 );
nor \U$46300 ( \46643 , \46640 , \46642 );
xor \U$46301 ( \46644 , \46643 , RI9873558_190);
and \U$46302 ( \46645 , \13882 , RI986e1e8_12);
and \U$46303 ( \46646 , RI986e0f8_10, \13880 );
nor \U$46304 ( \46647 , \46645 , \46646 );
and \U$46305 ( \46648 , \46647 , \13359 );
not \U$46306 ( \46649 , \46647 );
and \U$46307 ( \46650 , \46649 , \13358 );
nor \U$46308 ( \46651 , \46648 , \46650 );
and \U$46309 ( \46652 , \46644 , \46651 );
and \U$46310 ( \46653 , \46643 , RI9873558_190);
or \U$46311 ( \46654 , \46652 , \46653 );
or \U$46312 ( \46655 , \46636 , \46654 );
not \U$46313 ( \46656 , \46654 );
not \U$46314 ( \46657 , \46636 );
or \U$46315 ( \46658 , \46656 , \46657 );
and \U$46316 ( \46659 , \13045 , RI986de28_4);
and \U$46317 ( \46660 , RI986dd38_2, \13043 );
nor \U$46318 ( \46661 , \46659 , \46660 );
and \U$46319 ( \46662 , \46661 , \13047 );
not \U$46320 ( \46663 , \46661 );
and \U$46321 ( \46664 , \46663 , \12619 );
nor \U$46322 ( \46665 , \46662 , \46664 );
and \U$46323 ( \46666 , \11696 , RI986f598_54);
and \U$46324 ( \46667 , RI986f688_56, \11694 );
nor \U$46325 ( \46668 , \46666 , \46667 );
and \U$46326 ( \46669 , \46668 , \10965 );
not \U$46327 ( \46670 , \46668 );
and \U$46328 ( \46671 , \46670 , \11702 );
nor \U$46329 ( \46672 , \46669 , \46671 );
xor \U$46330 ( \46673 , \46665 , \46672 );
and \U$46331 ( \46674 , \12293 , RI986e008_8);
and \U$46332 ( \46675 , RI986df18_6, \12291 );
nor \U$46333 ( \46676 , \46674 , \46675 );
and \U$46334 ( \46677 , \46676 , \11687 );
not \U$46335 ( \46678 , \46676 );
and \U$46336 ( \46679 , \46678 , \11686 );
nor \U$46337 ( \46680 , \46677 , \46679 );
and \U$46338 ( \46681 , \46673 , \46680 );
and \U$46339 ( \46682 , \46665 , \46672 );
or \U$46340 ( \46683 , \46681 , \46682 );
nand \U$46341 ( \46684 , \46658 , \46683 );
nand \U$46342 ( \46685 , \46655 , \46684 );
xor \U$46343 ( \46686 , \46611 , \46685 );
and \U$46344 ( \46687 , \2464 , RI9871398_118);
and \U$46345 ( \46688 , RI9871488_120, \2462 );
nor \U$46346 ( \46689 , \46687 , \46688 );
and \U$46347 ( \46690 , \46689 , \2263 );
not \U$46348 ( \46691 , \46689 );
and \U$46349 ( \46692 , \46691 , \2468 );
nor \U$46350 ( \46693 , \46690 , \46692 );
and \U$46351 ( \46694 , \3254 , RI9871758_126);
and \U$46352 ( \46695 , RI9871848_128, \3252 );
nor \U$46353 ( \46696 , \46694 , \46695 );
not \U$46354 ( \46697 , \46696 );
not \U$46355 ( \46698 , \2935 );
and \U$46356 ( \46699 , \46697 , \46698 );
and \U$46357 ( \46700 , \46696 , \2935 );
nor \U$46358 ( \46701 , \46699 , \46700 );
xor \U$46359 ( \46702 , \46693 , \46701 );
and \U$46360 ( \46703 , \2274 , RI98712a8_116);
and \U$46361 ( \46704 , RI98711b8_114, \2272 );
nor \U$46362 ( \46705 , \46703 , \46704 );
and \U$46363 ( \46706 , \46705 , \2031 );
not \U$46364 ( \46707 , \46705 );
and \U$46365 ( \46708 , \46707 , \2030 );
nor \U$46366 ( \46709 , \46706 , \46708 );
and \U$46367 ( \46710 , \46702 , \46709 );
and \U$46368 ( \46711 , \46693 , \46701 );
nor \U$46369 ( \46712 , \46710 , \46711 );
and \U$46370 ( \46713 , \1311 , RI9870ee8_108);
and \U$46371 ( \46714 , RI9870c18_102, \1309 );
nor \U$46372 ( \46715 , \46713 , \46714 );
and \U$46373 ( \46716 , \46715 , \1315 );
not \U$46374 ( \46717 , \46715 );
and \U$46375 ( \46718 , \46717 , \1319 );
nor \U$46376 ( \46719 , \46716 , \46718 );
and \U$46377 ( \46720 , \2042 , RI98710c8_112);
and \U$46378 ( \46721 , RI9870d08_104, \2040 );
nor \U$46379 ( \46722 , \46720 , \46721 );
not \U$46380 ( \46723 , \46722 );
not \U$46381 ( \46724 , \1462 );
and \U$46382 ( \46725 , \46723 , \46724 );
and \U$46383 ( \46726 , \46722 , \1462 );
nor \U$46384 ( \46727 , \46725 , \46726 );
xor \U$46385 ( \46728 , \46719 , \46727 );
and \U$46386 ( \46729 , \1329 , RI9870df8_106);
and \U$46387 ( \46730 , RI9870a38_98, \1327 );
nor \U$46388 ( \46731 , \46729 , \46730 );
and \U$46389 ( \46732 , \46731 , \1337 );
not \U$46390 ( \46733 , \46731 );
and \U$46391 ( \46734 , \46733 , \1336 );
nor \U$46392 ( \46735 , \46732 , \46734 );
and \U$46393 ( \46736 , \46728 , \46735 );
and \U$46394 ( \46737 , \46719 , \46727 );
nor \U$46395 ( \46738 , \46736 , \46737 );
xor \U$46396 ( \46739 , \46712 , \46738 );
and \U$46397 ( \46740 , \776 , RI98700d8_78);
and \U$46398 ( \46741 , RI98701c8_80, \774 );
nor \U$46399 ( \46742 , \46740 , \46741 );
and \U$46400 ( \46743 , \46742 , \474 );
not \U$46401 ( \46744 , \46742 );
and \U$46402 ( \46745 , \46744 , \451 );
nor \U$46403 ( \46746 , \46743 , \46745 );
and \U$46404 ( \46747 , \438 , RI986ffe8_76);
and \U$46405 ( \46748 , RI986fef8_74, \436 );
nor \U$46406 ( \46749 , \46747 , \46748 );
and \U$46407 ( \46750 , \46749 , \444 );
not \U$46408 ( \46751 , \46749 );
and \U$46409 ( \46752 , \46751 , \443 );
nor \U$46410 ( \46753 , \46750 , \46752 );
xor \U$46411 ( \46754 , \46746 , \46753 );
not \U$46412 ( \46755 , \1301 );
and \U$46413 ( \46756 , \1293 , RI9870fd8_110);
and \U$46414 ( \46757 , RI9870b28_100, \1291 );
nor \U$46415 ( \46758 , \46756 , \46757 );
not \U$46416 ( \46759 , \46758 );
or \U$46417 ( \46760 , \46755 , \46759 );
or \U$46418 ( \46761 , \46758 , \1128 );
nand \U$46419 ( \46762 , \46760 , \46761 );
and \U$46420 ( \46763 , \46754 , \46762 );
and \U$46421 ( \46764 , \46746 , \46753 );
or \U$46422 ( \46765 , \46763 , \46764 );
and \U$46423 ( \46766 , \46739 , \46765 );
and \U$46424 ( \46767 , \46712 , \46738 );
or \U$46425 ( \46768 , \46766 , \46767 );
and \U$46426 ( \46769 , \46686 , \46768 );
and \U$46427 ( \46770 , \46611 , \46685 );
or \U$46428 ( \46771 , \46769 , \46770 );
xor \U$46429 ( \46772 , \46526 , \46771 );
xor \U$46430 ( \46773 , \46375 , \46382 );
xor \U$46431 ( \46774 , \46773 , \46390 );
xor \U$46432 ( \46775 , \46215 , \46222 );
xor \U$46433 ( \46776 , \46775 , \46230 );
xor \U$46434 ( \46777 , \46774 , \46776 );
xor \U$46435 ( \46778 , \46241 , \46248 );
xor \U$46436 ( \46779 , \46778 , \46256 );
and \U$46437 ( \46780 , \46777 , \46779 );
and \U$46438 ( \46781 , \46774 , \46776 );
nor \U$46439 ( \46782 , \46780 , \46781 );
xor \U$46440 ( \46783 , \46143 , \46145 );
xor \U$46441 ( \46784 , \46782 , \46783 );
xor \U$46442 ( \46785 , \45833 , \45840 );
xor \U$46443 ( \46786 , \46785 , \45848 );
xor \U$46444 ( \46787 , \46131 , \46136 );
xor \U$46445 ( \46788 , \46786 , \46787 );
and \U$46446 ( \46789 , \46784 , \46788 );
and \U$46447 ( \46790 , \46782 , \46783 );
or \U$46448 ( \46791 , \46789 , \46790 );
and \U$46449 ( \46792 , \46772 , \46791 );
and \U$46450 ( \46793 , \46526 , \46771 );
nor \U$46451 ( \46794 , \46792 , \46793 );
not \U$46452 ( \46795 , \46794 );
nand \U$46453 ( \46796 , \46439 , \46795 );
nand \U$46454 ( \46797 , \46438 , \46796 );
xor \U$46455 ( \46798 , \45658 , \45660 );
xor \U$46456 ( \46799 , \46798 , \45675 );
xor \U$46457 ( \46800 , \46797 , \46799 );
xor \U$46458 ( \46801 , \45782 , \45854 );
xor \U$46459 ( \46802 , \46801 , \45937 );
xor \U$46460 ( \46803 , \45990 , \45992 );
xor \U$46461 ( \46804 , \46803 , \45995 );
and \U$46462 ( \46805 , \46157 , \46804 );
xor \U$46463 ( \46806 , \45990 , \45992 );
xor \U$46464 ( \46807 , \46806 , \45995 );
and \U$46465 ( \46808 , \46161 , \46807 );
and \U$46466 ( \46809 , \46157 , \46161 );
or \U$46467 ( \46810 , \46805 , \46808 , \46809 );
xor \U$46468 ( \46811 , \45807 , \45825 );
xor \U$46469 ( \46812 , \46811 , \45851 );
and \U$46470 ( \46813 , \46429 , \46812 );
xor \U$46471 ( \46814 , \45807 , \45825 );
xor \U$46472 ( \46815 , \46814 , \45851 );
and \U$46473 ( \46816 , \46431 , \46815 );
and \U$46474 ( \46817 , \46429 , \46431 );
or \U$46475 ( \46818 , \46813 , \46816 , \46817 );
xor \U$46476 ( \46819 , \46810 , \46818 );
xor \U$46477 ( \46820 , \45402 , \45428 );
xor \U$46478 ( \46821 , \46820 , \45456 );
xor \U$46479 ( \46822 , \45648 , \45653 );
xor \U$46480 ( \46823 , \46821 , \46822 );
xor \U$46481 ( \46824 , \46819 , \46823 );
and \U$46482 ( \46825 , \46802 , \46824 );
xor \U$46483 ( \46826 , \45953 , \45987 );
xor \U$46484 ( \46827 , \46826 , \45998 );
xor \U$46485 ( \46828 , \45690 , \45692 );
xor \U$46486 ( \46829 , \46828 , \45697 );
xor \U$46487 ( \46830 , \45283 , \45285 );
xor \U$46488 ( \46831 , \46830 , \45288 );
xor \U$46489 ( \46832 , \45663 , \45670 );
xor \U$46490 ( \46833 , \46831 , \46832 );
xor \U$46491 ( \46834 , \46829 , \46833 );
xor \U$46492 ( \46835 , \46827 , \46834 );
xor \U$46493 ( \46836 , \46810 , \46818 );
xor \U$46494 ( \46837 , \46836 , \46823 );
and \U$46495 ( \46838 , \46835 , \46837 );
and \U$46496 ( \46839 , \46802 , \46835 );
or \U$46497 ( \46840 , \46825 , \46838 , \46839 );
xor \U$46498 ( \46841 , \46800 , \46840 );
xor \U$46499 ( \46842 , \46260 , \46340 );
xor \U$46500 ( \46843 , \46842 , \46421 );
not \U$46501 ( \46844 , \46843 );
xor \U$46502 ( \46845 , \46553 , \46580 );
xor \U$46503 ( \46846 , \46845 , \46608 );
xor \U$46504 ( \46847 , \46712 , \46738 );
xor \U$46505 ( \46848 , \46847 , \46765 );
and \U$46506 ( \46849 , \46846 , \46848 );
xor \U$46507 ( \46850 , \46478 , \46480 );
xor \U$46508 ( \46851 , \46850 , \46509 );
xor \U$46509 ( \46852 , \46712 , \46738 );
xor \U$46510 ( \46853 , \46852 , \46765 );
and \U$46511 ( \46854 , \46851 , \46853 );
and \U$46512 ( \46855 , \46846 , \46851 );
or \U$46513 ( \46856 , \46849 , \46854 , \46855 );
not \U$46514 ( \46857 , \46856 );
not \U$46515 ( \46858 , \46857 );
and \U$46516 ( \46859 , \46844 , \46858 );
and \U$46517 ( \46860 , \46843 , \46857 );
xor \U$46518 ( \46861 , \46449 , \46451 );
xor \U$46519 ( \46862 , \46861 , \46454 );
not \U$46520 ( \46863 , \46862 );
xor \U$46521 ( \46864 , \46774 , \46776 );
xor \U$46522 ( \46865 , \46864 , \46779 );
not \U$46523 ( \46866 , \46865 );
and \U$46524 ( \46867 , \46863 , \46866 );
and \U$46525 ( \46868 , \46862 , \46865 );
xor \U$46526 ( \46869 , \46515 , \46517 );
xor \U$46527 ( \46870 , \46869 , \46520 );
nor \U$46528 ( \46871 , \46868 , \46870 );
nor \U$46529 ( \46872 , \46867 , \46871 );
nor \U$46530 ( \46873 , \46860 , \46872 );
nor \U$46531 ( \46874 , \46859 , \46873 );
and \U$46532 ( \46875 , \1311 , RI9870a38_98);
and \U$46533 ( \46876 , RI9870ee8_108, \1309 );
nor \U$46534 ( \46877 , \46875 , \46876 );
and \U$46535 ( \46878 , \46877 , \1315 );
not \U$46536 ( \46879 , \46877 );
and \U$46537 ( \46880 , \46879 , \1458 );
nor \U$46538 ( \46881 , \46878 , \46880 );
and \U$46539 ( \46882 , \2042 , RI9870c18_102);
and \U$46540 ( \46883 , RI98710c8_112, \2040 );
nor \U$46541 ( \46884 , \46882 , \46883 );
not \U$46542 ( \46885 , \46884 );
not \U$46543 ( \46886 , \2034 );
and \U$46544 ( \46887 , \46885 , \46886 );
and \U$46545 ( \46888 , \46884 , \2034 );
nor \U$46546 ( \46889 , \46887 , \46888 );
xor \U$46547 ( \46890 , \46881 , \46889 );
and \U$46548 ( \46891 , \2274 , RI9870d08_104);
and \U$46549 ( \46892 , RI98712a8_116, \2272 );
nor \U$46550 ( \46893 , \46891 , \46892 );
and \U$46551 ( \46894 , \46893 , \2031 );
not \U$46552 ( \46895 , \46893 );
and \U$46553 ( \46896 , \46895 , \2030 );
nor \U$46554 ( \46897 , \46894 , \46896 );
and \U$46555 ( \46898 , \46890 , \46897 );
and \U$46556 ( \46899 , \46881 , \46889 );
or \U$46557 ( \46900 , \46898 , \46899 );
and \U$46558 ( \46901 , \2464 , RI98711b8_114);
and \U$46559 ( \46902 , RI9871398_118, \2462 );
nor \U$46560 ( \46903 , \46901 , \46902 );
and \U$46561 ( \46904 , \46903 , \2263 );
not \U$46562 ( \46905 , \46903 );
and \U$46563 ( \46906 , \46905 , \2468 );
nor \U$46564 ( \46907 , \46904 , \46906 );
and \U$46565 ( \46908 , \3254 , RI9871488_120);
and \U$46566 ( \46909 , RI9871758_126, \3252 );
nor \U$46567 ( \46910 , \46908 , \46909 );
not \U$46568 ( \46911 , \46910 );
not \U$46569 ( \46912 , \2935 );
and \U$46570 ( \46913 , \46911 , \46912 );
and \U$46571 ( \46914 , \46910 , \3406 );
nor \U$46572 ( \46915 , \46913 , \46914 );
xor \U$46573 ( \46916 , \46907 , \46915 );
and \U$46574 ( \46917 , \3683 , RI9871848_128);
and \U$46575 ( \46918 , RI9871578_122, \3681 );
nor \U$46576 ( \46919 , \46917 , \46918 );
not \U$46577 ( \46920 , \46919 );
not \U$46578 ( \46921 , \3918 );
and \U$46579 ( \46922 , \46920 , \46921 );
and \U$46580 ( \46923 , \46919 , \3918 );
nor \U$46581 ( \46924 , \46922 , \46923 );
and \U$46582 ( \46925 , \46916 , \46924 );
and \U$46583 ( \46926 , \46907 , \46915 );
or \U$46584 ( \46927 , \46925 , \46926 );
or \U$46585 ( \46928 , \46900 , \46927 );
not \U$46586 ( \46929 , \46900 );
not \U$46587 ( \46930 , \46927 );
or \U$46588 ( \46931 , \46929 , \46930 );
and \U$46589 ( \46932 , \1293 , RI98701c8_80);
and \U$46590 ( \46933 , RI9870fd8_110, \1291 );
nor \U$46591 ( \46934 , \46932 , \46933 );
not \U$46592 ( \46935 , \46934 );
not \U$46593 ( \46936 , \1128 );
and \U$46594 ( \46937 , \46935 , \46936 );
and \U$46595 ( \46938 , \46934 , \1128 );
nor \U$46596 ( \46939 , \46937 , \46938 );
and \U$46597 ( \46940 , \1329 , RI9870b28_100);
and \U$46598 ( \46941 , RI9870df8_106, \1327 );
nor \U$46599 ( \46942 , \46940 , \46941 );
and \U$46600 ( \46943 , \46942 , \1337 );
not \U$46601 ( \46944 , \46942 );
and \U$46602 ( \46945 , \46944 , \1336 );
nor \U$46603 ( \46946 , \46943 , \46945 );
xor \U$46604 ( \46947 , \46939 , \46946 );
and \U$46605 ( \46948 , \776 , RI986fef8_74);
and \U$46606 ( \46949 , RI98700d8_78, \774 );
nor \U$46607 ( \46950 , \46948 , \46949 );
and \U$46608 ( \46951 , \46950 , \451 );
not \U$46609 ( \46952 , \46950 );
and \U$46610 ( \46953 , \46952 , \474 );
nor \U$46611 ( \46954 , \46951 , \46953 );
and \U$46612 ( \46955 , \46947 , \46954 );
and \U$46613 ( \46956 , \46939 , \46946 );
nor \U$46614 ( \46957 , \46955 , \46956 );
nand \U$46615 ( \46958 , \46931 , \46957 );
nand \U$46616 ( \46959 , \46928 , \46958 );
and \U$46617 ( \46960 , \7079 , RI986eff8_42);
and \U$46618 ( \46961 , RI986f2c8_48, \7077 );
nor \U$46619 ( \46962 , \46960 , \46961 );
and \U$46620 ( \46963 , \46962 , \6709 );
not \U$46621 ( \46964 , \46962 );
and \U$46622 ( \46965 , \46964 , \6710 );
nor \U$46623 ( \46966 , \46963 , \46965 );
and \U$46624 ( \46967 , \5881 , RI986ee18_38);
and \U$46625 ( \46968 , RI986ec38_34, \5879 );
nor \U$46626 ( \46969 , \46967 , \46968 );
and \U$46627 ( \46970 , \46969 , \5885 );
not \U$46628 ( \46971 , \46969 );
and \U$46629 ( \46972 , \46971 , \5594 );
nor \U$46630 ( \46973 , \46970 , \46972 );
xor \U$46631 ( \46974 , \46966 , \46973 );
and \U$46632 ( \46975 , \6453 , RI986ed28_36);
and \U$46633 ( \46976 , RI986f0e8_44, \6451 );
nor \U$46634 ( \46977 , \46975 , \46976 );
and \U$46635 ( \46978 , \46977 , \6180 );
not \U$46636 ( \46979 , \46977 );
and \U$46637 ( \46980 , \46979 , \6190 );
nor \U$46638 ( \46981 , \46978 , \46980 );
and \U$46639 ( \46982 , \46974 , \46981 );
and \U$46640 ( \46983 , \46966 , \46973 );
or \U$46641 ( \46984 , \46982 , \46983 );
and \U$46642 ( \46985 , \9237 , RI986e698_22);
and \U$46643 ( \46986 , RI986f868_60, \9235 );
nor \U$46644 ( \46987 , \46985 , \46986 );
and \U$46645 ( \46988 , \46987 , \8836 );
not \U$46646 ( \46989 , \46987 );
and \U$46647 ( \46990 , \46989 , \9241 );
nor \U$46648 ( \46991 , \46988 , \46990 );
and \U$46649 ( \46992 , \7729 , RI986f1d8_46);
and \U$46650 ( \46993 , RI986e5a8_20, \7727 );
nor \U$46651 ( \46994 , \46992 , \46993 );
and \U$46652 ( \46995 , \46994 , \7733 );
not \U$46653 ( \46996 , \46994 );
and \U$46654 ( \46997 , \46996 , \7480 );
nor \U$46655 ( \46998 , \46995 , \46997 );
xor \U$46656 ( \46999 , \46991 , \46998 );
and \U$46657 ( \47000 , \8486 , RI986e4b8_18);
and \U$46658 ( \47001 , RI986e788_24, \8484 );
nor \U$46659 ( \47002 , \47000 , \47001 );
and \U$46660 ( \47003 , \47002 , \8051 );
not \U$46661 ( \47004 , \47002 );
and \U$46662 ( \47005 , \47004 , \8050 );
nor \U$46663 ( \47006 , \47003 , \47005 );
and \U$46664 ( \47007 , \46999 , \47006 );
and \U$46665 ( \47008 , \46991 , \46998 );
or \U$46666 ( \47009 , \47007 , \47008 );
or \U$46667 ( \47010 , \46984 , \47009 );
not \U$46668 ( \47011 , \46984 );
not \U$46669 ( \47012 , \47009 );
or \U$46670 ( \47013 , \47011 , \47012 );
and \U$46671 ( \47014 , \4203 , RI9871668_124);
and \U$46672 ( \47015 , RI986eb48_32, \4201 );
nor \U$46673 ( \47016 , \47014 , \47015 );
and \U$46674 ( \47017 , \47016 , \3923 );
not \U$46675 ( \47018 , \47016 );
and \U$46676 ( \47019 , \47018 , \4207 );
nor \U$46677 ( \47020 , \47017 , \47019 );
and \U$46678 ( \47021 , \4710 , RI986ea58_30);
and \U$46679 ( \47022 , RI986e968_28, \4708 );
nor \U$46680 ( \47023 , \47021 , \47022 );
not \U$46681 ( \47024 , \47023 );
not \U$46682 ( \47025 , \4521 );
and \U$46683 ( \47026 , \47024 , \47025 );
and \U$46684 ( \47027 , \47023 , \4519 );
nor \U$46685 ( \47028 , \47026 , \47027 );
or \U$46686 ( \47029 , \47020 , \47028 );
not \U$46687 ( \47030 , \47028 );
not \U$46688 ( \47031 , \47020 );
or \U$46689 ( \47032 , \47030 , \47031 );
and \U$46690 ( \47033 , \5318 , RI986e878_26);
and \U$46691 ( \47034 , RI986ef08_40, \5316 );
nor \U$46692 ( \47035 , \47033 , \47034 );
and \U$46693 ( \47036 , \47035 , \5052 );
not \U$46694 ( \47037 , \47035 );
and \U$46695 ( \47038 , \47037 , \5322 );
nor \U$46696 ( \47039 , \47036 , \47038 );
nand \U$46697 ( \47040 , \47032 , \47039 );
nand \U$46698 ( \47041 , \47029 , \47040 );
nand \U$46699 ( \47042 , \47013 , \47041 );
nand \U$46700 ( \47043 , \47010 , \47042 );
and \U$46701 ( \47044 , \46959 , \47043 );
not \U$46702 ( \47045 , \47043 );
not \U$46703 ( \47046 , \46959 );
and \U$46704 ( \47047 , \47045 , \47046 );
and \U$46705 ( \47048 , \13882 , RI986dd38_2);
and \U$46706 ( \47049 , RI986e1e8_12, \13880 );
nor \U$46707 ( \47050 , \47048 , \47049 );
and \U$46708 ( \47051 , \47050 , \13359 );
not \U$46709 ( \47052 , \47050 );
and \U$46710 ( \47053 , \47052 , \13358 );
nor \U$46711 ( \47054 , \47051 , \47053 );
and \U$46712 ( \47055 , \12293 , RI986f688_56);
and \U$46713 ( \47056 , RI986e008_8, \12291 );
nor \U$46714 ( \47057 , \47055 , \47056 );
and \U$46715 ( \47058 , \47057 , \11686 );
not \U$46716 ( \47059 , \47057 );
and \U$46717 ( \47060 , \47059 , \11687 );
nor \U$46718 ( \47061 , \47058 , \47060 );
xor \U$46719 ( \47062 , \47054 , \47061 );
and \U$46720 ( \47063 , \13045 , RI986df18_6);
and \U$46721 ( \47064 , RI986de28_4, \13043 );
nor \U$46722 ( \47065 , \47063 , \47064 );
and \U$46723 ( \47066 , \47065 , \12619 );
not \U$46724 ( \47067 , \47065 );
and \U$46725 ( \47068 , \47067 , \13047 );
nor \U$46726 ( \47069 , \47066 , \47068 );
and \U$46727 ( \47070 , \47062 , \47069 );
and \U$46728 ( \47071 , \47054 , \47061 );
or \U$46729 ( \47072 , \47070 , \47071 );
and \U$46730 ( \47073 , \14937 , RI986e0f8_10);
and \U$46731 ( \47074 , RI986e2d8_14, \14935 );
nor \U$46732 ( \47075 , \47073 , \47074 );
and \U$46733 ( \47076 , \47075 , \14538 );
not \U$46734 ( \47077 , \47075 );
and \U$46735 ( \47078 , \47077 , \14539 );
nor \U$46736 ( \47079 , \47076 , \47078 );
not \U$46737 ( \47080 , \47079 );
and \U$46738 ( \47081 , \15780 , RI986e3c8_16);
nor \U$46739 ( \47082 , \47081 , \14932 );
nand \U$46740 ( \47083 , \47080 , \47082 );
xor \U$46741 ( \47084 , \47072 , \47083 );
and \U$46742 ( \47085 , \11696 , RI986f3b8_50);
and \U$46743 ( \47086 , RI986f598_54, \11694 );
nor \U$46744 ( \47087 , \47085 , \47086 );
and \U$46745 ( \47088 , \47087 , \11702 );
not \U$46746 ( \47089 , \47087 );
and \U$46747 ( \47090 , \47089 , \10965 );
nor \U$46748 ( \47091 , \47088 , \47090 );
and \U$46749 ( \47092 , \9505 , RI986f778_58);
and \U$46750 ( \47093 , RI986fa48_64, \9503 );
nor \U$46751 ( \47094 , \47092 , \47093 );
and \U$46752 ( \47095 , \47094 , \9513 );
not \U$46753 ( \47096 , \47094 );
and \U$46754 ( \47097 , \47096 , \9510 );
nor \U$46755 ( \47098 , \47095 , \47097 );
xor \U$46756 ( \47099 , \47091 , \47098 );
and \U$46757 ( \47100 , \10424 , RI986f958_62);
and \U$46758 ( \47101 , RI986f4a8_52, \10422 );
nor \U$46759 ( \47102 , \47100 , \47101 );
and \U$46760 ( \47103 , \47102 , \10428 );
not \U$46761 ( \47104 , \47102 );
and \U$46762 ( \47105 , \47104 , \9840 );
nor \U$46763 ( \47106 , \47103 , \47105 );
and \U$46764 ( \47107 , \47099 , \47106 );
and \U$46765 ( \47108 , \47091 , \47098 );
or \U$46766 ( \47109 , \47107 , \47108 );
and \U$46767 ( \47110 , \47084 , \47109 );
and \U$46768 ( \47111 , \47072 , \47083 );
or \U$46769 ( \47112 , \47110 , \47111 );
nor \U$46770 ( \47113 , \47047 , \47112 );
nor \U$46771 ( \47114 , \47044 , \47113 );
xor \U$46772 ( \47115 , \46665 , \46672 );
xor \U$46773 ( \47116 , \47115 , \46680 );
not \U$46774 ( \47117 , \47116 );
xor \U$46775 ( \47118 , \46643 , RI9873558_190);
xor \U$46776 ( \47119 , \47118 , \46651 );
nor \U$46777 ( \47120 , \47117 , \47119 );
not \U$46778 ( \47121 , \46190 );
xor \U$46779 ( \47122 , \46206 , \46198 );
not \U$46780 ( \47123 , \47122 );
or \U$46781 ( \47124 , \47121 , \47123 );
or \U$46782 ( \47125 , \47122 , \46190 );
nand \U$46783 ( \47126 , \47124 , \47125 );
and \U$46784 ( \47127 , \47120 , \47126 );
not \U$46785 ( \47128 , \47120 );
not \U$46786 ( \47129 , \47126 );
and \U$46787 ( \47130 , \47128 , \47129 );
not \U$46788 ( \47131 , \46540 );
not \U$46789 ( \47132 , \46551 );
or \U$46790 ( \47133 , \47131 , \47132 );
or \U$46791 ( \47134 , \46540 , \46551 );
nand \U$46792 ( \47135 , \47133 , \47134 );
not \U$46793 ( \47136 , \47135 );
not \U$46794 ( \47137 , \46533 );
and \U$46795 ( \47138 , \47136 , \47137 );
and \U$46796 ( \47139 , \47135 , \46533 );
nor \U$46797 ( \47140 , \47138 , \47139 );
not \U$46798 ( \47141 , \46595 );
not \U$46799 ( \47142 , \46606 );
or \U$46800 ( \47143 , \47141 , \47142 );
or \U$46801 ( \47144 , \46595 , \46606 );
nand \U$46802 ( \47145 , \47143 , \47144 );
not \U$46803 ( \47146 , \47145 );
not \U$46804 ( \47147 , \46588 );
and \U$46805 ( \47148 , \47146 , \47147 );
and \U$46806 ( \47149 , \47145 , \46588 );
nor \U$46807 ( \47150 , \47148 , \47149 );
xor \U$46808 ( \47151 , \47140 , \47150 );
xor \U$46809 ( \47152 , \46618 , \46625 );
xor \U$46810 ( \47153 , \47152 , \46633 );
and \U$46811 ( \47154 , \47151 , \47153 );
and \U$46812 ( \47155 , \47140 , \47150 );
or \U$46813 ( \47156 , \47154 , \47155 );
nor \U$46814 ( \47157 , \47130 , \47156 );
nor \U$46815 ( \47158 , \47127 , \47157 );
xor \U$46816 ( \47159 , \47114 , \47158 );
xor \U$46817 ( \47160 , \46489 , \46497 );
xor \U$46818 ( \47161 , \47160 , \46506 );
xor \U$46819 ( \47162 , \46464 , \46466 );
xor \U$46820 ( \47163 , \47162 , \46475 );
xor \U$46821 ( \47164 , \47161 , \47163 );
xor \U$46822 ( \47165 , \46746 , \46753 );
xor \U$46823 ( \47166 , \47165 , \46762 );
and \U$46824 ( \47167 , \47164 , \47166 );
and \U$46825 ( \47168 , \47161 , \47163 );
nor \U$46826 ( \47169 , \47167 , \47168 );
not \U$46827 ( \47170 , \47169 );
and \U$46828 ( \47171 , \465 , RI986fc28_68);
and \U$46829 ( \47172 , RI986fe08_72, \463 );
nor \U$46830 ( \47173 , \47171 , \47172 );
not \U$46831 ( \47174 , \47173 );
not \U$46832 ( \47175 , \456 );
and \U$46833 ( \47176 , \47174 , \47175 );
and \U$46834 ( \47177 , \47173 , \454 );
nor \U$46835 ( \47178 , \47176 , \47177 );
and \U$46836 ( \47179 , \438 , RI986fd18_70);
and \U$46837 ( \47180 , RI986ffe8_76, \436 );
nor \U$46838 ( \47181 , \47179 , \47180 );
and \U$46839 ( \47182 , \47181 , \443 );
not \U$46840 ( \47183 , \47181 );
and \U$46841 ( \47184 , \47183 , \444 );
nor \U$46842 ( \47185 , \47182 , \47184 );
xor \U$46843 ( \47186 , \47178 , \47185 );
and \U$46844 ( \47187 , \376 , RI9870858_94);
and \U$46845 ( \47188 , RI986fb38_66, \374 );
nor \U$46846 ( \47189 , \47187 , \47188 );
not \U$46847 ( \47190 , \47189 );
not \U$46848 ( \47191 , \367 );
and \U$46849 ( \47192 , \47190 , \47191 );
and \U$46850 ( \47193 , \47189 , \365 );
nor \U$46851 ( \47194 , \47192 , \47193 );
and \U$46852 ( \47195 , \47186 , \47194 );
and \U$46853 ( \47196 , \47178 , \47185 );
nor \U$46854 ( \47197 , \47195 , \47196 );
and \U$46855 ( \47198 , \354 , RI98702b8_82);
and \U$46856 ( \47199 , RI9870768_92, \352 );
nor \U$46857 ( \47200 , \47198 , \47199 );
not \U$46858 ( \47201 , \47200 );
not \U$46859 ( \47202 , \345 );
and \U$46860 ( \47203 , \47201 , \47202 );
and \U$46861 ( \47204 , \47200 , \361 );
nor \U$46862 ( \47205 , \47203 , \47204 );
and \U$46863 ( \47206 , \416 , RI9870588_88);
and \U$46864 ( \47207 , RI98703a8_84, \414 );
nor \U$46865 ( \47208 , \47206 , \47207 );
and \U$46866 ( \47209 , \47208 , \421 );
not \U$46867 ( \47210 , \47208 );
and \U$46868 ( \47211 , \47210 , \422 );
nor \U$46869 ( \47212 , \47209 , \47211 );
or \U$46870 ( \47213 , \47205 , \47212 );
not \U$46871 ( \47214 , \47212 );
not \U$46872 ( \47215 , \47205 );
or \U$46873 ( \47216 , \47214 , \47215 );
not \U$46874 ( \47217 , \386 );
and \U$46875 ( \47218 , \395 , RI9870678_90);
and \U$46876 ( \47219 , RI9870948_96, \393 );
nor \U$46877 ( \47220 , \47218 , \47219 );
not \U$46878 ( \47221 , \47220 );
or \U$46879 ( \47222 , \47217 , \47221 );
or \U$46880 ( \47223 , \47220 , \386 );
nand \U$46881 ( \47224 , \47222 , \47223 );
nand \U$46882 ( \47225 , \47216 , \47224 );
nand \U$46883 ( \47226 , \47213 , \47225 );
nor \U$46884 ( \47227 , \47197 , \47226 );
not \U$46885 ( \47228 , \47227 );
and \U$46886 ( \47229 , \47170 , \47228 );
and \U$46887 ( \47230 , \47169 , \47227 );
xor \U$46888 ( \47231 , \46719 , \46727 );
xor \U$46889 ( \47232 , \47231 , \46735 );
xor \U$46890 ( \47233 , \46693 , \46701 );
xor \U$46891 ( \47234 , \47233 , \46709 );
xor \U$46892 ( \47235 , \47232 , \47234 );
xor \U$46893 ( \47236 , \46560 , \46568 );
xor \U$46894 ( \47237 , \47236 , \46577 );
and \U$46895 ( \47238 , \47235 , \47237 );
and \U$46896 ( \47239 , \47232 , \47234 );
or \U$46897 ( \47240 , \47238 , \47239 );
nor \U$46898 ( \47241 , \47230 , \47240 );
nor \U$46899 ( \47242 , \47229 , \47241 );
and \U$46900 ( \47243 , \47159 , \47242 );
and \U$46901 ( \47244 , \47114 , \47158 );
or \U$46902 ( \47245 , \47243 , \47244 );
or \U$46903 ( \47246 , \46874 , \47245 );
not \U$46904 ( \47247 , \47245 );
not \U$46905 ( \47248 , \46874 );
or \U$46906 ( \47249 , \47247 , \47248 );
xor \U$46907 ( \47250 , \46457 , \46512 );
xor \U$46908 ( \47251 , \47250 , \46523 );
xor \U$46909 ( \47252 , \46782 , \46783 );
xor \U$46910 ( \47253 , \47252 , \46788 );
and \U$46911 ( \47254 , \47251 , \47253 );
xor \U$46912 ( \47255 , \46057 , \46059 );
xor \U$46913 ( \47256 , \47255 , \46062 );
xor \U$46914 ( \47257 , \46171 , \46178 );
xor \U$46915 ( \47258 , \47256 , \47257 );
xor \U$46916 ( \47259 , \46782 , \46783 );
xor \U$46917 ( \47260 , \47259 , \46788 );
and \U$46918 ( \47261 , \47258 , \47260 );
and \U$46919 ( \47262 , \47251 , \47258 );
or \U$46920 ( \47263 , \47254 , \47261 , \47262 );
nand \U$46921 ( \47264 , \47249 , \47263 );
nand \U$46922 ( \47265 , \47246 , \47264 );
xor \U$46923 ( \47266 , \46065 , \46115 );
and \U$46924 ( \47267 , \47266 , \46128 );
and \U$46925 ( \47268 , \46065 , \46115 );
or \U$46926 ( \47269 , \47267 , \47268 );
xor \U$46927 ( \47270 , \46286 , \46312 );
and \U$46928 ( \47271 , \47270 , \46339 );
and \U$46929 ( \47272 , \46286 , \46312 );
nor \U$46930 ( \47273 , \47271 , \47272 );
xor \U$46931 ( \47274 , \46208 , \46233 );
and \U$46932 ( \47275 , \47274 , \46259 );
and \U$46933 ( \47276 , \46208 , \46233 );
nor \U$46934 ( \47277 , \47275 , \47276 );
xor \U$46935 ( \47278 , \47273 , \47277 );
xor \U$46936 ( \47279 , \46368 , \46393 );
and \U$46937 ( \47280 , \47279 , \46420 );
and \U$46938 ( \47281 , \46368 , \46393 );
nor \U$46939 ( \47282 , \47280 , \47281 );
and \U$46940 ( \47283 , \47278 , \47282 );
and \U$46941 ( \47284 , \47273 , \47277 );
or \U$46942 ( \47285 , \47283 , \47284 );
xor \U$46943 ( \47286 , \47269 , \47285 );
xor \U$46944 ( \47287 , \46141 , \46146 );
and \U$46945 ( \47288 , \47287 , \46151 );
and \U$46946 ( \47289 , \46141 , \46146 );
or \U$46947 ( \47290 , \47288 , \47289 );
xor \U$46948 ( \47291 , \47286 , \47290 );
xor \U$46949 ( \47292 , \47265 , \47291 );
xor \U$46950 ( \47293 , \47273 , \47277 );
xor \U$46951 ( \47294 , \47293 , \47282 );
xor \U$46952 ( \47295 , \46183 , \46424 );
xor \U$46953 ( \47296 , \47295 , \46433 );
and \U$46954 ( \47297 , \47294 , \47296 );
xor \U$46955 ( \47298 , \46141 , \46146 );
xor \U$46956 ( \47299 , \47298 , \46151 );
xor \U$46957 ( \47300 , \46129 , \46163 );
xor \U$46958 ( \47301 , \47299 , \47300 );
xor \U$46959 ( \47302 , \46183 , \46424 );
xor \U$46960 ( \47303 , \47302 , \46433 );
and \U$46961 ( \47304 , \47301 , \47303 );
and \U$46962 ( \47305 , \47294 , \47301 );
or \U$46963 ( \47306 , \47297 , \47304 , \47305 );
and \U$46964 ( \47307 , \47292 , \47306 );
and \U$46965 ( \47308 , \47265 , \47291 );
or \U$46966 ( \47309 , \47307 , \47308 );
xor \U$46967 ( \47310 , \45245 , \45280 );
xor \U$46968 ( \47311 , \47310 , \45291 );
xor \U$46969 ( \47312 , \45376 , \45459 );
xor \U$46970 ( \47313 , \47312 , \45537 );
xor \U$46971 ( \47314 , \47311 , \47313 );
xor \U$46972 ( \47315 , \45571 , \45573 );
xor \U$46973 ( \47316 , \47315 , \45578 );
xor \U$46974 ( \47317 , \46007 , \46014 );
xor \U$46975 ( \47318 , \47316 , \47317 );
xor \U$46976 ( \47319 , \47314 , \47318 );
xor \U$46977 ( \47320 , \45700 , \45940 );
xor \U$46978 ( \47321 , \47320 , \46001 );
xor \U$46979 ( \47322 , \46810 , \46818 );
and \U$46980 ( \47323 , \47322 , \46823 );
and \U$46981 ( \47324 , \46810 , \46818 );
or \U$46982 ( \47325 , \47323 , \47324 );
xor \U$46983 ( \47326 , \47269 , \47285 );
and \U$46984 ( \47327 , \47326 , \47290 );
and \U$46985 ( \47328 , \47269 , \47285 );
or \U$46986 ( \47329 , \47327 , \47328 );
xor \U$46987 ( \47330 , \47325 , \47329 );
xor \U$46988 ( \47331 , \45953 , \45987 );
xor \U$46989 ( \47332 , \47331 , \45998 );
and \U$46990 ( \47333 , \46829 , \47332 );
xor \U$46991 ( \47334 , \45953 , \45987 );
xor \U$46992 ( \47335 , \47334 , \45998 );
and \U$46993 ( \47336 , \46833 , \47335 );
and \U$46994 ( \47337 , \46829 , \46833 );
or \U$46995 ( \47338 , \47333 , \47336 , \47337 );
xor \U$46996 ( \47339 , \47330 , \47338 );
xor \U$46997 ( \47340 , \47321 , \47339 );
xor \U$46998 ( \47341 , \47319 , \47340 );
xor \U$46999 ( \47342 , \47309 , \47341 );
xor \U$47000 ( \47343 , \46841 , \47342 );
not \U$47001 ( \47344 , \47343 );
not \U$47002 ( \47345 , \46436 );
not \U$47003 ( \47346 , \46794 );
and \U$47004 ( \47347 , \47345 , \47346 );
and \U$47005 ( \47348 , \46436 , \46794 );
nor \U$47006 ( \47349 , \47347 , \47348 );
not \U$47007 ( \47350 , \47349 );
not \U$47008 ( \47351 , \46168 );
and \U$47009 ( \47352 , \47350 , \47351 );
and \U$47010 ( \47353 , \47349 , \46168 );
nor \U$47011 ( \47354 , \47352 , \47353 );
not \U$47012 ( \47355 , \47354 );
xor \U$47013 ( \47356 , \47265 , \47291 );
xor \U$47014 ( \47357 , \47356 , \47306 );
nand \U$47015 ( \47358 , \47355 , \47357 );
xor \U$47016 ( \47359 , \46810 , \46818 );
xor \U$47017 ( \47360 , \47359 , \46823 );
xor \U$47018 ( \47361 , \46802 , \46835 );
xor \U$47019 ( \47362 , \47360 , \47361 );
not \U$47020 ( \47363 , \47362 );
xnor \U$47021 ( \47364 , \47245 , \46874 );
not \U$47022 ( \47365 , \47364 );
not \U$47023 ( \47366 , \47263 );
and \U$47024 ( \47367 , \47365 , \47366 );
and \U$47025 ( \47368 , \47364 , \47263 );
nor \U$47026 ( \47369 , \47367 , \47368 );
not \U$47027 ( \47370 , \47369 );
xor \U$47028 ( \47371 , \46183 , \46424 );
xor \U$47029 ( \47372 , \47371 , \46433 );
xor \U$47030 ( \47373 , \47294 , \47301 );
xor \U$47031 ( \47374 , \47372 , \47373 );
nand \U$47032 ( \47375 , \47370 , \47374 );
nand \U$47033 ( \47376 , \47363 , \47375 );
not \U$47034 ( \47377 , \46957 );
not \U$47035 ( \47378 , \46900 );
or \U$47036 ( \47379 , \47377 , \47378 );
or \U$47037 ( \47380 , \46900 , \46957 );
nand \U$47038 ( \47381 , \47379 , \47380 );
not \U$47039 ( \47382 , \47381 );
not \U$47040 ( \47383 , \46927 );
and \U$47041 ( \47384 , \47382 , \47383 );
and \U$47042 ( \47385 , \47381 , \46927 );
nor \U$47043 ( \47386 , \47384 , \47385 );
xor \U$47044 ( \47387 , \47072 , \47083 );
xor \U$47045 ( \47388 , \47387 , \47109 );
and \U$47046 ( \47389 , \47386 , \47388 );
not \U$47047 ( \47390 , \47041 );
not \U$47048 ( \47391 , \46984 );
or \U$47049 ( \47392 , \47390 , \47391 );
or \U$47050 ( \47393 , \46984 , \47041 );
nand \U$47051 ( \47394 , \47392 , \47393 );
not \U$47052 ( \47395 , \47394 );
not \U$47053 ( \47396 , \47009 );
and \U$47054 ( \47397 , \47395 , \47396 );
and \U$47055 ( \47398 , \47394 , \47009 );
nor \U$47056 ( \47399 , \47397 , \47398 );
xor \U$47057 ( \47400 , \47072 , \47083 );
xor \U$47058 ( \47401 , \47400 , \47109 );
and \U$47059 ( \47402 , \47399 , \47401 );
and \U$47060 ( \47403 , \47386 , \47399 );
or \U$47061 ( \47404 , \47389 , \47402 , \47403 );
not \U$47062 ( \47405 , \46683 );
not \U$47063 ( \47406 , \46654 );
or \U$47064 ( \47407 , \47405 , \47406 );
or \U$47065 ( \47408 , \46654 , \46683 );
nand \U$47066 ( \47409 , \47407 , \47408 );
not \U$47067 ( \47410 , \47409 );
not \U$47068 ( \47411 , \46636 );
and \U$47069 ( \47412 , \47410 , \47411 );
and \U$47070 ( \47413 , \47409 , \46636 );
nor \U$47071 ( \47414 , \47412 , \47413 );
or \U$47072 ( \47415 , \47404 , \47414 );
not \U$47073 ( \47416 , \47414 );
not \U$47074 ( \47417 , \47404 );
or \U$47075 ( \47418 , \47416 , \47417 );
xor \U$47076 ( \47419 , \47232 , \47234 );
xor \U$47077 ( \47420 , \47419 , \47237 );
and \U$47078 ( \47421 , \47197 , \47226 );
nor \U$47079 ( \47422 , \47421 , \47227 );
or \U$47080 ( \47423 , \47420 , \47422 );
not \U$47081 ( \47424 , \47422 );
not \U$47082 ( \47425 , \47420 );
or \U$47083 ( \47426 , \47424 , \47425 );
xor \U$47084 ( \47427 , \47161 , \47163 );
xor \U$47085 ( \47428 , \47427 , \47166 );
nand \U$47086 ( \47429 , \47426 , \47428 );
nand \U$47087 ( \47430 , \47423 , \47429 );
nand \U$47088 ( \47431 , \47418 , \47430 );
nand \U$47089 ( \47432 , \47415 , \47431 );
and \U$47090 ( \47433 , \7729 , RI986f2c8_48);
and \U$47091 ( \47434 , RI986f1d8_46, \7727 );
nor \U$47092 ( \47435 , \47433 , \47434 );
and \U$47093 ( \47436 , \47435 , \7480 );
not \U$47094 ( \47437 , \47435 );
and \U$47095 ( \47438 , \47437 , \7733 );
nor \U$47096 ( \47439 , \47436 , \47438 );
and \U$47097 ( \47440 , \8486 , RI986e5a8_20);
and \U$47098 ( \47441 , RI986e4b8_18, \8484 );
nor \U$47099 ( \47442 , \47440 , \47441 );
and \U$47100 ( \47443 , \47442 , \8050 );
not \U$47101 ( \47444 , \47442 );
and \U$47102 ( \47445 , \47444 , \8051 );
nor \U$47103 ( \47446 , \47443 , \47445 );
xor \U$47104 ( \47447 , \47439 , \47446 );
and \U$47105 ( \47448 , \7079 , RI986f0e8_44);
and \U$47106 ( \47449 , RI986eff8_42, \7077 );
nor \U$47107 ( \47450 , \47448 , \47449 );
and \U$47108 ( \47451 , \47450 , \6710 );
not \U$47109 ( \47452 , \47450 );
and \U$47110 ( \47453 , \47452 , \6709 );
nor \U$47111 ( \47454 , \47451 , \47453 );
and \U$47112 ( \47455 , \47447 , \47454 );
and \U$47113 ( \47456 , \47439 , \47446 );
nor \U$47114 ( \47457 , \47455 , \47456 );
and \U$47115 ( \47458 , \5318 , RI986e968_28);
and \U$47116 ( \47459 , RI986e878_26, \5316 );
nor \U$47117 ( \47460 , \47458 , \47459 );
and \U$47118 ( \47461 , \47460 , \5322 );
not \U$47119 ( \47462 , \47460 );
and \U$47120 ( \47463 , \47462 , \5052 );
nor \U$47121 ( \47464 , \47461 , \47463 );
not \U$47122 ( \47465 , \47464 );
and \U$47123 ( \47466 , \5881 , RI986ef08_40);
and \U$47124 ( \47467 , RI986ee18_38, \5879 );
nor \U$47125 ( \47468 , \47466 , \47467 );
and \U$47126 ( \47469 , \47468 , \5885 );
not \U$47127 ( \47470 , \47468 );
and \U$47128 ( \47471 , \47470 , \5594 );
nor \U$47129 ( \47472 , \47469 , \47471 );
not \U$47130 ( \47473 , \47472 );
and \U$47131 ( \47474 , \47465 , \47473 );
and \U$47132 ( \47475 , \47472 , \47464 );
and \U$47133 ( \47476 , \6453 , RI986ec38_34);
and \U$47134 ( \47477 , RI986ed28_36, \6451 );
nor \U$47135 ( \47478 , \47476 , \47477 );
and \U$47136 ( \47479 , \47478 , \6180 );
not \U$47137 ( \47480 , \47478 );
and \U$47138 ( \47481 , \47480 , \6190 );
nor \U$47139 ( \47482 , \47479 , \47481 );
nor \U$47140 ( \47483 , \47475 , \47482 );
nor \U$47141 ( \47484 , \47474 , \47483 );
xor \U$47142 ( \47485 , \47457 , \47484 );
and \U$47143 ( \47486 , \4203 , RI9871578_122);
and \U$47144 ( \47487 , RI9871668_124, \4201 );
nor \U$47145 ( \47488 , \47486 , \47487 );
and \U$47146 ( \47489 , \47488 , \4207 );
not \U$47147 ( \47490 , \47488 );
and \U$47148 ( \47491 , \47490 , \3923 );
nor \U$47149 ( \47492 , \47489 , \47491 );
not \U$47150 ( \47493 , \4521 );
and \U$47151 ( \47494 , \4710 , RI986eb48_32);
and \U$47152 ( \47495 , RI986ea58_30, \4708 );
nor \U$47153 ( \47496 , \47494 , \47495 );
not \U$47154 ( \47497 , \47496 );
or \U$47155 ( \47498 , \47493 , \47497 );
or \U$47156 ( \47499 , \47496 , \4521 );
nand \U$47157 ( \47500 , \47498 , \47499 );
xor \U$47158 ( \47501 , \47492 , \47500 );
not \U$47159 ( \47502 , \3412 );
and \U$47160 ( \47503 , \3683 , RI9871758_126);
and \U$47161 ( \47504 , RI9871848_128, \3681 );
nor \U$47162 ( \47505 , \47503 , \47504 );
not \U$47163 ( \47506 , \47505 );
or \U$47164 ( \47507 , \47502 , \47506 );
or \U$47165 ( \47508 , \47505 , \3412 );
nand \U$47166 ( \47509 , \47507 , \47508 );
and \U$47167 ( \47510 , \47501 , \47509 );
and \U$47168 ( \47511 , \47492 , \47500 );
nor \U$47169 ( \47512 , \47510 , \47511 );
and \U$47170 ( \47513 , \47485 , \47512 );
and \U$47171 ( \47514 , \47457 , \47484 );
or \U$47172 ( \47515 , \47513 , \47514 );
and \U$47173 ( \47516 , \2274 , RI98710c8_112);
and \U$47174 ( \47517 , RI9870d08_104, \2272 );
nor \U$47175 ( \47518 , \47516 , \47517 );
and \U$47176 ( \47519 , \47518 , \2031 );
not \U$47177 ( \47520 , \47518 );
and \U$47178 ( \47521 , \47520 , \2030 );
nor \U$47179 ( \47522 , \47519 , \47521 );
not \U$47180 ( \47523 , \47522 );
and \U$47181 ( \47524 , \2464 , RI98712a8_116);
and \U$47182 ( \47525 , RI98711b8_114, \2462 );
nor \U$47183 ( \47526 , \47524 , \47525 );
and \U$47184 ( \47527 , \47526 , \2263 );
not \U$47185 ( \47528 , \47526 );
and \U$47186 ( \47529 , \47528 , \2468 );
nor \U$47187 ( \47530 , \47527 , \47529 );
not \U$47188 ( \47531 , \47530 );
and \U$47189 ( \47532 , \47523 , \47531 );
and \U$47190 ( \47533 , \47530 , \47522 );
and \U$47191 ( \47534 , \3254 , RI9871398_118);
and \U$47192 ( \47535 , RI9871488_120, \3252 );
nor \U$47193 ( \47536 , \47534 , \47535 );
not \U$47194 ( \47537 , \47536 );
not \U$47195 ( \47538 , \2935 );
and \U$47196 ( \47539 , \47537 , \47538 );
and \U$47197 ( \47540 , \47536 , \2935 );
nor \U$47198 ( \47541 , \47539 , \47540 );
nor \U$47199 ( \47542 , \47533 , \47541 );
nor \U$47200 ( \47543 , \47532 , \47542 );
and \U$47201 ( \47544 , \1311 , RI9870df8_106);
and \U$47202 ( \47545 , RI9870a38_98, \1309 );
nor \U$47203 ( \47546 , \47544 , \47545 );
and \U$47204 ( \47547 , \47546 , \1319 );
not \U$47205 ( \47548 , \47546 );
and \U$47206 ( \47549 , \47548 , \1318 );
nor \U$47207 ( \47550 , \47547 , \47549 );
not \U$47208 ( \47551 , \2034 );
and \U$47209 ( \47552 , \2042 , RI9870ee8_108);
and \U$47210 ( \47553 , RI9870c18_102, \2040 );
nor \U$47211 ( \47554 , \47552 , \47553 );
not \U$47212 ( \47555 , \47554 );
or \U$47213 ( \47556 , \47551 , \47555 );
or \U$47214 ( \47557 , \47554 , \1462 );
nand \U$47215 ( \47558 , \47556 , \47557 );
xor \U$47216 ( \47559 , \47550 , \47558 );
and \U$47217 ( \47560 , \1329 , RI9870fd8_110);
and \U$47218 ( \47561 , RI9870b28_100, \1327 );
nor \U$47219 ( \47562 , \47560 , \47561 );
and \U$47220 ( \47563 , \47562 , \1336 );
not \U$47221 ( \47564 , \47562 );
and \U$47222 ( \47565 , \47564 , \1337 );
nor \U$47223 ( \47566 , \47563 , \47565 );
and \U$47224 ( \47567 , \47559 , \47566 );
and \U$47225 ( \47568 , \47550 , \47558 );
nor \U$47226 ( \47569 , \47567 , \47568 );
xor \U$47227 ( \47570 , \47543 , \47569 );
and \U$47228 ( \47571 , \776 , RI986ffe8_76);
and \U$47229 ( \47572 , RI986fef8_74, \774 );
nor \U$47230 ( \47573 , \47571 , \47572 );
and \U$47231 ( \47574 , \47573 , \451 );
not \U$47232 ( \47575 , \47573 );
and \U$47233 ( \47576 , \47575 , \474 );
nor \U$47234 ( \47577 , \47574 , \47576 );
not \U$47235 ( \47578 , \47577 );
and \U$47236 ( \47579 , \438 , RI986fe08_72);
and \U$47237 ( \47580 , RI986fd18_70, \436 );
nor \U$47238 ( \47581 , \47579 , \47580 );
and \U$47239 ( \47582 , \47581 , \443 );
not \U$47240 ( \47583 , \47581 );
and \U$47241 ( \47584 , \47583 , \444 );
nor \U$47242 ( \47585 , \47582 , \47584 );
not \U$47243 ( \47586 , \47585 );
and \U$47244 ( \47587 , \47578 , \47586 );
and \U$47245 ( \47588 , \47585 , \47577 );
and \U$47246 ( \47589 , \1293 , RI98700d8_78);
and \U$47247 ( \47590 , RI98701c8_80, \1291 );
nor \U$47248 ( \47591 , \47589 , \47590 );
not \U$47249 ( \47592 , \47591 );
not \U$47250 ( \47593 , \1301 );
and \U$47251 ( \47594 , \47592 , \47593 );
and \U$47252 ( \47595 , \47591 , \1128 );
nor \U$47253 ( \47596 , \47594 , \47595 );
nor \U$47254 ( \47597 , \47588 , \47596 );
nor \U$47255 ( \47598 , \47587 , \47597 );
and \U$47256 ( \47599 , \47570 , \47598 );
and \U$47257 ( \47600 , \47543 , \47569 );
or \U$47258 ( \47601 , \47599 , \47600 );
xor \U$47259 ( \47602 , \47515 , \47601 );
and \U$47260 ( \47603 , \9237 , RI986e788_24);
and \U$47261 ( \47604 , RI986e698_22, \9235 );
nor \U$47262 ( \47605 , \47603 , \47604 );
and \U$47263 ( \47606 , \47605 , \8836 );
not \U$47264 ( \47607 , \47605 );
and \U$47265 ( \47608 , \47607 , \9241 );
nor \U$47266 ( \47609 , \47606 , \47608 );
not \U$47267 ( \47610 , \47609 );
and \U$47268 ( \47611 , \10424 , RI986fa48_64);
and \U$47269 ( \47612 , RI986f958_62, \10422 );
nor \U$47270 ( \47613 , \47611 , \47612 );
and \U$47271 ( \47614 , \47613 , \10428 );
not \U$47272 ( \47615 , \47613 );
and \U$47273 ( \47616 , \47615 , \9840 );
nor \U$47274 ( \47617 , \47614 , \47616 );
not \U$47275 ( \47618 , \47617 );
and \U$47276 ( \47619 , \47610 , \47618 );
and \U$47277 ( \47620 , \47617 , \47609 );
and \U$47278 ( \47621 , \9505 , RI986f868_60);
and \U$47279 ( \47622 , RI986f778_58, \9503 );
nor \U$47280 ( \47623 , \47621 , \47622 );
and \U$47281 ( \47624 , \47623 , \9513 );
not \U$47282 ( \47625 , \47623 );
and \U$47283 ( \47626 , \47625 , \9510 );
nor \U$47284 ( \47627 , \47624 , \47626 );
nor \U$47285 ( \47628 , \47620 , \47627 );
nor \U$47286 ( \47629 , \47619 , \47628 );
and \U$47287 ( \47630 , \13882 , RI986de28_4);
and \U$47288 ( \47631 , RI986dd38_2, \13880 );
nor \U$47289 ( \47632 , \47630 , \47631 );
and \U$47290 ( \47633 , \47632 , \13359 );
not \U$47291 ( \47634 , \47632 );
and \U$47292 ( \47635 , \47634 , \13358 );
nor \U$47293 ( \47636 , \47633 , \47635 );
and \U$47294 ( \47637 , \15780 , RI986e2d8_14);
and \U$47295 ( \47638 , RI986e3c8_16, RI9873648_192);
nor \U$47296 ( \47639 , \47637 , \47638 );
not \U$47297 ( \47640 , \47639 );
not \U$47298 ( \47641 , RI9873558_190);
and \U$47299 ( \47642 , \47640 , \47641 );
and \U$47300 ( \47643 , \47639 , RI9873558_190);
nor \U$47301 ( \47644 , \47642 , \47643 );
xor \U$47302 ( \47645 , \47636 , \47644 );
and \U$47303 ( \47646 , \14937 , RI986e1e8_12);
and \U$47304 ( \47647 , RI986e0f8_10, \14935 );
nor \U$47305 ( \47648 , \47646 , \47647 );
and \U$47306 ( \47649 , \47648 , \14538 );
nor \U$47307 ( \47650 , \47648 , \14538 );
nor \U$47308 ( \47651 , \47649 , \47650 );
and \U$47309 ( \47652 , \47645 , \47651 );
and \U$47310 ( \47653 , \47636 , \47644 );
or \U$47311 ( \47654 , \47652 , \47653 );
xor \U$47312 ( \47655 , \47629 , \47654 );
and \U$47313 ( \47656 , \11696 , RI986f4a8_52);
and \U$47314 ( \47657 , RI986f3b8_50, \11694 );
nor \U$47315 ( \47658 , \47656 , \47657 );
and \U$47316 ( \47659 , \47658 , \11702 );
not \U$47317 ( \47660 , \47658 );
and \U$47318 ( \47661 , \47660 , \10965 );
nor \U$47319 ( \47662 , \47659 , \47661 );
not \U$47320 ( \47663 , \47662 );
and \U$47321 ( \47664 , \13045 , RI986e008_8);
and \U$47322 ( \47665 , RI986df18_6, \13043 );
nor \U$47323 ( \47666 , \47664 , \47665 );
and \U$47324 ( \47667 , \47666 , \12619 );
not \U$47325 ( \47668 , \47666 );
and \U$47326 ( \47669 , \47668 , \13047 );
nor \U$47327 ( \47670 , \47667 , \47669 );
not \U$47328 ( \47671 , \47670 );
and \U$47329 ( \47672 , \47663 , \47671 );
and \U$47330 ( \47673 , \47670 , \47662 );
and \U$47331 ( \47674 , \12293 , RI986f598_54);
and \U$47332 ( \47675 , RI986f688_56, \12291 );
nor \U$47333 ( \47676 , \47674 , \47675 );
and \U$47334 ( \47677 , \47676 , \11686 );
not \U$47335 ( \47678 , \47676 );
and \U$47336 ( \47679 , \47678 , \11687 );
nor \U$47337 ( \47680 , \47677 , \47679 );
nor \U$47338 ( \47681 , \47673 , \47680 );
nor \U$47339 ( \47682 , \47672 , \47681 );
and \U$47340 ( \47683 , \47655 , \47682 );
and \U$47341 ( \47684 , \47629 , \47654 );
or \U$47342 ( \47685 , \47683 , \47684 );
and \U$47343 ( \47686 , \47602 , \47685 );
and \U$47344 ( \47687 , \47515 , \47601 );
or \U$47345 ( \47688 , \47686 , \47687 );
not \U$47346 ( \47689 , \47028 );
not \U$47347 ( \47690 , \47039 );
or \U$47348 ( \47691 , \47689 , \47690 );
or \U$47349 ( \47692 , \47028 , \47039 );
nand \U$47350 ( \47693 , \47691 , \47692 );
not \U$47351 ( \47694 , \47693 );
not \U$47352 ( \47695 , \47020 );
and \U$47353 ( \47696 , \47694 , \47695 );
and \U$47354 ( \47697 , \47693 , \47020 );
nor \U$47355 ( \47698 , \47696 , \47697 );
xor \U$47356 ( \47699 , \46907 , \46915 );
xor \U$47357 ( \47700 , \47699 , \46924 );
and \U$47358 ( \47701 , \47698 , \47700 );
xor \U$47359 ( \47702 , \46966 , \46973 );
xor \U$47360 ( \47703 , \47702 , \46981 );
xor \U$47361 ( \47704 , \46907 , \46915 );
xor \U$47362 ( \47705 , \47704 , \46924 );
and \U$47363 ( \47706 , \47703 , \47705 );
and \U$47364 ( \47707 , \47698 , \47703 );
or \U$47365 ( \47708 , \47701 , \47706 , \47707 );
and \U$47366 ( \47709 , \376 , RI9870948_96);
and \U$47367 ( \47710 , RI9870858_94, \374 );
nor \U$47368 ( \47711 , \47709 , \47710 );
not \U$47369 ( \47712 , \47711 );
not \U$47370 ( \47713 , \367 );
and \U$47371 ( \47714 , \47712 , \47713 );
and \U$47372 ( \47715 , \47711 , \367 );
nor \U$47373 ( \47716 , \47714 , \47715 );
not \U$47374 ( \47717 , \47716 );
and \U$47375 ( \47718 , \395 , RI9870768_92);
and \U$47376 ( \47719 , RI9870678_90, \393 );
nor \U$47377 ( \47720 , \47718 , \47719 );
not \U$47378 ( \47721 , \47720 );
not \U$47379 ( \47722 , \386 );
and \U$47380 ( \47723 , \47721 , \47722 );
and \U$47381 ( \47724 , \47720 , \487 );
nor \U$47382 ( \47725 , \47723 , \47724 );
not \U$47383 ( \47726 , \47725 );
and \U$47384 ( \47727 , \47717 , \47726 );
and \U$47385 ( \47728 , \47725 , \47716 );
and \U$47386 ( \47729 , \465 , RI986fb38_66);
and \U$47387 ( \47730 , RI986fc28_68, \463 );
nor \U$47388 ( \47731 , \47729 , \47730 );
not \U$47389 ( \47732 , \47731 );
not \U$47390 ( \47733 , \454 );
and \U$47391 ( \47734 , \47732 , \47733 );
and \U$47392 ( \47735 , \47731 , \456 );
nor \U$47393 ( \47736 , \47734 , \47735 );
nor \U$47394 ( \47737 , \47728 , \47736 );
nor \U$47395 ( \47738 , \47727 , \47737 );
nand \U$47396 ( \47739 , RI9870498_86, RI9871fc8_144);
xor \U$47397 ( \47740 , \47738 , \47739 );
not \U$47398 ( \47741 , \47205 );
not \U$47399 ( \47742 , \47224 );
or \U$47400 ( \47743 , \47741 , \47742 );
or \U$47401 ( \47744 , \47205 , \47224 );
nand \U$47402 ( \47745 , \47743 , \47744 );
not \U$47403 ( \47746 , \47745 );
not \U$47404 ( \47747 , \47212 );
and \U$47405 ( \47748 , \47746 , \47747 );
and \U$47406 ( \47749 , \47745 , \47212 );
nor \U$47407 ( \47750 , \47748 , \47749 );
and \U$47408 ( \47751 , \47740 , \47750 );
and \U$47409 ( \47752 , \47738 , \47739 );
or \U$47410 ( \47753 , \47751 , \47752 );
xor \U$47411 ( \47754 , \47708 , \47753 );
xor \U$47412 ( \47755 , \47178 , \47185 );
xor \U$47413 ( \47756 , \47755 , \47194 );
xor \U$47414 ( \47757 , \46939 , \46946 );
xor \U$47415 ( \47758 , \47757 , \46954 );
xor \U$47416 ( \47759 , \47756 , \47758 );
xor \U$47417 ( \47760 , \46881 , \46889 );
xor \U$47418 ( \47761 , \47760 , \46897 );
and \U$47419 ( \47762 , \47759 , \47761 );
and \U$47420 ( \47763 , \47756 , \47758 );
or \U$47421 ( \47764 , \47762 , \47763 );
and \U$47422 ( \47765 , \47754 , \47764 );
and \U$47423 ( \47766 , \47708 , \47753 );
or \U$47424 ( \47767 , \47765 , \47766 );
xor \U$47425 ( \47768 , \47688 , \47767 );
xor \U$47426 ( \47769 , \46991 , \46998 );
xor \U$47427 ( \47770 , \47769 , \47006 );
xor \U$47428 ( \47771 , \47091 , \47098 );
xor \U$47429 ( \47772 , \47771 , \47106 );
and \U$47430 ( \47773 , \47770 , \47772 );
xor \U$47431 ( \47774 , \47054 , \47061 );
xor \U$47432 ( \47775 , \47774 , \47069 );
xor \U$47433 ( \47776 , \47091 , \47098 );
xor \U$47434 ( \47777 , \47776 , \47106 );
and \U$47435 ( \47778 , \47775 , \47777 );
and \U$47436 ( \47779 , \47770 , \47775 );
or \U$47437 ( \47780 , \47773 , \47778 , \47779 );
not \U$47438 ( \47781 , \47119 );
not \U$47439 ( \47782 , \47116 );
and \U$47440 ( \47783 , \47781 , \47782 );
and \U$47441 ( \47784 , \47119 , \47116 );
nor \U$47442 ( \47785 , \47783 , \47784 );
xor \U$47443 ( \47786 , \47780 , \47785 );
xor \U$47444 ( \47787 , \47140 , \47150 );
xor \U$47445 ( \47788 , \47787 , \47153 );
and \U$47446 ( \47789 , \47786 , \47788 );
and \U$47447 ( \47790 , \47780 , \47785 );
or \U$47448 ( \47791 , \47789 , \47790 );
and \U$47449 ( \47792 , \47768 , \47791 );
and \U$47450 ( \47793 , \47688 , \47767 );
nor \U$47451 ( \47794 , \47792 , \47793 );
xor \U$47452 ( \47795 , \47432 , \47794 );
xor \U$47453 ( \47796 , \46712 , \46738 );
xor \U$47454 ( \47797 , \47796 , \46765 );
xor \U$47455 ( \47798 , \46846 , \46851 );
xor \U$47456 ( \47799 , \47797 , \47798 );
not \U$47457 ( \47800 , \47120 );
not \U$47458 ( \47801 , \47156 );
or \U$47459 ( \47802 , \47800 , \47801 );
or \U$47460 ( \47803 , \47156 , \47120 );
nand \U$47461 ( \47804 , \47802 , \47803 );
xor \U$47462 ( \47805 , \47126 , \47804 );
xor \U$47463 ( \47806 , \47799 , \47805 );
not \U$47464 ( \47807 , \46862 );
xor \U$47465 ( \47808 , \46870 , \46865 );
not \U$47466 ( \47809 , \47808 );
or \U$47467 ( \47810 , \47807 , \47809 );
or \U$47468 ( \47811 , \47808 , \46862 );
nand \U$47469 ( \47812 , \47810 , \47811 );
and \U$47470 ( \47813 , \47806 , \47812 );
and \U$47471 ( \47814 , \47799 , \47805 );
or \U$47472 ( \47815 , \47813 , \47814 );
and \U$47473 ( \47816 , \47795 , \47815 );
and \U$47474 ( \47817 , \47432 , \47794 );
or \U$47475 ( \47818 , \47816 , \47817 );
xor \U$47476 ( \47819 , \46526 , \46771 );
xor \U$47477 ( \47820 , \47819 , \46791 );
xor \U$47478 ( \47821 , \47818 , \47820 );
not \U$47479 ( \47822 , \46843 );
xor \U$47480 ( \47823 , \46857 , \46872 );
not \U$47481 ( \47824 , \47823 );
or \U$47482 ( \47825 , \47822 , \47824 );
or \U$47483 ( \47826 , \47823 , \46843 );
nand \U$47484 ( \47827 , \47825 , \47826 );
xor \U$47485 ( \47828 , \46611 , \46685 );
xor \U$47486 ( \47829 , \47828 , \46768 );
xor \U$47487 ( \47830 , \47827 , \47829 );
xor \U$47488 ( \47831 , \46782 , \46783 );
xor \U$47489 ( \47832 , \47831 , \46788 );
xor \U$47490 ( \47833 , \47251 , \47258 );
xor \U$47491 ( \47834 , \47832 , \47833 );
and \U$47492 ( \47835 , \47830 , \47834 );
and \U$47493 ( \47836 , \47827 , \47829 );
or \U$47494 ( \47837 , \47835 , \47836 );
and \U$47495 ( \47838 , \47821 , \47837 );
and \U$47496 ( \47839 , \47818 , \47820 );
or \U$47497 ( \47840 , \47838 , \47839 );
and \U$47498 ( \47841 , \47376 , \47840 );
not \U$47499 ( \47842 , \47375 );
and \U$47500 ( \47843 , \47362 , \47842 );
nor \U$47501 ( \47844 , \47841 , \47843 );
xnor \U$47502 ( \47845 , \47358 , \47844 );
not \U$47503 ( \47846 , \47845 );
and \U$47504 ( \47847 , \47344 , \47846 );
and \U$47505 ( \47848 , \47845 , \47343 );
nor \U$47506 ( \47849 , \47847 , \47848 );
not \U$47507 ( \47850 , \47362 );
not \U$47508 ( \47851 , \47840 );
not \U$47509 ( \47852 , \47375 );
and \U$47510 ( \47853 , \47851 , \47852 );
and \U$47511 ( \47854 , \47840 , \47375 );
nor \U$47512 ( \47855 , \47853 , \47854 );
not \U$47513 ( \47856 , \47855 );
or \U$47514 ( \47857 , \47850 , \47856 );
or \U$47515 ( \47858 , \47855 , \47362 );
nand \U$47516 ( \47859 , \47857 , \47858 );
not \U$47517 ( \47860 , \47354 );
not \U$47518 ( \47861 , \47357 );
or \U$47519 ( \47862 , \47860 , \47861 );
or \U$47520 ( \47863 , \47357 , \47354 );
nand \U$47521 ( \47864 , \47862 , \47863 );
and \U$47522 ( \47865 , \47859 , \47864 );
not \U$47523 ( \47866 , \47859 );
not \U$47524 ( \47867 , \47864 );
and \U$47525 ( \47868 , \47866 , \47867 );
xor \U$47526 ( \47869 , \47818 , \47820 );
xor \U$47527 ( \47870 , \47869 , \47837 );
not \U$47528 ( \47871 , \47369 );
not \U$47529 ( \47872 , \47374 );
or \U$47530 ( \47873 , \47871 , \47872 );
or \U$47531 ( \47874 , \47374 , \47369 );
nand \U$47532 ( \47875 , \47873 , \47874 );
and \U$47533 ( \47876 , \47870 , \47875 );
not \U$47534 ( \47877 , \47870 );
not \U$47535 ( \47878 , \47875 );
and \U$47536 ( \47879 , \47877 , \47878 );
xor \U$47537 ( \47880 , \46907 , \46915 );
xor \U$47538 ( \47881 , \47880 , \46924 );
xor \U$47539 ( \47882 , \47698 , \47703 );
xor \U$47540 ( \47883 , \47881 , \47882 );
xor \U$47541 ( \47884 , \47756 , \47758 );
xor \U$47542 ( \47885 , \47884 , \47761 );
and \U$47543 ( \47886 , \47883 , \47885 );
xor \U$47544 ( \47887 , \47091 , \47098 );
xor \U$47545 ( \47888 , \47887 , \47106 );
xor \U$47546 ( \47889 , \47770 , \47775 );
xor \U$47547 ( \47890 , \47888 , \47889 );
xor \U$47548 ( \47891 , \47756 , \47758 );
xor \U$47549 ( \47892 , \47891 , \47761 );
and \U$47550 ( \47893 , \47890 , \47892 );
and \U$47551 ( \47894 , \47883 , \47890 );
or \U$47552 ( \47895 , \47886 , \47893 , \47894 );
xor \U$47553 ( \47896 , \47738 , \47739 );
xor \U$47554 ( \47897 , \47896 , \47750 );
xor \U$47555 ( \47898 , \47543 , \47569 );
xor \U$47556 ( \47899 , \47898 , \47598 );
and \U$47557 ( \47900 , \47897 , \47899 );
xor \U$47558 ( \47901 , \47457 , \47484 );
xor \U$47559 ( \47902 , \47901 , \47512 );
xor \U$47560 ( \47903 , \47543 , \47569 );
xor \U$47561 ( \47904 , \47903 , \47598 );
and \U$47562 ( \47905 , \47902 , \47904 );
and \U$47563 ( \47906 , \47897 , \47902 );
or \U$47564 ( \47907 , \47900 , \47905 , \47906 );
xor \U$47565 ( \47908 , \47895 , \47907 );
xor \U$47566 ( \47909 , \47072 , \47083 );
xor \U$47567 ( \47910 , \47909 , \47109 );
xor \U$47568 ( \47911 , \47386 , \47399 );
xor \U$47569 ( \47912 , \47910 , \47911 );
and \U$47570 ( \47913 , \47908 , \47912 );
and \U$47571 ( \47914 , \47895 , \47907 );
or \U$47572 ( \47915 , \47913 , \47914 );
and \U$47573 ( \47916 , \1311 , RI9870b28_100);
and \U$47574 ( \47917 , RI9870df8_106, \1309 );
nor \U$47575 ( \47918 , \47916 , \47917 );
and \U$47576 ( \47919 , \47918 , \1315 );
not \U$47577 ( \47920 , \47918 );
and \U$47578 ( \47921 , \47920 , \1458 );
nor \U$47579 ( \47922 , \47919 , \47921 );
not \U$47580 ( \47923 , \47922 );
and \U$47581 ( \47924 , \2042 , RI9870a38_98);
and \U$47582 ( \47925 , RI9870ee8_108, \2040 );
nor \U$47583 ( \47926 , \47924 , \47925 );
not \U$47584 ( \47927 , \47926 );
not \U$47585 ( \47928 , \2034 );
and \U$47586 ( \47929 , \47927 , \47928 );
and \U$47587 ( \47930 , \47926 , \1462 );
nor \U$47588 ( \47931 , \47929 , \47930 );
not \U$47589 ( \47932 , \47931 );
and \U$47590 ( \47933 , \47923 , \47932 );
and \U$47591 ( \47934 , \47931 , \47922 );
and \U$47592 ( \47935 , \2274 , RI9870c18_102);
and \U$47593 ( \47936 , RI98710c8_112, \2272 );
nor \U$47594 ( \47937 , \47935 , \47936 );
and \U$47595 ( \47938 , \47937 , \2031 );
not \U$47596 ( \47939 , \47937 );
and \U$47597 ( \47940 , \47939 , \2030 );
nor \U$47598 ( \47941 , \47938 , \47940 );
nor \U$47599 ( \47942 , \47934 , \47941 );
nor \U$47600 ( \47943 , \47933 , \47942 );
not \U$47601 ( \47944 , \2935 );
and \U$47602 ( \47945 , \3254 , RI98711b8_114);
and \U$47603 ( \47946 , RI9871398_118, \3252 );
nor \U$47604 ( \47947 , \47945 , \47946 );
not \U$47605 ( \47948 , \47947 );
or \U$47606 ( \47949 , \47944 , \47948 );
or \U$47607 ( \47950 , \47947 , \3406 );
nand \U$47608 ( \47951 , \47949 , \47950 );
not \U$47609 ( \47952 , \3412 );
and \U$47610 ( \47953 , \3683 , RI9871488_120);
and \U$47611 ( \47954 , RI9871758_126, \3681 );
nor \U$47612 ( \47955 , \47953 , \47954 );
not \U$47613 ( \47956 , \47955 );
or \U$47614 ( \47957 , \47952 , \47956 );
or \U$47615 ( \47958 , \47955 , \3412 );
nand \U$47616 ( \47959 , \47957 , \47958 );
xor \U$47617 ( \47960 , \47951 , \47959 );
and \U$47618 ( \47961 , \2464 , RI9870d08_104);
and \U$47619 ( \47962 , RI98712a8_116, \2462 );
nor \U$47620 ( \47963 , \47961 , \47962 );
and \U$47621 ( \47964 , \47963 , \2468 );
not \U$47622 ( \47965 , \47963 );
and \U$47623 ( \47966 , \47965 , \2263 );
nor \U$47624 ( \47967 , \47964 , \47966 );
and \U$47625 ( \47968 , \47960 , \47967 );
and \U$47626 ( \47969 , \47951 , \47959 );
nor \U$47627 ( \47970 , \47968 , \47969 );
xor \U$47628 ( \47971 , \47943 , \47970 );
not \U$47629 ( \47972 , \1128 );
and \U$47630 ( \47973 , \1293 , RI986fef8_74);
and \U$47631 ( \47974 , RI98700d8_78, \1291 );
nor \U$47632 ( \47975 , \47973 , \47974 );
not \U$47633 ( \47976 , \47975 );
or \U$47634 ( \47977 , \47972 , \47976 );
or \U$47635 ( \47978 , \47975 , \1301 );
nand \U$47636 ( \47979 , \47977 , \47978 );
and \U$47637 ( \47980 , \1329 , RI98701c8_80);
and \U$47638 ( \47981 , RI9870fd8_110, \1327 );
nor \U$47639 ( \47982 , \47980 , \47981 );
and \U$47640 ( \47983 , \47982 , \1336 );
not \U$47641 ( \47984 , \47982 );
and \U$47642 ( \47985 , \47984 , \1337 );
nor \U$47643 ( \47986 , \47983 , \47985 );
xor \U$47644 ( \47987 , \47979 , \47986 );
and \U$47645 ( \47988 , \776 , RI986fd18_70);
and \U$47646 ( \47989 , RI986ffe8_76, \774 );
nor \U$47647 ( \47990 , \47988 , \47989 );
and \U$47648 ( \47991 , \47990 , \474 );
not \U$47649 ( \47992 , \47990 );
and \U$47650 ( \47993 , \47992 , \451 );
nor \U$47651 ( \47994 , \47991 , \47993 );
and \U$47652 ( \47995 , \47987 , \47994 );
and \U$47653 ( \47996 , \47979 , \47986 );
nor \U$47654 ( \47997 , \47995 , \47996 );
and \U$47655 ( \47998 , \47971 , \47997 );
and \U$47656 ( \47999 , \47943 , \47970 );
nor \U$47657 ( \48000 , \47998 , \47999 );
and \U$47658 ( \48001 , \15780 , RI986e0f8_10);
and \U$47659 ( \48002 , RI986e2d8_14, RI9873648_192);
nor \U$47660 ( \48003 , \48001 , \48002 );
not \U$47661 ( \48004 , \48003 );
not \U$47662 ( \48005 , RI9873558_190);
and \U$47663 ( \48006 , \48004 , \48005 );
and \U$47664 ( \48007 , \48003 , RI9873558_190);
nor \U$47665 ( \48008 , \48006 , \48007 );
not \U$47666 ( \48009 , \48008 );
not \U$47667 ( \48010 , \422 );
and \U$47668 ( \48011 , \48009 , \48010 );
and \U$47669 ( \48012 , \48008 , \422 );
and \U$47670 ( \48013 , \14937 , RI986dd38_2);
and \U$47671 ( \48014 , RI986e1e8_12, \14935 );
nor \U$47672 ( \48015 , \48013 , \48014 );
and \U$47673 ( \48016 , \48015 , \14538 );
not \U$47674 ( \48017 , \48015 );
and \U$47675 ( \48018 , \48017 , \14539 );
nor \U$47676 ( \48019 , \48016 , \48018 );
nor \U$47677 ( \48020 , \48012 , \48019 );
nor \U$47678 ( \48021 , \48011 , \48020 );
and \U$47679 ( \48022 , \9505 , RI986e698_22);
and \U$47680 ( \48023 , RI986f868_60, \9503 );
nor \U$47681 ( \48024 , \48022 , \48023 );
and \U$47682 ( \48025 , \48024 , \9513 );
not \U$47683 ( \48026 , \48024 );
and \U$47684 ( \48027 , \48026 , \9510 );
nor \U$47685 ( \48028 , \48025 , \48027 );
not \U$47686 ( \48029 , \48028 );
and \U$47687 ( \48030 , \11696 , RI986f958_62);
and \U$47688 ( \48031 , RI986f4a8_52, \11694 );
nor \U$47689 ( \48032 , \48030 , \48031 );
and \U$47690 ( \48033 , \48032 , \11702 );
not \U$47691 ( \48034 , \48032 );
and \U$47692 ( \48035 , \48034 , \10965 );
nor \U$47693 ( \48036 , \48033 , \48035 );
not \U$47694 ( \48037 , \48036 );
and \U$47695 ( \48038 , \48029 , \48037 );
and \U$47696 ( \48039 , \48036 , \48028 );
and \U$47697 ( \48040 , \10424 , RI986f778_58);
and \U$47698 ( \48041 , RI986fa48_64, \10422 );
nor \U$47699 ( \48042 , \48040 , \48041 );
and \U$47700 ( \48043 , \48042 , \10428 );
not \U$47701 ( \48044 , \48042 );
and \U$47702 ( \48045 , \48044 , \9840 );
nor \U$47703 ( \48046 , \48043 , \48045 );
nor \U$47704 ( \48047 , \48039 , \48046 );
nor \U$47705 ( \48048 , \48038 , \48047 );
xor \U$47706 ( \48049 , \48021 , \48048 );
and \U$47707 ( \48050 , \12293 , RI986f3b8_50);
and \U$47708 ( \48051 , RI986f598_54, \12291 );
nor \U$47709 ( \48052 , \48050 , \48051 );
and \U$47710 ( \48053 , \48052 , \11686 );
not \U$47711 ( \48054 , \48052 );
and \U$47712 ( \48055 , \48054 , \11687 );
nor \U$47713 ( \48056 , \48053 , \48055 );
not \U$47714 ( \48057 , \48056 );
and \U$47715 ( \48058 , \13045 , RI986f688_56);
and \U$47716 ( \48059 , RI986e008_8, \13043 );
nor \U$47717 ( \48060 , \48058 , \48059 );
and \U$47718 ( \48061 , \48060 , \12619 );
not \U$47719 ( \48062 , \48060 );
and \U$47720 ( \48063 , \48062 , \13047 );
nor \U$47721 ( \48064 , \48061 , \48063 );
not \U$47722 ( \48065 , \48064 );
and \U$47723 ( \48066 , \48057 , \48065 );
and \U$47724 ( \48067 , \48064 , \48056 );
and \U$47725 ( \48068 , \13882 , RI986df18_6);
and \U$47726 ( \48069 , RI986de28_4, \13880 );
nor \U$47727 ( \48070 , \48068 , \48069 );
and \U$47728 ( \48071 , \48070 , \13359 );
not \U$47729 ( \48072 , \48070 );
and \U$47730 ( \48073 , \48072 , \13358 );
nor \U$47731 ( \48074 , \48071 , \48073 );
nor \U$47732 ( \48075 , \48067 , \48074 );
nor \U$47733 ( \48076 , \48066 , \48075 );
and \U$47734 ( \48077 , \48049 , \48076 );
and \U$47735 ( \48078 , \48021 , \48048 );
nor \U$47736 ( \48079 , \48077 , \48078 );
xor \U$47737 ( \48080 , \48000 , \48079 );
and \U$47738 ( \48081 , \5881 , RI986e878_26);
and \U$47739 ( \48082 , RI986ef08_40, \5879 );
nor \U$47740 ( \48083 , \48081 , \48082 );
and \U$47741 ( \48084 , \48083 , \5885 );
not \U$47742 ( \48085 , \48083 );
and \U$47743 ( \48086 , \48085 , \5594 );
nor \U$47744 ( \48087 , \48084 , \48086 );
not \U$47745 ( \48088 , \48087 );
and \U$47746 ( \48089 , \6453 , RI986ee18_38);
and \U$47747 ( \48090 , RI986ec38_34, \6451 );
nor \U$47748 ( \48091 , \48089 , \48090 );
and \U$47749 ( \48092 , \48091 , \6180 );
not \U$47750 ( \48093 , \48091 );
and \U$47751 ( \48094 , \48093 , \6190 );
nor \U$47752 ( \48095 , \48092 , \48094 );
not \U$47753 ( \48096 , \48095 );
and \U$47754 ( \48097 , \48088 , \48096 );
and \U$47755 ( \48098 , \48095 , \48087 );
and \U$47756 ( \48099 , \7079 , RI986ed28_36);
and \U$47757 ( \48100 , RI986f0e8_44, \7077 );
nor \U$47758 ( \48101 , \48099 , \48100 );
and \U$47759 ( \48102 , \48101 , \6709 );
not \U$47760 ( \48103 , \48101 );
and \U$47761 ( \48104 , \48103 , \6710 );
nor \U$47762 ( \48105 , \48102 , \48104 );
nor \U$47763 ( \48106 , \48098 , \48105 );
nor \U$47764 ( \48107 , \48097 , \48106 );
and \U$47765 ( \48108 , \8486 , RI986f1d8_46);
and \U$47766 ( \48109 , RI986e5a8_20, \8484 );
nor \U$47767 ( \48110 , \48108 , \48109 );
and \U$47768 ( \48111 , \48110 , \8050 );
not \U$47769 ( \48112 , \48110 );
and \U$47770 ( \48113 , \48112 , \8051 );
nor \U$47771 ( \48114 , \48111 , \48113 );
and \U$47772 ( \48115 , \9237 , RI986e4b8_18);
and \U$47773 ( \48116 , RI986e788_24, \9235 );
nor \U$47774 ( \48117 , \48115 , \48116 );
and \U$47775 ( \48118 , \48117 , \9241 );
not \U$47776 ( \48119 , \48117 );
and \U$47777 ( \48120 , \48119 , \8836 );
nor \U$47778 ( \48121 , \48118 , \48120 );
xor \U$47779 ( \48122 , \48114 , \48121 );
and \U$47780 ( \48123 , \7729 , RI986eff8_42);
and \U$47781 ( \48124 , RI986f2c8_48, \7727 );
nor \U$47782 ( \48125 , \48123 , \48124 );
and \U$47783 ( \48126 , \48125 , \7480 );
not \U$47784 ( \48127 , \48125 );
and \U$47785 ( \48128 , \48127 , \7733 );
nor \U$47786 ( \48129 , \48126 , \48128 );
and \U$47787 ( \48130 , \48122 , \48129 );
and \U$47788 ( \48131 , \48114 , \48121 );
nor \U$47789 ( \48132 , \48130 , \48131 );
xor \U$47790 ( \48133 , \48107 , \48132 );
not \U$47791 ( \48134 , \4519 );
and \U$47792 ( \48135 , \4710 , RI9871668_124);
and \U$47793 ( \48136 , RI986eb48_32, \4708 );
nor \U$47794 ( \48137 , \48135 , \48136 );
not \U$47795 ( \48138 , \48137 );
or \U$47796 ( \48139 , \48134 , \48138 );
or \U$47797 ( \48140 , \48137 , \4521 );
nand \U$47798 ( \48141 , \48139 , \48140 );
and \U$47799 ( \48142 , \5318 , RI986ea58_30);
and \U$47800 ( \48143 , RI986e968_28, \5316 );
nor \U$47801 ( \48144 , \48142 , \48143 );
and \U$47802 ( \48145 , \48144 , \5052 );
not \U$47803 ( \48146 , \48144 );
and \U$47804 ( \48147 , \48146 , \5322 );
nor \U$47805 ( \48148 , \48145 , \48147 );
xor \U$47806 ( \48149 , \48141 , \48148 );
and \U$47807 ( \48150 , \4203 , RI9871848_128);
and \U$47808 ( \48151 , RI9871578_122, \4201 );
nor \U$47809 ( \48152 , \48150 , \48151 );
and \U$47810 ( \48153 , \48152 , \4207 );
not \U$47811 ( \48154 , \48152 );
and \U$47812 ( \48155 , \48154 , \3922 );
nor \U$47813 ( \48156 , \48153 , \48155 );
and \U$47814 ( \48157 , \48149 , \48156 );
and \U$47815 ( \48158 , \48141 , \48148 );
nor \U$47816 ( \48159 , \48157 , \48158 );
and \U$47817 ( \48160 , \48133 , \48159 );
and \U$47818 ( \48161 , \48107 , \48132 );
nor \U$47819 ( \48162 , \48160 , \48161 );
and \U$47820 ( \48163 , \48080 , \48162 );
and \U$47821 ( \48164 , \48000 , \48079 );
nor \U$47822 ( \48165 , \48163 , \48164 );
not \U$47823 ( \48166 , \48165 );
xor \U$47824 ( \48167 , \47636 , \47644 );
xor \U$47825 ( \48168 , \48167 , \47651 );
not \U$47826 ( \48169 , \48168 );
not \U$47827 ( \48170 , \47662 );
xor \U$47828 ( \48171 , \47680 , \47670 );
not \U$47829 ( \48172 , \48171 );
or \U$47830 ( \48173 , \48170 , \48172 );
or \U$47831 ( \48174 , \48171 , \47662 );
nand \U$47832 ( \48175 , \48173 , \48174 );
nand \U$47833 ( \48176 , \48169 , \48175 );
not \U$47834 ( \48177 , \47079 );
not \U$47835 ( \48178 , \47082 );
and \U$47836 ( \48179 , \48177 , \48178 );
and \U$47837 ( \48180 , \47079 , \47082 );
nor \U$47838 ( \48181 , \48179 , \48180 );
xor \U$47839 ( \48182 , \48176 , \48181 );
not \U$47840 ( \48183 , \47464 );
xor \U$47841 ( \48184 , \47472 , \47482 );
not \U$47842 ( \48185 , \48184 );
or \U$47843 ( \48186 , \48183 , \48185 );
or \U$47844 ( \48187 , \48184 , \47464 );
nand \U$47845 ( \48188 , \48186 , \48187 );
xor \U$47846 ( \48189 , \47439 , \47446 );
xor \U$47847 ( \48190 , \48189 , \47454 );
xor \U$47848 ( \48191 , \48188 , \48190 );
not \U$47849 ( \48192 , \47609 );
xor \U$47850 ( \48193 , \47627 , \47617 );
not \U$47851 ( \48194 , \48193 );
or \U$47852 ( \48195 , \48192 , \48194 );
or \U$47853 ( \48196 , \48193 , \47609 );
nand \U$47854 ( \48197 , \48195 , \48196 );
and \U$47855 ( \48198 , \48191 , \48197 );
and \U$47856 ( \48199 , \48188 , \48190 );
nor \U$47857 ( \48200 , \48198 , \48199 );
and \U$47858 ( \48201 , \48182 , \48200 );
and \U$47859 ( \48202 , \48176 , \48181 );
or \U$47860 ( \48203 , \48201 , \48202 );
not \U$47861 ( \48204 , \48203 );
and \U$47862 ( \48205 , \48166 , \48204 );
and \U$47863 ( \48206 , \48165 , \48203 );
not \U$47864 ( \48207 , \47585 );
xor \U$47865 ( \48208 , \47577 , \47596 );
not \U$47866 ( \48209 , \48208 );
or \U$47867 ( \48210 , \48207 , \48209 );
or \U$47868 ( \48211 , \48208 , \47585 );
nand \U$47869 ( \48212 , \48210 , \48211 );
and \U$47870 ( \48213 , \416 , RI9870498_86);
and \U$47871 ( \48214 , RI9870588_88, \414 );
nor \U$47872 ( \48215 , \48213 , \48214 );
and \U$47873 ( \48216 , \48215 , \422 );
not \U$47874 ( \48217 , \48215 );
and \U$47875 ( \48218 , \48217 , \421 );
nor \U$47876 ( \48219 , \48216 , \48218 );
xor \U$47877 ( \48220 , \48212 , \48219 );
not \U$47878 ( \48221 , \47725 );
xor \U$47879 ( \48222 , \47736 , \47716 );
not \U$47880 ( \48223 , \48222 );
or \U$47881 ( \48224 , \48221 , \48223 );
or \U$47882 ( \48225 , \48222 , \47725 );
nand \U$47883 ( \48226 , \48224 , \48225 );
and \U$47884 ( \48227 , \48220 , \48226 );
and \U$47885 ( \48228 , \48212 , \48219 );
or \U$47886 ( \48229 , \48227 , \48228 );
not \U$47887 ( \48230 , \361 );
and \U$47888 ( \48231 , \354 , RI9870588_88);
and \U$47889 ( \48232 , RI98703a8_84, \352 );
nor \U$47890 ( \48233 , \48231 , \48232 );
not \U$47891 ( \48234 , \48233 );
or \U$47892 ( \48235 , \48230 , \48234 );
or \U$47893 ( \48236 , \48233 , \345 );
nand \U$47894 ( \48237 , \48235 , \48236 );
nand \U$47895 ( \48238 , RI9870498_86, \414 );
and \U$47896 ( \48239 , \48238 , \422 );
not \U$47897 ( \48240 , \48238 );
and \U$47898 ( \48241 , \48240 , \421 );
nor \U$47899 ( \48242 , \48239 , \48241 );
xor \U$47900 ( \48243 , \48237 , \48242 );
not \U$47901 ( \48244 , \487 );
and \U$47902 ( \48245 , \395 , RI98702b8_82);
and \U$47903 ( \48246 , RI9870768_92, \393 );
nor \U$47904 ( \48247 , \48245 , \48246 );
not \U$47905 ( \48248 , \48247 );
or \U$47906 ( \48249 , \48244 , \48248 );
or \U$47907 ( \48250 , \48247 , \487 );
nand \U$47908 ( \48251 , \48249 , \48250 );
and \U$47909 ( \48252 , \48243 , \48251 );
and \U$47910 ( \48253 , \48237 , \48242 );
or \U$47911 ( \48254 , \48252 , \48253 );
not \U$47912 ( \48255 , \345 );
and \U$47913 ( \48256 , \354 , RI98703a8_84);
and \U$47914 ( \48257 , RI98702b8_82, \352 );
nor \U$47915 ( \48258 , \48256 , \48257 );
not \U$47916 ( \48259 , \48258 );
or \U$47917 ( \48260 , \48255 , \48259 );
or \U$47918 ( \48261 , \48258 , \345 );
nand \U$47919 ( \48262 , \48260 , \48261 );
xor \U$47920 ( \48263 , \48254 , \48262 );
not \U$47921 ( \48264 , \367 );
and \U$47922 ( \48265 , \376 , RI9870678_90);
and \U$47923 ( \48266 , RI9870948_96, \374 );
nor \U$47924 ( \48267 , \48265 , \48266 );
not \U$47925 ( \48268 , \48267 );
or \U$47926 ( \48269 , \48264 , \48268 );
or \U$47927 ( \48270 , \48267 , \365 );
nand \U$47928 ( \48271 , \48269 , \48270 );
and \U$47929 ( \48272 , \438 , RI986fc28_68);
and \U$47930 ( \48273 , RI986fe08_72, \436 );
nor \U$47931 ( \48274 , \48272 , \48273 );
and \U$47932 ( \48275 , \48274 , \444 );
not \U$47933 ( \48276 , \48274 );
and \U$47934 ( \48277 , \48276 , \443 );
nor \U$47935 ( \48278 , \48275 , \48277 );
xor \U$47936 ( \48279 , \48271 , \48278 );
not \U$47937 ( \48280 , \456 );
and \U$47938 ( \48281 , \465 , RI9870858_94);
and \U$47939 ( \48282 , RI986fb38_66, \463 );
nor \U$47940 ( \48283 , \48281 , \48282 );
not \U$47941 ( \48284 , \48283 );
or \U$47942 ( \48285 , \48280 , \48284 );
or \U$47943 ( \48286 , \48283 , \454 );
nand \U$47944 ( \48287 , \48285 , \48286 );
and \U$47945 ( \48288 , \48279 , \48287 );
and \U$47946 ( \48289 , \48271 , \48278 );
or \U$47947 ( \48290 , \48288 , \48289 );
and \U$47948 ( \48291 , \48263 , \48290 );
and \U$47949 ( \48292 , \48254 , \48262 );
or \U$47950 ( \48293 , \48291 , \48292 );
xor \U$47951 ( \48294 , \48229 , \48293 );
not \U$47952 ( \48295 , \47522 );
xor \U$47953 ( \48296 , \47530 , \47541 );
not \U$47954 ( \48297 , \48296 );
or \U$47955 ( \48298 , \48295 , \48297 );
or \U$47956 ( \48299 , \48296 , \47522 );
nand \U$47957 ( \48300 , \48298 , \48299 );
xor \U$47958 ( \48301 , \47550 , \47558 );
xor \U$47959 ( \48302 , \48301 , \47566 );
xor \U$47960 ( \48303 , \48300 , \48302 );
xor \U$47961 ( \48304 , \47492 , \47500 );
xor \U$47962 ( \48305 , \48304 , \47509 );
and \U$47963 ( \48306 , \48303 , \48305 );
and \U$47964 ( \48307 , \48300 , \48302 );
or \U$47965 ( \48308 , \48306 , \48307 );
and \U$47966 ( \48309 , \48294 , \48308 );
and \U$47967 ( \48310 , \48229 , \48293 );
nor \U$47968 ( \48311 , \48309 , \48310 );
nor \U$47969 ( \48312 , \48206 , \48311 );
nor \U$47970 ( \48313 , \48205 , \48312 );
xor \U$47971 ( \48314 , \47915 , \48313 );
not \U$47972 ( \48315 , \47420 );
not \U$47973 ( \48316 , \47428 );
or \U$47974 ( \48317 , \48315 , \48316 );
or \U$47975 ( \48318 , \47428 , \47420 );
nand \U$47976 ( \48319 , \48317 , \48318 );
not \U$47977 ( \48320 , \48319 );
not \U$47978 ( \48321 , \47422 );
and \U$47979 ( \48322 , \48320 , \48321 );
and \U$47980 ( \48323 , \48319 , \47422 );
nor \U$47981 ( \48324 , \48322 , \48323 );
xor \U$47982 ( \48325 , \47708 , \47753 );
xor \U$47983 ( \48326 , \48325 , \47764 );
xor \U$47984 ( \48327 , \48324 , \48326 );
xor \U$47985 ( \48328 , \47780 , \47785 );
xor \U$47986 ( \48329 , \48328 , \47788 );
and \U$47987 ( \48330 , \48327 , \48329 );
and \U$47988 ( \48331 , \48324 , \48326 );
or \U$47989 ( \48332 , \48330 , \48331 );
and \U$47990 ( \48333 , \48314 , \48332 );
and \U$47991 ( \48334 , \47915 , \48313 );
or \U$47992 ( \48335 , \48333 , \48334 );
not \U$47993 ( \48336 , \48335 );
xor \U$47994 ( \48337 , \47114 , \47158 );
xor \U$47995 ( \48338 , \48337 , \47242 );
not \U$47996 ( \48339 , \48338 );
and \U$47997 ( \48340 , \48336 , \48339 );
and \U$47998 ( \48341 , \48335 , \48338 );
not \U$47999 ( \48342 , \47112 );
xor \U$48000 ( \48343 , \47043 , \46959 );
not \U$48001 ( \48344 , \48343 );
or \U$48002 ( \48345 , \48342 , \48344 );
or \U$48003 ( \48346 , \48343 , \47112 );
nand \U$48004 ( \48347 , \48345 , \48346 );
not \U$48005 ( \48348 , \47227 );
xor \U$48006 ( \48349 , \47169 , \47240 );
not \U$48007 ( \48350 , \48349 );
or \U$48008 ( \48351 , \48348 , \48350 );
or \U$48009 ( \48352 , \48349 , \47227 );
nand \U$48010 ( \48353 , \48351 , \48352 );
xor \U$48011 ( \48354 , \48347 , \48353 );
xor \U$48012 ( \48355 , \47799 , \47805 );
xor \U$48013 ( \48356 , \48355 , \47812 );
and \U$48014 ( \48357 , \48354 , \48356 );
and \U$48015 ( \48358 , \48347 , \48353 );
nor \U$48016 ( \48359 , \48357 , \48358 );
nor \U$48017 ( \48360 , \48341 , \48359 );
nor \U$48018 ( \48361 , \48340 , \48360 );
nor \U$48019 ( \48362 , \47879 , \48361 );
nor \U$48020 ( \48363 , \47876 , \48362 );
nor \U$48021 ( \48364 , \47868 , \48363 );
nor \U$48022 ( \48365 , \47865 , \48364 );
xor \U$48023 ( \48366 , \47849 , \48365 );
xor \U$48024 ( \48367 , \48141 , \48148 );
xor \U$48025 ( \48368 , \48367 , \48156 );
not \U$48026 ( \48369 , \48087 );
xor \U$48027 ( \48370 , \48095 , \48105 );
not \U$48028 ( \48371 , \48370 );
or \U$48029 ( \48372 , \48369 , \48371 );
or \U$48030 ( \48373 , \48370 , \48087 );
nand \U$48031 ( \48374 , \48372 , \48373 );
xor \U$48032 ( \48375 , \48368 , \48374 );
xor \U$48033 ( \48376 , \48114 , \48121 );
xor \U$48034 ( \48377 , \48376 , \48129 );
and \U$48035 ( \48378 , \48375 , \48377 );
and \U$48036 ( \48379 , \48368 , \48374 );
or \U$48037 ( \48380 , \48378 , \48379 );
not \U$48038 ( \48381 , \367 );
and \U$48039 ( \48382 , \376 , RI9870768_92);
and \U$48040 ( \48383 , RI9870678_90, \374 );
nor \U$48041 ( \48384 , \48382 , \48383 );
not \U$48042 ( \48385 , \48384 );
or \U$48043 ( \48386 , \48381 , \48385 );
or \U$48044 ( \48387 , \48384 , \365 );
nand \U$48045 ( \48388 , \48386 , \48387 );
not \U$48046 ( \48389 , \454 );
and \U$48047 ( \48390 , \465 , RI9870948_96);
and \U$48048 ( \48391 , RI9870858_94, \463 );
nor \U$48049 ( \48392 , \48390 , \48391 );
not \U$48050 ( \48393 , \48392 );
or \U$48051 ( \48394 , \48389 , \48393 );
or \U$48052 ( \48395 , \48392 , \454 );
nand \U$48053 ( \48396 , \48394 , \48395 );
xor \U$48054 ( \48397 , \48388 , \48396 );
not \U$48055 ( \48398 , \487 );
and \U$48056 ( \48399 , \395 , RI98703a8_84);
and \U$48057 ( \48400 , RI98702b8_82, \393 );
nor \U$48058 ( \48401 , \48399 , \48400 );
not \U$48059 ( \48402 , \48401 );
or \U$48060 ( \48403 , \48398 , \48402 );
or \U$48061 ( \48404 , \48401 , \487 );
nand \U$48062 ( \48405 , \48403 , \48404 );
and \U$48063 ( \48406 , \48397 , \48405 );
and \U$48064 ( \48407 , \48388 , \48396 );
or \U$48065 ( \48408 , \48406 , \48407 );
xor \U$48066 ( \48409 , \48237 , \48242 );
xor \U$48067 ( \48410 , \48409 , \48251 );
and \U$48068 ( \48411 , \48408 , \48410 );
xor \U$48069 ( \48412 , \48271 , \48278 );
xor \U$48070 ( \48413 , \48412 , \48287 );
xor \U$48071 ( \48414 , \48237 , \48242 );
xor \U$48072 ( \48415 , \48414 , \48251 );
and \U$48073 ( \48416 , \48413 , \48415 );
and \U$48074 ( \48417 , \48408 , \48413 );
or \U$48075 ( \48418 , \48411 , \48416 , \48417 );
xor \U$48076 ( \48419 , \48380 , \48418 );
not \U$48077 ( \48420 , \47922 );
xor \U$48078 ( \48421 , \47931 , \47941 );
not \U$48079 ( \48422 , \48421 );
or \U$48080 ( \48423 , \48420 , \48422 );
or \U$48081 ( \48424 , \48421 , \47922 );
nand \U$48082 ( \48425 , \48423 , \48424 );
xor \U$48083 ( \48426 , \47979 , \47986 );
xor \U$48084 ( \48427 , \48426 , \47994 );
xor \U$48085 ( \48428 , \48425 , \48427 );
xor \U$48086 ( \48429 , \47951 , \47959 );
xor \U$48087 ( \48430 , \48429 , \47967 );
and \U$48088 ( \48431 , \48428 , \48430 );
and \U$48089 ( \48432 , \48425 , \48427 );
or \U$48090 ( \48433 , \48431 , \48432 );
and \U$48091 ( \48434 , \48419 , \48433 );
and \U$48092 ( \48435 , \48380 , \48418 );
or \U$48093 ( \48436 , \48434 , \48435 );
and \U$48094 ( \48437 , \8486 , RI986f2c8_48);
and \U$48095 ( \48438 , RI986f1d8_46, \8484 );
nor \U$48096 ( \48439 , \48437 , \48438 );
and \U$48097 ( \48440 , \48439 , \8050 );
not \U$48098 ( \48441 , \48439 );
and \U$48099 ( \48442 , \48441 , \8051 );
nor \U$48100 ( \48443 , \48440 , \48442 );
and \U$48101 ( \48444 , \7079 , RI986ec38_34);
and \U$48102 ( \48445 , RI986ed28_36, \7077 );
nor \U$48103 ( \48446 , \48444 , \48445 );
and \U$48104 ( \48447 , \48446 , \6710 );
not \U$48105 ( \48448 , \48446 );
and \U$48106 ( \48449 , \48448 , \6709 );
nor \U$48107 ( \48450 , \48447 , \48449 );
xor \U$48108 ( \48451 , \48443 , \48450 );
and \U$48109 ( \48452 , \7729 , RI986f0e8_44);
and \U$48110 ( \48453 , RI986eff8_42, \7727 );
nor \U$48111 ( \48454 , \48452 , \48453 );
and \U$48112 ( \48455 , \48454 , \7480 );
not \U$48113 ( \48456 , \48454 );
and \U$48114 ( \48457 , \48456 , \7733 );
nor \U$48115 ( \48458 , \48455 , \48457 );
and \U$48116 ( \48459 , \48451 , \48458 );
and \U$48117 ( \48460 , \48443 , \48450 );
or \U$48118 ( \48461 , \48459 , \48460 );
not \U$48119 ( \48462 , \3918 );
and \U$48120 ( \48463 , \3683 , RI9871398_118);
and \U$48121 ( \48464 , RI9871488_120, \3681 );
nor \U$48122 ( \48465 , \48463 , \48464 );
not \U$48123 ( \48466 , \48465 );
or \U$48124 ( \48467 , \48462 , \48466 );
or \U$48125 ( \48468 , \48465 , \3412 );
nand \U$48126 ( \48469 , \48467 , \48468 );
and \U$48127 ( \48470 , \4203 , RI9871758_126);
and \U$48128 ( \48471 , RI9871848_128, \4201 );
nor \U$48129 ( \48472 , \48470 , \48471 );
and \U$48130 ( \48473 , \48472 , \4207 );
not \U$48131 ( \48474 , \48472 );
and \U$48132 ( \48475 , \48474 , \3922 );
nor \U$48133 ( \48476 , \48473 , \48475 );
xor \U$48134 ( \48477 , \48469 , \48476 );
not \U$48135 ( \48478 , \4519 );
and \U$48136 ( \48479 , \4710 , RI9871578_122);
and \U$48137 ( \48480 , RI9871668_124, \4708 );
nor \U$48138 ( \48481 , \48479 , \48480 );
not \U$48139 ( \48482 , \48481 );
or \U$48140 ( \48483 , \48478 , \48482 );
or \U$48141 ( \48484 , \48481 , \4521 );
nand \U$48142 ( \48485 , \48483 , \48484 );
and \U$48143 ( \48486 , \48477 , \48485 );
and \U$48144 ( \48487 , \48469 , \48476 );
or \U$48145 ( \48488 , \48486 , \48487 );
xor \U$48146 ( \48489 , \48461 , \48488 );
and \U$48147 ( \48490 , \5318 , RI986eb48_32);
and \U$48148 ( \48491 , RI986ea58_30, \5316 );
nor \U$48149 ( \48492 , \48490 , \48491 );
and \U$48150 ( \48493 , \48492 , \5052 );
not \U$48151 ( \48494 , \48492 );
and \U$48152 ( \48495 , \48494 , \5322 );
nor \U$48153 ( \48496 , \48493 , \48495 );
and \U$48154 ( \48497 , \5881 , RI986e968_28);
and \U$48155 ( \48498 , RI986e878_26, \5879 );
nor \U$48156 ( \48499 , \48497 , \48498 );
and \U$48157 ( \48500 , \48499 , \5594 );
not \U$48158 ( \48501 , \48499 );
and \U$48159 ( \48502 , \48501 , \5885 );
nor \U$48160 ( \48503 , \48500 , \48502 );
xor \U$48161 ( \48504 , \48496 , \48503 );
and \U$48162 ( \48505 , \6453 , RI986ef08_40);
and \U$48163 ( \48506 , RI986ee18_38, \6451 );
nor \U$48164 ( \48507 , \48505 , \48506 );
and \U$48165 ( \48508 , \48507 , \6190 );
not \U$48166 ( \48509 , \48507 );
and \U$48167 ( \48510 , \48509 , \6180 );
nor \U$48168 ( \48511 , \48508 , \48510 );
and \U$48169 ( \48512 , \48504 , \48511 );
and \U$48170 ( \48513 , \48496 , \48503 );
or \U$48171 ( \48514 , \48512 , \48513 );
and \U$48172 ( \48515 , \48489 , \48514 );
and \U$48173 ( \48516 , \48461 , \48488 );
or \U$48174 ( \48517 , \48515 , \48516 );
and \U$48175 ( \48518 , \11696 , RI986fa48_64);
and \U$48176 ( \48519 , RI986f958_62, \11694 );
nor \U$48177 ( \48520 , \48518 , \48519 );
and \U$48178 ( \48521 , \48520 , \10965 );
not \U$48179 ( \48522 , \48520 );
and \U$48180 ( \48523 , \48522 , \11702 );
nor \U$48181 ( \48524 , \48521 , \48523 );
and \U$48182 ( \48525 , \12293 , RI986f4a8_52);
and \U$48183 ( \48526 , RI986f3b8_50, \12291 );
nor \U$48184 ( \48527 , \48525 , \48526 );
and \U$48185 ( \48528 , \48527 , \11687 );
not \U$48186 ( \48529 , \48527 );
and \U$48187 ( \48530 , \48529 , \11686 );
nor \U$48188 ( \48531 , \48528 , \48530 );
xor \U$48189 ( \48532 , \48524 , \48531 );
and \U$48190 ( \48533 , \13045 , RI986f598_54);
and \U$48191 ( \48534 , RI986f688_56, \13043 );
nor \U$48192 ( \48535 , \48533 , \48534 );
and \U$48193 ( \48536 , \48535 , \13047 );
not \U$48194 ( \48537 , \48535 );
and \U$48195 ( \48538 , \48537 , \12619 );
nor \U$48196 ( \48539 , \48536 , \48538 );
and \U$48197 ( \48540 , \48532 , \48539 );
and \U$48198 ( \48541 , \48524 , \48531 );
or \U$48199 ( \48542 , \48540 , \48541 );
and \U$48200 ( \48543 , \13882 , RI986e008_8);
and \U$48201 ( \48544 , RI986df18_6, \13880 );
nor \U$48202 ( \48545 , \48543 , \48544 );
and \U$48203 ( \48546 , \48545 , \13358 );
not \U$48204 ( \48547 , \48545 );
and \U$48205 ( \48548 , \48547 , \13359 );
nor \U$48206 ( \48549 , \48546 , \48548 );
not \U$48207 ( \48550 , RI9873558_190);
and \U$48208 ( \48551 , \15780 , RI986e1e8_12);
and \U$48209 ( \48552 , RI986e0f8_10, RI9873648_192);
nor \U$48210 ( \48553 , \48551 , \48552 );
not \U$48211 ( \48554 , \48553 );
or \U$48212 ( \48555 , \48550 , \48554 );
or \U$48213 ( \48556 , \48553 , RI9873558_190);
nand \U$48214 ( \48557 , \48555 , \48556 );
xor \U$48215 ( \48558 , \48549 , \48557 );
and \U$48216 ( \48559 , \14937 , RI986de28_4);
and \U$48217 ( \48560 , RI986dd38_2, \14935 );
nor \U$48218 ( \48561 , \48559 , \48560 );
and \U$48219 ( \48562 , \48561 , \14539 );
not \U$48220 ( \48563 , \48561 );
and \U$48221 ( \48564 , \48563 , \14538 );
nor \U$48222 ( \48565 , \48562 , \48564 );
and \U$48223 ( \48566 , \48558 , \48565 );
and \U$48224 ( \48567 , \48549 , \48557 );
or \U$48225 ( \48568 , \48566 , \48567 );
xor \U$48226 ( \48569 , \48542 , \48568 );
and \U$48227 ( \48570 , \9237 , RI986e5a8_20);
and \U$48228 ( \48571 , RI986e4b8_18, \9235 );
nor \U$48229 ( \48572 , \48570 , \48571 );
and \U$48230 ( \48573 , \48572 , \9241 );
not \U$48231 ( \48574 , \48572 );
and \U$48232 ( \48575 , \48574 , \8836 );
nor \U$48233 ( \48576 , \48573 , \48575 );
and \U$48234 ( \48577 , \9505 , RI986e788_24);
and \U$48235 ( \48578 , RI986e698_22, \9503 );
nor \U$48236 ( \48579 , \48577 , \48578 );
and \U$48237 ( \48580 , \48579 , \9510 );
not \U$48238 ( \48581 , \48579 );
and \U$48239 ( \48582 , \48581 , \9513 );
nor \U$48240 ( \48583 , \48580 , \48582 );
xor \U$48241 ( \48584 , \48576 , \48583 );
and \U$48242 ( \48585 , \10424 , RI986f868_60);
and \U$48243 ( \48586 , RI986f778_58, \10422 );
nor \U$48244 ( \48587 , \48585 , \48586 );
and \U$48245 ( \48588 , \48587 , \9840 );
not \U$48246 ( \48589 , \48587 );
and \U$48247 ( \48590 , \48589 , \10428 );
nor \U$48248 ( \48591 , \48588 , \48590 );
and \U$48249 ( \48592 , \48584 , \48591 );
and \U$48250 ( \48593 , \48576 , \48583 );
or \U$48251 ( \48594 , \48592 , \48593 );
and \U$48252 ( \48595 , \48569 , \48594 );
and \U$48253 ( \48596 , \48542 , \48568 );
or \U$48254 ( \48597 , \48595 , \48596 );
xor \U$48255 ( \48598 , \48517 , \48597 );
and \U$48256 ( \48599 , \2274 , RI9870ee8_108);
and \U$48257 ( \48600 , RI9870c18_102, \2272 );
nor \U$48258 ( \48601 , \48599 , \48600 );
and \U$48259 ( \48602 , \48601 , \2030 );
not \U$48260 ( \48603 , \48601 );
and \U$48261 ( \48604 , \48603 , \2031 );
nor \U$48262 ( \48605 , \48602 , \48604 );
and \U$48263 ( \48606 , \2464 , RI98710c8_112);
and \U$48264 ( \48607 , RI9870d08_104, \2462 );
nor \U$48265 ( \48608 , \48606 , \48607 );
and \U$48266 ( \48609 , \48608 , \2468 );
not \U$48267 ( \48610 , \48608 );
and \U$48268 ( \48611 , \48610 , \2263 );
nor \U$48269 ( \48612 , \48609 , \48611 );
xor \U$48270 ( \48613 , \48605 , \48612 );
not \U$48271 ( \48614 , \3406 );
and \U$48272 ( \48615 , \3254 , RI98712a8_116);
and \U$48273 ( \48616 , RI98711b8_114, \3252 );
nor \U$48274 ( \48617 , \48615 , \48616 );
not \U$48275 ( \48618 , \48617 );
or \U$48276 ( \48619 , \48614 , \48618 );
or \U$48277 ( \48620 , \48617 , \2935 );
nand \U$48278 ( \48621 , \48619 , \48620 );
and \U$48279 ( \48622 , \48613 , \48621 );
and \U$48280 ( \48623 , \48605 , \48612 );
or \U$48281 ( \48624 , \48622 , \48623 );
and \U$48282 ( \48625 , \1329 , RI98700d8_78);
and \U$48283 ( \48626 , RI98701c8_80, \1327 );
nor \U$48284 ( \48627 , \48625 , \48626 );
and \U$48285 ( \48628 , \48627 , \1336 );
not \U$48286 ( \48629 , \48627 );
and \U$48287 ( \48630 , \48629 , \1337 );
nor \U$48288 ( \48631 , \48628 , \48630 );
and \U$48289 ( \48632 , \1311 , RI9870fd8_110);
and \U$48290 ( \48633 , RI9870b28_100, \1309 );
nor \U$48291 ( \48634 , \48632 , \48633 );
and \U$48292 ( \48635 , \48634 , \1458 );
not \U$48293 ( \48636 , \48634 );
and \U$48294 ( \48637 , \48636 , \1318 );
nor \U$48295 ( \48638 , \48635 , \48637 );
xor \U$48296 ( \48639 , \48631 , \48638 );
not \U$48297 ( \48640 , \2034 );
and \U$48298 ( \48641 , \2042 , RI9870df8_106);
and \U$48299 ( \48642 , RI9870a38_98, \2040 );
nor \U$48300 ( \48643 , \48641 , \48642 );
not \U$48301 ( \48644 , \48643 );
or \U$48302 ( \48645 , \48640 , \48644 );
or \U$48303 ( \48646 , \48643 , \2034 );
nand \U$48304 ( \48647 , \48645 , \48646 );
and \U$48305 ( \48648 , \48639 , \48647 );
and \U$48306 ( \48649 , \48631 , \48638 );
or \U$48307 ( \48650 , \48648 , \48649 );
xor \U$48308 ( \48651 , \48624 , \48650 );
and \U$48309 ( \48652 , \776 , RI986fe08_72);
and \U$48310 ( \48653 , RI986fd18_70, \774 );
nor \U$48311 ( \48654 , \48652 , \48653 );
and \U$48312 ( \48655 , \48654 , \474 );
not \U$48313 ( \48656 , \48654 );
and \U$48314 ( \48657 , \48656 , \451 );
nor \U$48315 ( \48658 , \48655 , \48657 );
and \U$48316 ( \48659 , \438 , RI986fb38_66);
and \U$48317 ( \48660 , RI986fc28_68, \436 );
nor \U$48318 ( \48661 , \48659 , \48660 );
and \U$48319 ( \48662 , \48661 , \444 );
not \U$48320 ( \48663 , \48661 );
and \U$48321 ( \48664 , \48663 , \443 );
nor \U$48322 ( \48665 , \48662 , \48664 );
xor \U$48323 ( \48666 , \48658 , \48665 );
not \U$48324 ( \48667 , \1301 );
and \U$48325 ( \48668 , \1293 , RI986ffe8_76);
and \U$48326 ( \48669 , RI986fef8_74, \1291 );
nor \U$48327 ( \48670 , \48668 , \48669 );
not \U$48328 ( \48671 , \48670 );
or \U$48329 ( \48672 , \48667 , \48671 );
or \U$48330 ( \48673 , \48670 , \1128 );
nand \U$48331 ( \48674 , \48672 , \48673 );
and \U$48332 ( \48675 , \48666 , \48674 );
and \U$48333 ( \48676 , \48658 , \48665 );
or \U$48334 ( \48677 , \48675 , \48676 );
and \U$48335 ( \48678 , \48651 , \48677 );
and \U$48336 ( \48679 , \48624 , \48650 );
or \U$48337 ( \48680 , \48678 , \48679 );
and \U$48338 ( \48681 , \48598 , \48680 );
and \U$48339 ( \48682 , \48517 , \48597 );
or \U$48340 ( \48683 , \48681 , \48682 );
xor \U$48341 ( \48684 , \48436 , \48683 );
not \U$48342 ( \48685 , \48028 );
xor \U$48343 ( \48686 , \48046 , \48036 );
not \U$48344 ( \48687 , \48686 );
or \U$48345 ( \48688 , \48685 , \48687 );
or \U$48346 ( \48689 , \48686 , \48028 );
nand \U$48347 ( \48690 , \48688 , \48689 );
not \U$48348 ( \48691 , \48056 );
xor \U$48349 ( \48692 , \48064 , \48074 );
not \U$48350 ( \48693 , \48692 );
or \U$48351 ( \48694 , \48691 , \48693 );
or \U$48352 ( \48695 , \48692 , \48056 );
nand \U$48353 ( \48696 , \48694 , \48695 );
xor \U$48354 ( \48697 , \48690 , \48696 );
not \U$48355 ( \48698 , \421 );
xnor \U$48356 ( \48699 , \48019 , \48008 );
not \U$48357 ( \48700 , \48699 );
or \U$48358 ( \48701 , \48698 , \48700 );
or \U$48359 ( \48702 , \48699 , \421 );
nand \U$48360 ( \48703 , \48701 , \48702 );
and \U$48361 ( \48704 , \48697 , \48703 );
and \U$48362 ( \48705 , \48690 , \48696 );
or \U$48363 ( \48706 , \48704 , \48705 );
not \U$48364 ( \48707 , \48175 );
not \U$48365 ( \48708 , \48168 );
or \U$48366 ( \48709 , \48707 , \48708 );
or \U$48367 ( \48710 , \48168 , \48175 );
nand \U$48368 ( \48711 , \48709 , \48710 );
xor \U$48369 ( \48712 , \48706 , \48711 );
xor \U$48370 ( \48713 , \48188 , \48190 );
xor \U$48371 ( \48714 , \48713 , \48197 );
and \U$48372 ( \48715 , \48712 , \48714 );
and \U$48373 ( \48716 , \48706 , \48711 );
or \U$48374 ( \48717 , \48715 , \48716 );
and \U$48375 ( \48718 , \48684 , \48717 );
and \U$48376 ( \48719 , \48436 , \48683 );
nor \U$48377 ( \48720 , \48718 , \48719 );
xor \U$48378 ( \48721 , \47943 , \47970 );
xor \U$48379 ( \48722 , \48721 , \47997 );
not \U$48380 ( \48723 , \48722 );
xor \U$48381 ( \48724 , \48107 , \48132 );
xor \U$48382 ( \48725 , \48724 , \48159 );
not \U$48383 ( \48726 , \48725 );
and \U$48384 ( \48727 , \48723 , \48726 );
and \U$48385 ( \48728 , \48725 , \48722 );
xor \U$48386 ( \48729 , \48021 , \48048 );
xor \U$48387 ( \48730 , \48729 , \48076 );
nor \U$48388 ( \48731 , \48728 , \48730 );
nor \U$48389 ( \48732 , \48727 , \48731 );
not \U$48390 ( \48733 , \48732 );
xor \U$48391 ( \48734 , \47629 , \47654 );
xor \U$48392 ( \48735 , \48734 , \47682 );
not \U$48393 ( \48736 , \48735 );
and \U$48394 ( \48737 , \48733 , \48736 );
and \U$48395 ( \48738 , \48732 , \48735 );
xor \U$48396 ( \48739 , \48254 , \48262 );
xor \U$48397 ( \48740 , \48739 , \48290 );
xor \U$48398 ( \48741 , \48212 , \48219 );
xor \U$48399 ( \48742 , \48741 , \48226 );
and \U$48400 ( \48743 , \48740 , \48742 );
xor \U$48401 ( \48744 , \48300 , \48302 );
xor \U$48402 ( \48745 , \48744 , \48305 );
xor \U$48403 ( \48746 , \48212 , \48219 );
xor \U$48404 ( \48747 , \48746 , \48226 );
and \U$48405 ( \48748 , \48745 , \48747 );
and \U$48406 ( \48749 , \48740 , \48745 );
or \U$48407 ( \48750 , \48743 , \48748 , \48749 );
not \U$48408 ( \48751 , \48750 );
nor \U$48409 ( \48752 , \48738 , \48751 );
nor \U$48410 ( \48753 , \48737 , \48752 );
xor \U$48411 ( \48754 , \48720 , \48753 );
xor \U$48412 ( \48755 , \47543 , \47569 );
xor \U$48413 ( \48756 , \48755 , \47598 );
xor \U$48414 ( \48757 , \47897 , \47902 );
xor \U$48415 ( \48758 , \48756 , \48757 );
not \U$48416 ( \48759 , \48758 );
xor \U$48417 ( \48760 , \48176 , \48181 );
xor \U$48418 ( \48761 , \48760 , \48200 );
not \U$48419 ( \48762 , \48761 );
and \U$48420 ( \48763 , \48759 , \48762 );
and \U$48421 ( \48764 , \48758 , \48761 );
xor \U$48422 ( \48765 , \47756 , \47758 );
xor \U$48423 ( \48766 , \48765 , \47761 );
xor \U$48424 ( \48767 , \47883 , \47890 );
xor \U$48425 ( \48768 , \48766 , \48767 );
nor \U$48426 ( \48769 , \48764 , \48768 );
nor \U$48427 ( \48770 , \48763 , \48769 );
and \U$48428 ( \48771 , \48754 , \48770 );
and \U$48429 ( \48772 , \48720 , \48753 );
or \U$48430 ( \48773 , \48771 , \48772 );
not \U$48431 ( \48774 , \47430 );
not \U$48432 ( \48775 , \47404 );
or \U$48433 ( \48776 , \48774 , \48775 );
or \U$48434 ( \48777 , \47404 , \47430 );
nand \U$48435 ( \48778 , \48776 , \48777 );
not \U$48436 ( \48779 , \48778 );
not \U$48437 ( \48780 , \47414 );
and \U$48438 ( \48781 , \48779 , \48780 );
and \U$48439 ( \48782 , \48778 , \47414 );
nor \U$48440 ( \48783 , \48781 , \48782 );
or \U$48441 ( \48784 , \48773 , \48783 );
not \U$48442 ( \48785 , \48783 );
not \U$48443 ( \48786 , \48773 );
or \U$48444 ( \48787 , \48785 , \48786 );
xor \U$48445 ( \48788 , \47515 , \47601 );
xor \U$48446 ( \48789 , \48788 , \47685 );
xor \U$48447 ( \48790 , \47895 , \47907 );
xor \U$48448 ( \48791 , \48790 , \47912 );
xor \U$48449 ( \48792 , \48789 , \48791 );
xor \U$48450 ( \48793 , \48324 , \48326 );
xor \U$48451 ( \48794 , \48793 , \48329 );
and \U$48452 ( \48795 , \48792 , \48794 );
and \U$48453 ( \48796 , \48789 , \48791 );
nor \U$48454 ( \48797 , \48795 , \48796 );
nand \U$48455 ( \48798 , \48787 , \48797 );
nand \U$48456 ( \48799 , \48784 , \48798 );
xor \U$48457 ( \48800 , \47827 , \47829 );
xor \U$48458 ( \48801 , \48800 , \47834 );
xor \U$48459 ( \48802 , \48799 , \48801 );
xor \U$48460 ( \48803 , \47915 , \48313 );
xor \U$48461 ( \48804 , \48803 , \48332 );
xor \U$48462 ( \48805 , \47688 , \47767 );
xor \U$48463 ( \48806 , \48805 , \47791 );
or \U$48464 ( \48807 , \48804 , \48806 );
not \U$48465 ( \48808 , \48806 );
not \U$48466 ( \48809 , \48804 );
or \U$48467 ( \48810 , \48808 , \48809 );
xor \U$48468 ( \48811 , \48347 , \48353 );
xor \U$48469 ( \48812 , \48811 , \48356 );
nand \U$48470 ( \48813 , \48810 , \48812 );
nand \U$48471 ( \48814 , \48807 , \48813 );
and \U$48472 ( \48815 , \48802 , \48814 );
and \U$48473 ( \48816 , \48799 , \48801 );
or \U$48474 ( \48817 , \48815 , \48816 );
xor \U$48475 ( \48818 , \47432 , \47794 );
xor \U$48476 ( \48819 , \48818 , \47815 );
not \U$48477 ( \48820 , \48338 );
xor \U$48478 ( \48821 , \48335 , \48359 );
not \U$48479 ( \48822 , \48821 );
or \U$48480 ( \48823 , \48820 , \48822 );
or \U$48481 ( \48824 , \48821 , \48338 );
nand \U$48482 ( \48825 , \48823 , \48824 );
and \U$48483 ( \48826 , \48819 , \48825 );
xor \U$48484 ( \48827 , \48817 , \48826 );
not \U$48485 ( \48828 , \47875 );
not \U$48486 ( \48829 , \47870 );
not \U$48487 ( \48830 , \48361 );
and \U$48488 ( \48831 , \48829 , \48830 );
and \U$48489 ( \48832 , \47870 , \48361 );
nor \U$48490 ( \48833 , \48831 , \48832 );
not \U$48491 ( \48834 , \48833 );
or \U$48492 ( \48835 , \48828 , \48834 );
or \U$48493 ( \48836 , \48833 , \47875 );
nand \U$48494 ( \48837 , \48835 , \48836 );
xor \U$48495 ( \48838 , \48827 , \48837 );
xor \U$48496 ( \48839 , \48819 , \48825 );
not \U$48497 ( \48840 , \48839 );
xor \U$48498 ( \48841 , \48799 , \48801 );
xor \U$48499 ( \48842 , \48841 , \48814 );
not \U$48500 ( \48843 , \48842 );
or \U$48501 ( \48844 , \48840 , \48843 );
or \U$48502 ( \48845 , \48842 , \48839 );
not \U$48503 ( \48846 , \48773 );
not \U$48504 ( \48847 , \48797 );
or \U$48505 ( \48848 , \48846 , \48847 );
or \U$48506 ( \48849 , \48797 , \48773 );
nand \U$48507 ( \48850 , \48848 , \48849 );
not \U$48508 ( \48851 , \48850 );
not \U$48509 ( \48852 , \48783 );
and \U$48510 ( \48853 , \48851 , \48852 );
and \U$48511 ( \48854 , \48850 , \48783 );
nor \U$48512 ( \48855 , \48853 , \48854 );
xnor \U$48513 ( \48856 , \48806 , \48804 );
not \U$48514 ( \48857 , \48856 );
not \U$48515 ( \48858 , \48812 );
and \U$48516 ( \48859 , \48857 , \48858 );
and \U$48517 ( \48860 , \48856 , \48812 );
nor \U$48518 ( \48861 , \48859 , \48860 );
or \U$48519 ( \48862 , \48855 , \48861 );
not \U$48520 ( \48863 , \48861 );
not \U$48521 ( \48864 , \48855 );
or \U$48522 ( \48865 , \48863 , \48864 );
xor \U$48523 ( \48866 , \48229 , \48293 );
xor \U$48524 ( \48867 , \48866 , \48308 );
xor \U$48525 ( \48868 , \48000 , \48079 );
xor \U$48526 ( \48869 , \48868 , \48162 );
xor \U$48527 ( \48870 , \48867 , \48869 );
not \U$48528 ( \48871 , \48761 );
xor \U$48529 ( \48872 , \48758 , \48768 );
not \U$48530 ( \48873 , \48872 );
or \U$48531 ( \48874 , \48871 , \48873 );
or \U$48532 ( \48875 , \48872 , \48761 );
nand \U$48533 ( \48876 , \48874 , \48875 );
and \U$48534 ( \48877 , \48870 , \48876 );
and \U$48535 ( \48878 , \48867 , \48869 );
or \U$48536 ( \48879 , \48877 , \48878 );
not \U$48537 ( \48880 , \48203 );
xor \U$48538 ( \48881 , \48165 , \48311 );
not \U$48539 ( \48882 , \48881 );
or \U$48540 ( \48883 , \48880 , \48882 );
or \U$48541 ( \48884 , \48881 , \48203 );
nand \U$48542 ( \48885 , \48883 , \48884 );
xor \U$48543 ( \48886 , \48879 , \48885 );
xor \U$48544 ( \48887 , \48380 , \48418 );
xor \U$48545 ( \48888 , \48887 , \48433 );
xor \U$48546 ( \48889 , \48517 , \48597 );
xor \U$48547 ( \48890 , \48889 , \48680 );
xor \U$48548 ( \48891 , \48888 , \48890 );
xor \U$48549 ( \48892 , \48706 , \48711 );
xor \U$48550 ( \48893 , \48892 , \48714 );
and \U$48551 ( \48894 , \48891 , \48893 );
and \U$48552 ( \48895 , \48888 , \48890 );
or \U$48553 ( \48896 , \48894 , \48895 );
xor \U$48554 ( \48897 , \48631 , \48638 );
xor \U$48555 ( \48898 , \48897 , \48647 );
xor \U$48556 ( \48899 , \48388 , \48396 );
xor \U$48557 ( \48900 , \48899 , \48405 );
xor \U$48558 ( \48901 , \48898 , \48900 );
xor \U$48559 ( \48902 , \48658 , \48665 );
xor \U$48560 ( \48903 , \48902 , \48674 );
and \U$48561 ( \48904 , \48901 , \48903 );
and \U$48562 ( \48905 , \48898 , \48900 );
or \U$48563 ( \48906 , \48904 , \48905 );
nand \U$48564 ( \48907 , RI9870498_86, \352 );
not \U$48565 ( \48908 , \48907 );
not \U$48566 ( \48909 , \361 );
or \U$48567 ( \48910 , \48908 , \48909 );
or \U$48568 ( \48911 , \345 , \48907 );
nand \U$48569 ( \48912 , \48910 , \48911 );
not \U$48570 ( \48913 , \487 );
and \U$48571 ( \48914 , \395 , RI9870588_88);
and \U$48572 ( \48915 , RI98703a8_84, \393 );
nor \U$48573 ( \48916 , \48914 , \48915 );
not \U$48574 ( \48917 , \48916 );
or \U$48575 ( \48918 , \48913 , \48917 );
or \U$48576 ( \48919 , \48916 , \386 );
nand \U$48577 ( \48920 , \48918 , \48919 );
and \U$48578 ( \48921 , \48912 , \48920 );
not \U$48579 ( \48922 , \345 );
and \U$48580 ( \48923 , \354 , RI9870498_86);
and \U$48581 ( \48924 , RI9870588_88, \352 );
nor \U$48582 ( \48925 , \48923 , \48924 );
not \U$48583 ( \48926 , \48925 );
or \U$48584 ( \48927 , \48922 , \48926 );
or \U$48585 ( \48928 , \48925 , \345 );
nand \U$48586 ( \48929 , \48927 , \48928 );
xor \U$48587 ( \48930 , \48921 , \48929 );
not \U$48588 ( \48931 , \365 );
and \U$48589 ( \48932 , \376 , RI98702b8_82);
and \U$48590 ( \48933 , RI9870768_92, \374 );
nor \U$48591 ( \48934 , \48932 , \48933 );
not \U$48592 ( \48935 , \48934 );
or \U$48593 ( \48936 , \48931 , \48935 );
or \U$48594 ( \48937 , \48934 , \367 );
nand \U$48595 ( \48938 , \48936 , \48937 );
and \U$48596 ( \48939 , \438 , RI9870858_94);
and \U$48597 ( \48940 , RI986fb38_66, \436 );
nor \U$48598 ( \48941 , \48939 , \48940 );
and \U$48599 ( \48942 , \48941 , \444 );
not \U$48600 ( \48943 , \48941 );
and \U$48601 ( \48944 , \48943 , \443 );
nor \U$48602 ( \48945 , \48942 , \48944 );
xor \U$48603 ( \48946 , \48938 , \48945 );
not \U$48604 ( \48947 , \456 );
and \U$48605 ( \48948 , \465 , RI9870678_90);
and \U$48606 ( \48949 , RI9870948_96, \463 );
nor \U$48607 ( \48950 , \48948 , \48949 );
not \U$48608 ( \48951 , \48950 );
or \U$48609 ( \48952 , \48947 , \48951 );
or \U$48610 ( \48953 , \48950 , \456 );
nand \U$48611 ( \48954 , \48952 , \48953 );
and \U$48612 ( \48955 , \48946 , \48954 );
and \U$48613 ( \48956 , \48938 , \48945 );
or \U$48614 ( \48957 , \48955 , \48956 );
and \U$48615 ( \48958 , \48930 , \48957 );
and \U$48616 ( \48959 , \48921 , \48929 );
or \U$48617 ( \48960 , \48958 , \48959 );
xor \U$48618 ( \48961 , \48906 , \48960 );
xor \U$48619 ( \48962 , \48605 , \48612 );
xor \U$48620 ( \48963 , \48962 , \48621 );
xor \U$48621 ( \48964 , \48496 , \48503 );
xor \U$48622 ( \48965 , \48964 , \48511 );
and \U$48623 ( \48966 , \48963 , \48965 );
xor \U$48624 ( \48967 , \48469 , \48476 );
xor \U$48625 ( \48968 , \48967 , \48485 );
xor \U$48626 ( \48969 , \48496 , \48503 );
xor \U$48627 ( \48970 , \48969 , \48511 );
and \U$48628 ( \48971 , \48968 , \48970 );
and \U$48629 ( \48972 , \48963 , \48968 );
or \U$48630 ( \48973 , \48966 , \48971 , \48972 );
and \U$48631 ( \48974 , \48961 , \48973 );
and \U$48632 ( \48975 , \48906 , \48960 );
or \U$48633 ( \48976 , \48974 , \48975 );
not \U$48634 ( \48977 , \3412 );
and \U$48635 ( \48978 , \3683 , RI98711b8_114);
and \U$48636 ( \48979 , RI9871398_118, \3681 );
nor \U$48637 ( \48980 , \48978 , \48979 );
not \U$48638 ( \48981 , \48980 );
or \U$48639 ( \48982 , \48977 , \48981 );
or \U$48640 ( \48983 , \48980 , \3412 );
nand \U$48641 ( \48984 , \48982 , \48983 );
and \U$48642 ( \48985 , \2464 , RI9870c18_102);
and \U$48643 ( \48986 , RI98710c8_112, \2462 );
nor \U$48644 ( \48987 , \48985 , \48986 );
and \U$48645 ( \48988 , \48987 , \2468 );
not \U$48646 ( \48989 , \48987 );
and \U$48647 ( \48990 , \48989 , \2263 );
nor \U$48648 ( \48991 , \48988 , \48990 );
xor \U$48649 ( \48992 , \48984 , \48991 );
not \U$48650 ( \48993 , \3406 );
and \U$48651 ( \48994 , \3254 , RI9870d08_104);
and \U$48652 ( \48995 , RI98712a8_116, \3252 );
nor \U$48653 ( \48996 , \48994 , \48995 );
not \U$48654 ( \48997 , \48996 );
or \U$48655 ( \48998 , \48993 , \48997 );
or \U$48656 ( \48999 , \48996 , \3406 );
nand \U$48657 ( \49000 , \48998 , \48999 );
and \U$48658 ( \49001 , \48992 , \49000 );
and \U$48659 ( \49002 , \48984 , \48991 );
or \U$48660 ( \49003 , \49001 , \49002 );
and \U$48661 ( \49004 , \776 , RI986fc28_68);
and \U$48662 ( \49005 , RI986fe08_72, \774 );
nor \U$48663 ( \49006 , \49004 , \49005 );
and \U$48664 ( \49007 , \49006 , \474 );
not \U$48665 ( \49008 , \49006 );
and \U$48666 ( \49009 , \49008 , \451 );
nor \U$48667 ( \49010 , \49007 , \49009 );
not \U$48668 ( \49011 , \1128 );
and \U$48669 ( \49012 , \1293 , RI986fd18_70);
and \U$48670 ( \49013 , RI986ffe8_76, \1291 );
nor \U$48671 ( \49014 , \49012 , \49013 );
not \U$48672 ( \49015 , \49014 );
or \U$48673 ( \49016 , \49011 , \49015 );
or \U$48674 ( \49017 , \49014 , \1128 );
nand \U$48675 ( \49018 , \49016 , \49017 );
xor \U$48676 ( \49019 , \49010 , \49018 );
and \U$48677 ( \49020 , \1329 , RI986fef8_74);
and \U$48678 ( \49021 , RI98700d8_78, \1327 );
nor \U$48679 ( \49022 , \49020 , \49021 );
and \U$48680 ( \49023 , \49022 , \1336 );
not \U$48681 ( \49024 , \49022 );
and \U$48682 ( \49025 , \49024 , \1337 );
nor \U$48683 ( \49026 , \49023 , \49025 );
and \U$48684 ( \49027 , \49019 , \49026 );
and \U$48685 ( \49028 , \49010 , \49018 );
or \U$48686 ( \49029 , \49027 , \49028 );
xor \U$48687 ( \49030 , \49003 , \49029 );
not \U$48688 ( \49031 , \1462 );
and \U$48689 ( \49032 , \2042 , RI9870b28_100);
and \U$48690 ( \49033 , RI9870df8_106, \2040 );
nor \U$48691 ( \49034 , \49032 , \49033 );
not \U$48692 ( \49035 , \49034 );
or \U$48693 ( \49036 , \49031 , \49035 );
or \U$48694 ( \49037 , \49034 , \2034 );
nand \U$48695 ( \49038 , \49036 , \49037 );
and \U$48696 ( \49039 , \1311 , RI98701c8_80);
and \U$48697 ( \49040 , RI9870fd8_110, \1309 );
nor \U$48698 ( \49041 , \49039 , \49040 );
and \U$48699 ( \49042 , \49041 , \1458 );
not \U$48700 ( \49043 , \49041 );
and \U$48701 ( \49044 , \49043 , \1318 );
nor \U$48702 ( \49045 , \49042 , \49044 );
xor \U$48703 ( \49046 , \49038 , \49045 );
and \U$48704 ( \49047 , \2274 , RI9870a38_98);
and \U$48705 ( \49048 , RI9870ee8_108, \2272 );
nor \U$48706 ( \49049 , \49047 , \49048 );
and \U$48707 ( \49050 , \49049 , \2030 );
not \U$48708 ( \49051 , \49049 );
and \U$48709 ( \49052 , \49051 , \2031 );
nor \U$48710 ( \49053 , \49050 , \49052 );
and \U$48711 ( \49054 , \49046 , \49053 );
and \U$48712 ( \49055 , \49038 , \49045 );
or \U$48713 ( \49056 , \49054 , \49055 );
and \U$48714 ( \49057 , \49030 , \49056 );
and \U$48715 ( \49058 , \49003 , \49029 );
or \U$48716 ( \49059 , \49057 , \49058 );
and \U$48717 ( \49060 , \9505 , RI986e4b8_18);
and \U$48718 ( \49061 , RI986e788_24, \9503 );
nor \U$48719 ( \49062 , \49060 , \49061 );
and \U$48720 ( \49063 , \49062 , \9510 );
not \U$48721 ( \49064 , \49062 );
and \U$48722 ( \49065 , \49064 , \9513 );
nor \U$48723 ( \49066 , \49063 , \49065 );
and \U$48724 ( \49067 , \10424 , RI986e698_22);
and \U$48725 ( \49068 , RI986f868_60, \10422 );
nor \U$48726 ( \49069 , \49067 , \49068 );
and \U$48727 ( \49070 , \49069 , \9840 );
not \U$48728 ( \49071 , \49069 );
and \U$48729 ( \49072 , \49071 , \10428 );
nor \U$48730 ( \49073 , \49070 , \49072 );
xor \U$48731 ( \49074 , \49066 , \49073 );
and \U$48732 ( \49075 , \11696 , RI986f778_58);
and \U$48733 ( \49076 , RI986fa48_64, \11694 );
nor \U$48734 ( \49077 , \49075 , \49076 );
and \U$48735 ( \49078 , \49077 , \10965 );
not \U$48736 ( \49079 , \49077 );
and \U$48737 ( \49080 , \49079 , \11702 );
nor \U$48738 ( \49081 , \49078 , \49080 );
and \U$48739 ( \49082 , \49074 , \49081 );
and \U$48740 ( \49083 , \49066 , \49073 );
or \U$48741 ( \49084 , \49082 , \49083 );
not \U$48742 ( \49085 , RI9873558_190);
and \U$48743 ( \49086 , \15780 , RI986dd38_2);
and \U$48744 ( \49087 , RI986e1e8_12, RI9873648_192);
nor \U$48745 ( \49088 , \49086 , \49087 );
not \U$48746 ( \49089 , \49088 );
or \U$48747 ( \49090 , \49085 , \49089 );
or \U$48748 ( \49091 , \49088 , RI9873558_190);
nand \U$48749 ( \49092 , \49090 , \49091 );
xor \U$48750 ( \49093 , \49092 , \361 );
and \U$48751 ( \49094 , \14937 , RI986df18_6);
and \U$48752 ( \49095 , RI986de28_4, \14935 );
nor \U$48753 ( \49096 , \49094 , \49095 );
and \U$48754 ( \49097 , \49096 , \14539 );
not \U$48755 ( \49098 , \49096 );
and \U$48756 ( \49099 , \49098 , \14538 );
nor \U$48757 ( \49100 , \49097 , \49099 );
and \U$48758 ( \49101 , \49093 , \49100 );
and \U$48759 ( \49102 , \49092 , \361 );
or \U$48760 ( \49103 , \49101 , \49102 );
xor \U$48761 ( \49104 , \49084 , \49103 );
and \U$48762 ( \49105 , \13882 , RI986f688_56);
and \U$48763 ( \49106 , RI986e008_8, \13880 );
nor \U$48764 ( \49107 , \49105 , \49106 );
and \U$48765 ( \49108 , \49107 , \13358 );
not \U$48766 ( \49109 , \49107 );
and \U$48767 ( \49110 , \49109 , \13359 );
nor \U$48768 ( \49111 , \49108 , \49110 );
and \U$48769 ( \49112 , \12293 , RI986f958_62);
and \U$48770 ( \49113 , RI986f4a8_52, \12291 );
nor \U$48771 ( \49114 , \49112 , \49113 );
and \U$48772 ( \49115 , \49114 , \11687 );
not \U$48773 ( \49116 , \49114 );
and \U$48774 ( \49117 , \49116 , \11686 );
nor \U$48775 ( \49118 , \49115 , \49117 );
xor \U$48776 ( \49119 , \49111 , \49118 );
and \U$48777 ( \49120 , \13045 , RI986f3b8_50);
and \U$48778 ( \49121 , RI986f598_54, \13043 );
nor \U$48779 ( \49122 , \49120 , \49121 );
and \U$48780 ( \49123 , \49122 , \13047 );
not \U$48781 ( \49124 , \49122 );
and \U$48782 ( \49125 , \49124 , \12619 );
nor \U$48783 ( \49126 , \49123 , \49125 );
and \U$48784 ( \49127 , \49119 , \49126 );
and \U$48785 ( \49128 , \49111 , \49118 );
or \U$48786 ( \49129 , \49127 , \49128 );
and \U$48787 ( \49130 , \49104 , \49129 );
and \U$48788 ( \49131 , \49084 , \49103 );
or \U$48789 ( \49132 , \49130 , \49131 );
xor \U$48790 ( \49133 , \49059 , \49132 );
and \U$48791 ( \49134 , \9237 , RI986f1d8_46);
and \U$48792 ( \49135 , RI986e5a8_20, \9235 );
nor \U$48793 ( \49136 , \49134 , \49135 );
and \U$48794 ( \49137 , \49136 , \9241 );
not \U$48795 ( \49138 , \49136 );
and \U$48796 ( \49139 , \49138 , \8836 );
nor \U$48797 ( \49140 , \49137 , \49139 );
and \U$48798 ( \49141 , \7729 , RI986ed28_36);
and \U$48799 ( \49142 , RI986f0e8_44, \7727 );
nor \U$48800 ( \49143 , \49141 , \49142 );
and \U$48801 ( \49144 , \49143 , \7480 );
not \U$48802 ( \49145 , \49143 );
and \U$48803 ( \49146 , \49145 , \7733 );
nor \U$48804 ( \49147 , \49144 , \49146 );
xor \U$48805 ( \49148 , \49140 , \49147 );
and \U$48806 ( \49149 , \8486 , RI986eff8_42);
and \U$48807 ( \49150 , RI986f2c8_48, \8484 );
nor \U$48808 ( \49151 , \49149 , \49150 );
and \U$48809 ( \49152 , \49151 , \8050 );
not \U$48810 ( \49153 , \49151 );
and \U$48811 ( \49154 , \49153 , \8051 );
nor \U$48812 ( \49155 , \49152 , \49154 );
and \U$48813 ( \49156 , \49148 , \49155 );
and \U$48814 ( \49157 , \49140 , \49147 );
or \U$48815 ( \49158 , \49156 , \49157 );
and \U$48816 ( \49159 , \5881 , RI986ea58_30);
and \U$48817 ( \49160 , RI986e968_28, \5879 );
nor \U$48818 ( \49161 , \49159 , \49160 );
and \U$48819 ( \49162 , \49161 , \5594 );
not \U$48820 ( \49163 , \49161 );
and \U$48821 ( \49164 , \49163 , \5885 );
nor \U$48822 ( \49165 , \49162 , \49164 );
and \U$48823 ( \49166 , \6453 , RI986e878_26);
and \U$48824 ( \49167 , RI986ef08_40, \6451 );
nor \U$48825 ( \49168 , \49166 , \49167 );
and \U$48826 ( \49169 , \49168 , \6190 );
not \U$48827 ( \49170 , \49168 );
and \U$48828 ( \49171 , \49170 , \6180 );
nor \U$48829 ( \49172 , \49169 , \49171 );
xor \U$48830 ( \49173 , \49165 , \49172 );
and \U$48831 ( \49174 , \7079 , RI986ee18_38);
and \U$48832 ( \49175 , RI986ec38_34, \7077 );
nor \U$48833 ( \49176 , \49174 , \49175 );
and \U$48834 ( \49177 , \49176 , \6710 );
not \U$48835 ( \49178 , \49176 );
and \U$48836 ( \49179 , \49178 , \6709 );
nor \U$48837 ( \49180 , \49177 , \49179 );
and \U$48838 ( \49181 , \49173 , \49180 );
and \U$48839 ( \49182 , \49165 , \49172 );
or \U$48840 ( \49183 , \49181 , \49182 );
xor \U$48841 ( \49184 , \49158 , \49183 );
not \U$48842 ( \49185 , \4521 );
and \U$48843 ( \49186 , \4710 , RI9871848_128);
and \U$48844 ( \49187 , RI9871578_122, \4708 );
nor \U$48845 ( \49188 , \49186 , \49187 );
not \U$48846 ( \49189 , \49188 );
or \U$48847 ( \49190 , \49185 , \49189 );
or \U$48848 ( \49191 , \49188 , \4521 );
nand \U$48849 ( \49192 , \49190 , \49191 );
and \U$48850 ( \49193 , \4203 , RI9871488_120);
and \U$48851 ( \49194 , RI9871758_126, \4201 );
nor \U$48852 ( \49195 , \49193 , \49194 );
and \U$48853 ( \49196 , \49195 , \4207 );
not \U$48854 ( \49197 , \49195 );
and \U$48855 ( \49198 , \49197 , \3923 );
nor \U$48856 ( \49199 , \49196 , \49198 );
xor \U$48857 ( \49200 , \49192 , \49199 );
and \U$48858 ( \49201 , \5318 , RI9871668_124);
and \U$48859 ( \49202 , RI986eb48_32, \5316 );
nor \U$48860 ( \49203 , \49201 , \49202 );
and \U$48861 ( \49204 , \49203 , \5052 );
not \U$48862 ( \49205 , \49203 );
and \U$48863 ( \49206 , \49205 , \5322 );
nor \U$48864 ( \49207 , \49204 , \49206 );
and \U$48865 ( \49208 , \49200 , \49207 );
and \U$48866 ( \49209 , \49192 , \49199 );
or \U$48867 ( \49210 , \49208 , \49209 );
and \U$48868 ( \49211 , \49184 , \49210 );
and \U$48869 ( \49212 , \49158 , \49183 );
or \U$48870 ( \49213 , \49211 , \49212 );
and \U$48871 ( \49214 , \49133 , \49213 );
and \U$48872 ( \49215 , \49059 , \49132 );
or \U$48873 ( \49216 , \49214 , \49215 );
xor \U$48874 ( \49217 , \48976 , \49216 );
xor \U$48875 ( \49218 , \48443 , \48450 );
xor \U$48876 ( \49219 , \49218 , \48458 );
xor \U$48877 ( \49220 , \48576 , \48583 );
xor \U$48878 ( \49221 , \49220 , \48591 );
and \U$48879 ( \49222 , \49219 , \49221 );
xor \U$48880 ( \49223 , \48524 , \48531 );
xor \U$48881 ( \49224 , \49223 , \48539 );
xor \U$48882 ( \49225 , \48576 , \48583 );
xor \U$48883 ( \49226 , \49225 , \48591 );
and \U$48884 ( \49227 , \49224 , \49226 );
and \U$48885 ( \49228 , \49219 , \49224 );
or \U$48886 ( \49229 , \49222 , \49227 , \49228 );
xor \U$48887 ( \49230 , \48690 , \48696 );
xor \U$48888 ( \49231 , \49230 , \48703 );
and \U$48889 ( \49232 , \49229 , \49231 );
xor \U$48890 ( \49233 , \48368 , \48374 );
xor \U$48891 ( \49234 , \49233 , \48377 );
xor \U$48892 ( \49235 , \48690 , \48696 );
xor \U$48893 ( \49236 , \49235 , \48703 );
and \U$48894 ( \49237 , \49234 , \49236 );
and \U$48895 ( \49238 , \49229 , \49234 );
or \U$48896 ( \49239 , \49232 , \49237 , \49238 );
and \U$48897 ( \49240 , \49217 , \49239 );
and \U$48898 ( \49241 , \48976 , \49216 );
or \U$48899 ( \49242 , \49240 , \49241 );
xor \U$48900 ( \49243 , \48896 , \49242 );
not \U$48901 ( \49244 , \48725 );
xor \U$48902 ( \49245 , \48730 , \48722 );
not \U$48903 ( \49246 , \49245 );
or \U$48904 ( \49247 , \49244 , \49246 );
or \U$48905 ( \49248 , \49245 , \48725 );
nand \U$48906 ( \49249 , \49247 , \49248 );
xor \U$48907 ( \49250 , \48237 , \48242 );
xor \U$48908 ( \49251 , \49250 , \48251 );
xor \U$48909 ( \49252 , \48408 , \48413 );
xor \U$48910 ( \49253 , \49251 , \49252 );
xor \U$48911 ( \49254 , \48624 , \48650 );
xor \U$48912 ( \49255 , \49254 , \48677 );
xor \U$48913 ( \49256 , \49253 , \49255 );
xor \U$48914 ( \49257 , \48425 , \48427 );
xor \U$48915 ( \49258 , \49257 , \48430 );
and \U$48916 ( \49259 , \49256 , \49258 );
and \U$48917 ( \49260 , \49253 , \49255 );
or \U$48918 ( \49261 , \49259 , \49260 );
xor \U$48919 ( \49262 , \49249 , \49261 );
xor \U$48920 ( \49263 , \48212 , \48219 );
xor \U$48921 ( \49264 , \49263 , \48226 );
xor \U$48922 ( \49265 , \48740 , \48745 );
xor \U$48923 ( \49266 , \49264 , \49265 );
and \U$48924 ( \49267 , \49262 , \49266 );
and \U$48925 ( \49268 , \49249 , \49261 );
or \U$48926 ( \49269 , \49267 , \49268 );
and \U$48927 ( \49270 , \49243 , \49269 );
and \U$48928 ( \49271 , \48896 , \49242 );
or \U$48929 ( \49272 , \49270 , \49271 );
and \U$48930 ( \49273 , \48886 , \49272 );
and \U$48931 ( \49274 , \48879 , \48885 );
or \U$48932 ( \49275 , \49273 , \49274 );
nand \U$48933 ( \49276 , \48865 , \49275 );
nand \U$48934 ( \49277 , \48862 , \49276 );
nand \U$48935 ( \49278 , \48845 , \49277 );
nand \U$48936 ( \49279 , \48844 , \49278 );
and \U$48937 ( \49280 , \48838 , \49279 );
xor \U$48938 ( \49281 , \49279 , \48838 );
xnor \U$48939 ( \49282 , \48842 , \49277 );
not \U$48940 ( \49283 , \49282 );
not \U$48941 ( \49284 , \48839 );
and \U$48942 ( \49285 , \49283 , \49284 );
and \U$48943 ( \49286 , \49282 , \48839 );
nor \U$48944 ( \49287 , \49285 , \49286 );
not \U$48945 ( \49288 , \49275 );
not \U$48946 ( \49289 , \48855 );
or \U$48947 ( \49290 , \49288 , \49289 );
or \U$48948 ( \49291 , \48855 , \49275 );
nand \U$48949 ( \49292 , \49290 , \49291 );
not \U$48950 ( \49293 , \49292 );
not \U$48951 ( \49294 , \48861 );
and \U$48952 ( \49295 , \49293 , \49294 );
and \U$48953 ( \49296 , \49292 , \48861 );
nor \U$48954 ( \49297 , \49295 , \49296 );
not \U$48955 ( \49298 , \49297 );
xor \U$48956 ( \49299 , \48720 , \48753 );
xor \U$48957 ( \49300 , \49299 , \48770 );
not \U$48958 ( \49301 , \49300 );
xor \U$48959 ( \49302 , \48879 , \48885 );
xor \U$48960 ( \49303 , \49302 , \49272 );
nand \U$48961 ( \49304 , \49301 , \49303 );
not \U$48962 ( \49305 , \49304 );
and \U$48963 ( \49306 , \49298 , \49305 );
and \U$48964 ( \49307 , \49297 , \49304 );
not \U$48965 ( \49308 , \48735 );
xor \U$48966 ( \49309 , \48732 , \48751 );
not \U$48967 ( \49310 , \49309 );
or \U$48968 ( \49311 , \49308 , \49310 );
or \U$48969 ( \49312 , \49309 , \48735 );
nand \U$48970 ( \49313 , \49311 , \49312 );
xor \U$48971 ( \49314 , \49084 , \49103 );
xor \U$48972 ( \49315 , \49314 , \49129 );
xor \U$48973 ( \49316 , \49003 , \49029 );
xor \U$48974 ( \49317 , \49316 , \49056 );
and \U$48975 ( \49318 , \49315 , \49317 );
xor \U$48976 ( \49319 , \49158 , \49183 );
xor \U$48977 ( \49320 , \49319 , \49210 );
xor \U$48978 ( \49321 , \49003 , \49029 );
xor \U$48979 ( \49322 , \49321 , \49056 );
and \U$48980 ( \49323 , \49320 , \49322 );
and \U$48981 ( \49324 , \49315 , \49320 );
or \U$48982 ( \49325 , \49318 , \49323 , \49324 );
xor \U$48983 ( \49326 , \48461 , \48488 );
xor \U$48984 ( \49327 , \49326 , \48514 );
xor \U$48985 ( \49328 , \49325 , \49327 );
xor \U$48986 ( \49329 , \48921 , \48929 );
xor \U$48987 ( \49330 , \49329 , \48957 );
xor \U$48988 ( \49331 , \48898 , \48900 );
xor \U$48989 ( \49332 , \49331 , \48903 );
and \U$48990 ( \49333 , \49330 , \49332 );
xor \U$48991 ( \49334 , \48496 , \48503 );
xor \U$48992 ( \49335 , \49334 , \48511 );
xor \U$48993 ( \49336 , \48963 , \48968 );
xor \U$48994 ( \49337 , \49335 , \49336 );
xor \U$48995 ( \49338 , \48898 , \48900 );
xor \U$48996 ( \49339 , \49338 , \48903 );
and \U$48997 ( \49340 , \49337 , \49339 );
and \U$48998 ( \49341 , \49330 , \49337 );
or \U$48999 ( \49342 , \49333 , \49340 , \49341 );
and \U$49000 ( \49343 , \49328 , \49342 );
and \U$49001 ( \49344 , \49325 , \49327 );
or \U$49002 ( \49345 , \49343 , \49344 );
xor \U$49003 ( \49346 , \48984 , \48991 );
xor \U$49004 ( \49347 , \49346 , \49000 );
xor \U$49005 ( \49348 , \49010 , \49018 );
xor \U$49006 ( \49349 , \49348 , \49026 );
xor \U$49007 ( \49350 , \49347 , \49349 );
xor \U$49008 ( \49351 , \49038 , \49045 );
xor \U$49009 ( \49352 , \49351 , \49053 );
and \U$49010 ( \49353 , \49350 , \49352 );
and \U$49011 ( \49354 , \49347 , \49349 );
or \U$49012 ( \49355 , \49353 , \49354 );
not \U$49013 ( \49356 , \487 );
and \U$49014 ( \49357 , \395 , RI9870498_86);
and \U$49015 ( \49358 , RI9870588_88, \393 );
nor \U$49016 ( \49359 , \49357 , \49358 );
not \U$49017 ( \49360 , \49359 );
or \U$49018 ( \49361 , \49356 , \49360 );
or \U$49019 ( \49362 , \49359 , \386 );
nand \U$49020 ( \49363 , \49361 , \49362 );
not \U$49021 ( \49364 , \456 );
and \U$49022 ( \49365 , \465 , RI9870768_92);
and \U$49023 ( \49366 , RI9870678_90, \463 );
nor \U$49024 ( \49367 , \49365 , \49366 );
not \U$49025 ( \49368 , \49367 );
or \U$49026 ( \49369 , \49364 , \49368 );
or \U$49027 ( \49370 , \49367 , \456 );
nand \U$49028 ( \49371 , \49369 , \49370 );
xor \U$49029 ( \49372 , \49363 , \49371 );
not \U$49030 ( \49373 , \365 );
and \U$49031 ( \49374 , \376 , RI98703a8_84);
and \U$49032 ( \49375 , RI98702b8_82, \374 );
nor \U$49033 ( \49376 , \49374 , \49375 );
not \U$49034 ( \49377 , \49376 );
or \U$49035 ( \49378 , \49373 , \49377 );
or \U$49036 ( \49379 , \49376 , \365 );
nand \U$49037 ( \49380 , \49378 , \49379 );
and \U$49038 ( \49381 , \49372 , \49380 );
and \U$49039 ( \49382 , \49363 , \49371 );
or \U$49040 ( \49383 , \49381 , \49382 );
xor \U$49041 ( \49384 , \48912 , \48920 );
xor \U$49042 ( \49385 , \49383 , \49384 );
xor \U$49043 ( \49386 , \48938 , \48945 );
xor \U$49044 ( \49387 , \49386 , \48954 );
and \U$49045 ( \49388 , \49385 , \49387 );
and \U$49046 ( \49389 , \49383 , \49384 );
or \U$49047 ( \49390 , \49388 , \49389 );
xor \U$49048 ( \49391 , \49355 , \49390 );
xor \U$49049 ( \49392 , \49165 , \49172 );
xor \U$49050 ( \49393 , \49392 , \49180 );
xor \U$49051 ( \49394 , \49192 , \49199 );
xor \U$49052 ( \49395 , \49394 , \49207 );
and \U$49053 ( \49396 , \49393 , \49395 );
xor \U$49054 ( \49397 , \49140 , \49147 );
xor \U$49055 ( \49398 , \49397 , \49155 );
xor \U$49056 ( \49399 , \49192 , \49199 );
xor \U$49057 ( \49400 , \49399 , \49207 );
and \U$49058 ( \49401 , \49398 , \49400 );
and \U$49059 ( \49402 , \49393 , \49398 );
or \U$49060 ( \49403 , \49396 , \49401 , \49402 );
and \U$49061 ( \49404 , \49391 , \49403 );
and \U$49062 ( \49405 , \49355 , \49390 );
or \U$49063 ( \49406 , \49404 , \49405 );
and \U$49064 ( \49407 , \8486 , RI986f0e8_44);
and \U$49065 ( \49408 , RI986eff8_42, \8484 );
nor \U$49066 ( \49409 , \49407 , \49408 );
and \U$49067 ( \49410 , \49409 , \8050 );
not \U$49068 ( \49411 , \49409 );
and \U$49069 ( \49412 , \49411 , \8051 );
nor \U$49070 ( \49413 , \49410 , \49412 );
and \U$49071 ( \49414 , \7079 , RI986ef08_40);
and \U$49072 ( \49415 , RI986ee18_38, \7077 );
nor \U$49073 ( \49416 , \49414 , \49415 );
and \U$49074 ( \49417 , \49416 , \6710 );
not \U$49075 ( \49418 , \49416 );
and \U$49076 ( \49419 , \49418 , \6709 );
nor \U$49077 ( \49420 , \49417 , \49419 );
xor \U$49078 ( \49421 , \49413 , \49420 );
and \U$49079 ( \49422 , \7729 , RI986ec38_34);
and \U$49080 ( \49423 , RI986ed28_36, \7727 );
nor \U$49081 ( \49424 , \49422 , \49423 );
and \U$49082 ( \49425 , \49424 , \7480 );
not \U$49083 ( \49426 , \49424 );
and \U$49084 ( \49427 , \49426 , \7733 );
nor \U$49085 ( \49428 , \49425 , \49427 );
and \U$49086 ( \49429 , \49421 , \49428 );
and \U$49087 ( \49430 , \49413 , \49420 );
or \U$49088 ( \49431 , \49429 , \49430 );
not \U$49089 ( \49432 , \4519 );
and \U$49090 ( \49433 , \4710 , RI9871758_126);
and \U$49091 ( \49434 , RI9871848_128, \4708 );
nor \U$49092 ( \49435 , \49433 , \49434 );
not \U$49093 ( \49436 , \49435 );
or \U$49094 ( \49437 , \49432 , \49436 );
or \U$49095 ( \49438 , \49435 , \4521 );
nand \U$49096 ( \49439 , \49437 , \49438 );
not \U$49097 ( \49440 , \3412 );
and \U$49098 ( \49441 , \3683 , RI98712a8_116);
and \U$49099 ( \49442 , RI98711b8_114, \3681 );
nor \U$49100 ( \49443 , \49441 , \49442 );
not \U$49101 ( \49444 , \49443 );
or \U$49102 ( \49445 , \49440 , \49444 );
or \U$49103 ( \49446 , \49443 , \3412 );
nand \U$49104 ( \49447 , \49445 , \49446 );
xor \U$49105 ( \49448 , \49439 , \49447 );
and \U$49106 ( \49449 , \4203 , RI9871398_118);
and \U$49107 ( \49450 , RI9871488_120, \4201 );
nor \U$49108 ( \49451 , \49449 , \49450 );
and \U$49109 ( \49452 , \49451 , \4207 );
not \U$49110 ( \49453 , \49451 );
and \U$49111 ( \49454 , \49453 , \3922 );
nor \U$49112 ( \49455 , \49452 , \49454 );
and \U$49113 ( \49456 , \49448 , \49455 );
and \U$49114 ( \49457 , \49439 , \49447 );
or \U$49115 ( \49458 , \49456 , \49457 );
xor \U$49116 ( \49459 , \49431 , \49458 );
and \U$49117 ( \49460 , \5318 , RI9871578_122);
and \U$49118 ( \49461 , RI9871668_124, \5316 );
nor \U$49119 ( \49462 , \49460 , \49461 );
and \U$49120 ( \49463 , \49462 , \5052 );
not \U$49121 ( \49464 , \49462 );
and \U$49122 ( \49465 , \49464 , \5322 );
nor \U$49123 ( \49466 , \49463 , \49465 );
and \U$49124 ( \49467 , \5881 , RI986eb48_32);
and \U$49125 ( \49468 , RI986ea58_30, \5879 );
nor \U$49126 ( \49469 , \49467 , \49468 );
and \U$49127 ( \49470 , \49469 , \5594 );
not \U$49128 ( \49471 , \49469 );
and \U$49129 ( \49472 , \49471 , \5885 );
nor \U$49130 ( \49473 , \49470 , \49472 );
xor \U$49131 ( \49474 , \49466 , \49473 );
and \U$49132 ( \49475 , \6453 , RI986e968_28);
and \U$49133 ( \49476 , RI986e878_26, \6451 );
nor \U$49134 ( \49477 , \49475 , \49476 );
and \U$49135 ( \49478 , \49477 , \6190 );
not \U$49136 ( \49479 , \49477 );
and \U$49137 ( \49480 , \49479 , \6180 );
nor \U$49138 ( \49481 , \49478 , \49480 );
and \U$49139 ( \49482 , \49474 , \49481 );
and \U$49140 ( \49483 , \49466 , \49473 );
or \U$49141 ( \49484 , \49482 , \49483 );
and \U$49142 ( \49485 , \49459 , \49484 );
and \U$49143 ( \49486 , \49431 , \49458 );
or \U$49144 ( \49487 , \49485 , \49486 );
and \U$49145 ( \49488 , \2274 , RI9870df8_106);
and \U$49146 ( \49489 , RI9870a38_98, \2272 );
nor \U$49147 ( \49490 , \49488 , \49489 );
and \U$49148 ( \49491 , \49490 , \2030 );
not \U$49149 ( \49492 , \49490 );
and \U$49150 ( \49493 , \49492 , \2031 );
nor \U$49151 ( \49494 , \49491 , \49493 );
and \U$49152 ( \49495 , \2464 , RI9870ee8_108);
and \U$49153 ( \49496 , RI9870c18_102, \2462 );
nor \U$49154 ( \49497 , \49495 , \49496 );
and \U$49155 ( \49498 , \49497 , \2468 );
not \U$49156 ( \49499 , \49497 );
and \U$49157 ( \49500 , \49499 , \2263 );
nor \U$49158 ( \49501 , \49498 , \49500 );
xor \U$49159 ( \49502 , \49494 , \49501 );
not \U$49160 ( \49503 , \2935 );
and \U$49161 ( \49504 , \3254 , RI98710c8_112);
and \U$49162 ( \49505 , RI9870d08_104, \3252 );
nor \U$49163 ( \49506 , \49504 , \49505 );
not \U$49164 ( \49507 , \49506 );
or \U$49165 ( \49508 , \49503 , \49507 );
or \U$49166 ( \49509 , \49506 , \2935 );
nand \U$49167 ( \49510 , \49508 , \49509 );
and \U$49168 ( \49511 , \49502 , \49510 );
and \U$49169 ( \49512 , \49494 , \49501 );
or \U$49170 ( \49513 , \49511 , \49512 );
and \U$49171 ( \49514 , \1329 , RI986ffe8_76);
and \U$49172 ( \49515 , RI986fef8_74, \1327 );
nor \U$49173 ( \49516 , \49514 , \49515 );
and \U$49174 ( \49517 , \49516 , \1336 );
not \U$49175 ( \49518 , \49516 );
and \U$49176 ( \49519 , \49518 , \1337 );
nor \U$49177 ( \49520 , \49517 , \49519 );
and \U$49178 ( \49521 , \1311 , RI98700d8_78);
and \U$49179 ( \49522 , RI98701c8_80, \1309 );
nor \U$49180 ( \49523 , \49521 , \49522 );
and \U$49181 ( \49524 , \49523 , \1458 );
not \U$49182 ( \49525 , \49523 );
and \U$49183 ( \49526 , \49525 , \1318 );
nor \U$49184 ( \49527 , \49524 , \49526 );
xor \U$49185 ( \49528 , \49520 , \49527 );
not \U$49186 ( \49529 , \2034 );
and \U$49187 ( \49530 , \2042 , RI9870fd8_110);
and \U$49188 ( \49531 , RI9870b28_100, \2040 );
nor \U$49189 ( \49532 , \49530 , \49531 );
not \U$49190 ( \49533 , \49532 );
or \U$49191 ( \49534 , \49529 , \49533 );
or \U$49192 ( \49535 , \49532 , \2034 );
nand \U$49193 ( \49536 , \49534 , \49535 );
and \U$49194 ( \49537 , \49528 , \49536 );
and \U$49195 ( \49538 , \49520 , \49527 );
or \U$49196 ( \49539 , \49537 , \49538 );
xor \U$49197 ( \49540 , \49513 , \49539 );
and \U$49198 ( \49541 , \776 , RI986fb38_66);
and \U$49199 ( \49542 , RI986fc28_68, \774 );
nor \U$49200 ( \49543 , \49541 , \49542 );
and \U$49201 ( \49544 , \49543 , \474 );
not \U$49202 ( \49545 , \49543 );
and \U$49203 ( \49546 , \49545 , \451 );
nor \U$49204 ( \49547 , \49544 , \49546 );
and \U$49205 ( \49548 , \438 , RI9870948_96);
and \U$49206 ( \49549 , RI9870858_94, \436 );
nor \U$49207 ( \49550 , \49548 , \49549 );
and \U$49208 ( \49551 , \49550 , \444 );
not \U$49209 ( \49552 , \49550 );
and \U$49210 ( \49553 , \49552 , \443 );
nor \U$49211 ( \49554 , \49551 , \49553 );
xor \U$49212 ( \49555 , \49547 , \49554 );
not \U$49213 ( \49556 , \1128 );
and \U$49214 ( \49557 , \1293 , RI986fe08_72);
and \U$49215 ( \49558 , RI986fd18_70, \1291 );
nor \U$49216 ( \49559 , \49557 , \49558 );
not \U$49217 ( \49560 , \49559 );
or \U$49218 ( \49561 , \49556 , \49560 );
or \U$49219 ( \49562 , \49559 , \1128 );
nand \U$49220 ( \49563 , \49561 , \49562 );
and \U$49221 ( \49564 , \49555 , \49563 );
and \U$49222 ( \49565 , \49547 , \49554 );
or \U$49223 ( \49566 , \49564 , \49565 );
and \U$49224 ( \49567 , \49540 , \49566 );
and \U$49225 ( \49568 , \49513 , \49539 );
or \U$49226 ( \49569 , \49567 , \49568 );
xor \U$49227 ( \49570 , \49487 , \49569 );
and \U$49228 ( \49571 , \9237 , RI986f2c8_48);
and \U$49229 ( \49572 , RI986f1d8_46, \9235 );
nor \U$49230 ( \49573 , \49571 , \49572 );
and \U$49231 ( \49574 , \49573 , \9241 );
not \U$49232 ( \49575 , \49573 );
and \U$49233 ( \49576 , \49575 , \8836 );
nor \U$49234 ( \49577 , \49574 , \49576 );
and \U$49235 ( \49578 , \9505 , RI986e5a8_20);
and \U$49236 ( \49579 , RI986e4b8_18, \9503 );
nor \U$49237 ( \49580 , \49578 , \49579 );
and \U$49238 ( \49581 , \49580 , \9510 );
not \U$49239 ( \49582 , \49580 );
and \U$49240 ( \49583 , \49582 , \9513 );
nor \U$49241 ( \49584 , \49581 , \49583 );
xor \U$49242 ( \49585 , \49577 , \49584 );
and \U$49243 ( \49586 , \10424 , RI986e788_24);
and \U$49244 ( \49587 , RI986e698_22, \10422 );
nor \U$49245 ( \49588 , \49586 , \49587 );
and \U$49246 ( \49589 , \49588 , \9840 );
not \U$49247 ( \49590 , \49588 );
and \U$49248 ( \49591 , \49590 , \10428 );
nor \U$49249 ( \49592 , \49589 , \49591 );
and \U$49250 ( \49593 , \49585 , \49592 );
and \U$49251 ( \49594 , \49577 , \49584 );
or \U$49252 ( \49595 , \49593 , \49594 );
and \U$49253 ( \49596 , \14937 , RI986e008_8);
and \U$49254 ( \49597 , RI986df18_6, \14935 );
nor \U$49255 ( \49598 , \49596 , \49597 );
and \U$49256 ( \49599 , \49598 , \14539 );
not \U$49257 ( \49600 , \49598 );
and \U$49258 ( \49601 , \49600 , \14538 );
nor \U$49259 ( \49602 , \49599 , \49601 );
not \U$49260 ( \49603 , RI9873558_190);
and \U$49261 ( \49604 , \15780 , RI986de28_4);
and \U$49262 ( \49605 , RI986dd38_2, RI9873648_192);
nor \U$49263 ( \49606 , \49604 , \49605 );
not \U$49264 ( \49607 , \49606 );
or \U$49265 ( \49608 , \49603 , \49607 );
or \U$49266 ( \49609 , \49606 , RI9873558_190);
nand \U$49267 ( \49610 , \49608 , \49609 );
xor \U$49268 ( \49611 , \49602 , \49610 );
and \U$49269 ( \49612 , \13882 , RI986f598_54);
and \U$49270 ( \49613 , RI986f688_56, \13880 );
nor \U$49271 ( \49614 , \49612 , \49613 );
and \U$49272 ( \49615 , \49614 , \13358 );
not \U$49273 ( \49616 , \49614 );
and \U$49274 ( \49617 , \49616 , \13359 );
nor \U$49275 ( \49618 , \49615 , \49617 );
and \U$49276 ( \49619 , \49611 , \49618 );
and \U$49277 ( \49620 , \49602 , \49610 );
or \U$49278 ( \49621 , \49619 , \49620 );
xor \U$49279 ( \49622 , \49595 , \49621 );
and \U$49280 ( \49623 , \13045 , RI986f4a8_52);
and \U$49281 ( \49624 , RI986f3b8_50, \13043 );
nor \U$49282 ( \49625 , \49623 , \49624 );
and \U$49283 ( \49626 , \49625 , \13047 );
not \U$49284 ( \49627 , \49625 );
and \U$49285 ( \49628 , \49627 , \12619 );
nor \U$49286 ( \49629 , \49626 , \49628 );
and \U$49287 ( \49630 , \11696 , RI986f868_60);
and \U$49288 ( \49631 , RI986f778_58, \11694 );
nor \U$49289 ( \49632 , \49630 , \49631 );
and \U$49290 ( \49633 , \49632 , \10965 );
not \U$49291 ( \49634 , \49632 );
and \U$49292 ( \49635 , \49634 , \11702 );
nor \U$49293 ( \49636 , \49633 , \49635 );
xor \U$49294 ( \49637 , \49629 , \49636 );
and \U$49295 ( \49638 , \12293 , RI986fa48_64);
and \U$49296 ( \49639 , RI986f958_62, \12291 );
nor \U$49297 ( \49640 , \49638 , \49639 );
and \U$49298 ( \49641 , \49640 , \11687 );
not \U$49299 ( \49642 , \49640 );
and \U$49300 ( \49643 , \49642 , \11686 );
nor \U$49301 ( \49644 , \49641 , \49643 );
and \U$49302 ( \49645 , \49637 , \49644 );
and \U$49303 ( \49646 , \49629 , \49636 );
or \U$49304 ( \49647 , \49645 , \49646 );
and \U$49305 ( \49648 , \49622 , \49647 );
and \U$49306 ( \49649 , \49595 , \49621 );
or \U$49307 ( \49650 , \49648 , \49649 );
and \U$49308 ( \49651 , \49570 , \49650 );
and \U$49309 ( \49652 , \49487 , \49569 );
or \U$49310 ( \49653 , \49651 , \49652 );
xor \U$49311 ( \49654 , \49406 , \49653 );
xor \U$49312 ( \49655 , \49092 , \361 );
xor \U$49313 ( \49656 , \49655 , \49100 );
xor \U$49314 ( \49657 , \49111 , \49118 );
xor \U$49315 ( \49658 , \49657 , \49126 );
and \U$49316 ( \49659 , \49656 , \49658 );
xor \U$49317 ( \49660 , \49066 , \49073 );
xor \U$49318 ( \49661 , \49660 , \49081 );
xor \U$49319 ( \49662 , \49111 , \49118 );
xor \U$49320 ( \49663 , \49662 , \49126 );
and \U$49321 ( \49664 , \49661 , \49663 );
and \U$49322 ( \49665 , \49656 , \49661 );
or \U$49323 ( \49666 , \49659 , \49664 , \49665 );
xor \U$49324 ( \49667 , \48549 , \48557 );
xor \U$49325 ( \49668 , \49667 , \48565 );
xor \U$49326 ( \49669 , \49666 , \49668 );
xor \U$49327 ( \49670 , \48576 , \48583 );
xor \U$49328 ( \49671 , \49670 , \48591 );
xor \U$49329 ( \49672 , \49219 , \49224 );
xor \U$49330 ( \49673 , \49671 , \49672 );
and \U$49331 ( \49674 , \49669 , \49673 );
and \U$49332 ( \49675 , \49666 , \49668 );
or \U$49333 ( \49676 , \49674 , \49675 );
and \U$49334 ( \49677 , \49654 , \49676 );
and \U$49335 ( \49678 , \49406 , \49653 );
or \U$49336 ( \49679 , \49677 , \49678 );
xor \U$49337 ( \49680 , \49345 , \49679 );
xor \U$49338 ( \49681 , \48542 , \48568 );
xor \U$49339 ( \49682 , \49681 , \48594 );
xor \U$49340 ( \49683 , \49253 , \49255 );
xor \U$49341 ( \49684 , \49683 , \49258 );
and \U$49342 ( \49685 , \49682 , \49684 );
xor \U$49343 ( \49686 , \48690 , \48696 );
xor \U$49344 ( \49687 , \49686 , \48703 );
xor \U$49345 ( \49688 , \49229 , \49234 );
xor \U$49346 ( \49689 , \49687 , \49688 );
xor \U$49347 ( \49690 , \49253 , \49255 );
xor \U$49348 ( \49691 , \49690 , \49258 );
and \U$49349 ( \49692 , \49689 , \49691 );
and \U$49350 ( \49693 , \49682 , \49689 );
or \U$49351 ( \49694 , \49685 , \49692 , \49693 );
and \U$49352 ( \49695 , \49680 , \49694 );
and \U$49353 ( \49696 , \49345 , \49679 );
or \U$49354 ( \49697 , \49695 , \49696 );
xor \U$49355 ( \49698 , \49313 , \49697 );
xor \U$49356 ( \49699 , \48976 , \49216 );
xor \U$49357 ( \49700 , \49699 , \49239 );
xor \U$49358 ( \49701 , \48888 , \48890 );
xor \U$49359 ( \49702 , \49701 , \48893 );
and \U$49360 ( \49703 , \49700 , \49702 );
xor \U$49361 ( \49704 , \49249 , \49261 );
xor \U$49362 ( \49705 , \49704 , \49266 );
xor \U$49363 ( \49706 , \48888 , \48890 );
xor \U$49364 ( \49707 , \49706 , \48893 );
and \U$49365 ( \49708 , \49705 , \49707 );
and \U$49366 ( \49709 , \49700 , \49705 );
or \U$49367 ( \49710 , \49703 , \49708 , \49709 );
and \U$49368 ( \49711 , \49698 , \49710 );
and \U$49369 ( \49712 , \49313 , \49697 );
nor \U$49370 ( \49713 , \49711 , \49712 );
not \U$49371 ( \49714 , \49713 );
xor \U$49372 ( \49715 , \48789 , \48791 );
xor \U$49373 ( \49716 , \49715 , \48794 );
not \U$49374 ( \49717 , \49716 );
and \U$49375 ( \49718 , \49714 , \49717 );
and \U$49376 ( \49719 , \49713 , \49716 );
xor \U$49377 ( \49720 , \48867 , \48869 );
xor \U$49378 ( \49721 , \49720 , \48876 );
xor \U$49379 ( \49722 , \48896 , \49242 );
xor \U$49380 ( \49723 , \49722 , \49269 );
xor \U$49381 ( \49724 , \49721 , \49723 );
xor \U$49382 ( \49725 , \48436 , \48683 );
xor \U$49383 ( \49726 , \49725 , \48717 );
and \U$49384 ( \49727 , \49724 , \49726 );
and \U$49385 ( \49728 , \49721 , \49723 );
nor \U$49386 ( \49729 , \49727 , \49728 );
nor \U$49387 ( \49730 , \49719 , \49729 );
nor \U$49388 ( \49731 , \49718 , \49730 );
nor \U$49389 ( \49732 , \49307 , \49731 );
nor \U$49390 ( \49733 , \49306 , \49732 );
or \U$49391 ( \49734 , \49287 , \49733 );
xnor \U$49392 ( \49735 , \49733 , \49287 );
not \U$49393 ( \49736 , \49297 );
xor \U$49394 ( \49737 , \49304 , \49731 );
not \U$49395 ( \49738 , \49737 );
or \U$49396 ( \49739 , \49736 , \49738 );
or \U$49397 ( \49740 , \49737 , \49297 );
nand \U$49398 ( \49741 , \49739 , \49740 );
xor \U$49399 ( \49742 , \49721 , \49723 );
xor \U$49400 ( \49743 , \49742 , \49726 );
xor \U$49401 ( \49744 , \49003 , \49029 );
xor \U$49402 ( \49745 , \49744 , \49056 );
xor \U$49403 ( \49746 , \49315 , \49320 );
xor \U$49404 ( \49747 , \49745 , \49746 );
xor \U$49405 ( \49748 , \49513 , \49539 );
xor \U$49406 ( \49749 , \49748 , \49566 );
xor \U$49407 ( \49750 , \49431 , \49458 );
xor \U$49408 ( \49751 , \49750 , \49484 );
and \U$49409 ( \49752 , \49749 , \49751 );
xor \U$49410 ( \49753 , \49383 , \49384 );
xor \U$49411 ( \49754 , \49753 , \49387 );
xor \U$49412 ( \49755 , \49431 , \49458 );
xor \U$49413 ( \49756 , \49755 , \49484 );
and \U$49414 ( \49757 , \49754 , \49756 );
and \U$49415 ( \49758 , \49749 , \49754 );
or \U$49416 ( \49759 , \49752 , \49757 , \49758 );
xor \U$49417 ( \49760 , \49747 , \49759 );
xor \U$49418 ( \49761 , \48898 , \48900 );
xor \U$49419 ( \49762 , \49761 , \48903 );
xor \U$49420 ( \49763 , \49330 , \49337 );
xor \U$49421 ( \49764 , \49762 , \49763 );
and \U$49422 ( \49765 , \49760 , \49764 );
and \U$49423 ( \49766 , \49747 , \49759 );
or \U$49424 ( \49767 , \49765 , \49766 );
xor \U$49425 ( \49768 , \49466 , \49473 );
xor \U$49426 ( \49769 , \49768 , \49481 );
xor \U$49427 ( \49770 , \49413 , \49420 );
xor \U$49428 ( \49771 , \49770 , \49428 );
and \U$49429 ( \49772 , \49769 , \49771 );
xor \U$49430 ( \49773 , \49577 , \49584 );
xor \U$49431 ( \49774 , \49773 , \49592 );
xor \U$49432 ( \49775 , \49413 , \49420 );
xor \U$49433 ( \49776 , \49775 , \49428 );
and \U$49434 ( \49777 , \49774 , \49776 );
and \U$49435 ( \49778 , \49769 , \49774 );
or \U$49436 ( \49779 , \49772 , \49777 , \49778 );
xor \U$49437 ( \49780 , \49363 , \49371 );
xor \U$49438 ( \49781 , \49780 , \49380 );
not \U$49439 ( \49782 , \365 );
and \U$49440 ( \49783 , \376 , RI9870588_88);
and \U$49441 ( \49784 , RI98703a8_84, \374 );
nor \U$49442 ( \49785 , \49783 , \49784 );
not \U$49443 ( \49786 , \49785 );
or \U$49444 ( \49787 , \49782 , \49786 );
or \U$49445 ( \49788 , \49785 , \367 );
nand \U$49446 ( \49789 , \49787 , \49788 );
and \U$49447 ( \49790 , \438 , RI9870678_90);
and \U$49448 ( \49791 , RI9870948_96, \436 );
nor \U$49449 ( \49792 , \49790 , \49791 );
and \U$49450 ( \49793 , \49792 , \444 );
not \U$49451 ( \49794 , \49792 );
and \U$49452 ( \49795 , \49794 , \443 );
nor \U$49453 ( \49796 , \49793 , \49795 );
xor \U$49454 ( \49797 , \49789 , \49796 );
not \U$49455 ( \49798 , \454 );
and \U$49456 ( \49799 , \465 , RI98702b8_82);
and \U$49457 ( \49800 , RI9870768_92, \463 );
nor \U$49458 ( \49801 , \49799 , \49800 );
not \U$49459 ( \49802 , \49801 );
or \U$49460 ( \49803 , \49798 , \49802 );
or \U$49461 ( \49804 , \49801 , \456 );
nand \U$49462 ( \49805 , \49803 , \49804 );
and \U$49463 ( \49806 , \49797 , \49805 );
and \U$49464 ( \49807 , \49789 , \49796 );
or \U$49465 ( \49808 , \49806 , \49807 );
xor \U$49466 ( \49809 , \49781 , \49808 );
xor \U$49467 ( \49810 , \49547 , \49554 );
xor \U$49468 ( \49811 , \49810 , \49563 );
and \U$49469 ( \49812 , \49809 , \49811 );
and \U$49470 ( \49813 , \49781 , \49808 );
or \U$49471 ( \49814 , \49812 , \49813 );
xor \U$49472 ( \49815 , \49779 , \49814 );
xor \U$49473 ( \49816 , \49520 , \49527 );
xor \U$49474 ( \49817 , \49816 , \49536 );
xor \U$49475 ( \49818 , \49494 , \49501 );
xor \U$49476 ( \49819 , \49818 , \49510 );
and \U$49477 ( \49820 , \49817 , \49819 );
xor \U$49478 ( \49821 , \49439 , \49447 );
xor \U$49479 ( \49822 , \49821 , \49455 );
xor \U$49480 ( \49823 , \49494 , \49501 );
xor \U$49481 ( \49824 , \49823 , \49510 );
and \U$49482 ( \49825 , \49822 , \49824 );
and \U$49483 ( \49826 , \49817 , \49822 );
or \U$49484 ( \49827 , \49820 , \49825 , \49826 );
and \U$49485 ( \49828 , \49815 , \49827 );
and \U$49486 ( \49829 , \49779 , \49814 );
or \U$49487 ( \49830 , \49828 , \49829 );
not \U$49488 ( \49831 , \3406 );
and \U$49489 ( \49832 , \3254 , RI9870c18_102);
and \U$49490 ( \49833 , RI98710c8_112, \3252 );
nor \U$49491 ( \49834 , \49832 , \49833 );
not \U$49492 ( \49835 , \49834 );
or \U$49493 ( \49836 , \49831 , \49835 );
or \U$49494 ( \49837 , \49834 , \2935 );
nand \U$49495 ( \49838 , \49836 , \49837 );
and \U$49496 ( \49839 , \2464 , RI9870a38_98);
and \U$49497 ( \49840 , RI9870ee8_108, \2462 );
nor \U$49498 ( \49841 , \49839 , \49840 );
and \U$49499 ( \49842 , \49841 , \2468 );
not \U$49500 ( \49843 , \49841 );
and \U$49501 ( \49844 , \49843 , \2263 );
nor \U$49502 ( \49845 , \49842 , \49844 );
xor \U$49503 ( \49846 , \49838 , \49845 );
not \U$49504 ( \49847 , \3918 );
and \U$49505 ( \49848 , \3683 , RI9870d08_104);
and \U$49506 ( \49849 , RI98712a8_116, \3681 );
nor \U$49507 ( \49850 , \49848 , \49849 );
not \U$49508 ( \49851 , \49850 );
or \U$49509 ( \49852 , \49847 , \49851 );
or \U$49510 ( \49853 , \49850 , \3918 );
nand \U$49511 ( \49854 , \49852 , \49853 );
and \U$49512 ( \49855 , \49846 , \49854 );
and \U$49513 ( \49856 , \49838 , \49845 );
or \U$49514 ( \49857 , \49855 , \49856 );
and \U$49515 ( \49858 , \1329 , RI986fd18_70);
and \U$49516 ( \49859 , RI986ffe8_76, \1327 );
nor \U$49517 ( \49860 , \49858 , \49859 );
and \U$49518 ( \49861 , \49860 , \1336 );
not \U$49519 ( \49862 , \49860 );
and \U$49520 ( \49863 , \49862 , \1337 );
nor \U$49521 ( \49864 , \49861 , \49863 );
and \U$49522 ( \49865 , \776 , RI9870858_94);
and \U$49523 ( \49866 , RI986fb38_66, \774 );
nor \U$49524 ( \49867 , \49865 , \49866 );
and \U$49525 ( \49868 , \49867 , \474 );
not \U$49526 ( \49869 , \49867 );
and \U$49527 ( \49870 , \49869 , \451 );
nor \U$49528 ( \49871 , \49868 , \49870 );
xor \U$49529 ( \49872 , \49864 , \49871 );
not \U$49530 ( \49873 , \1301 );
and \U$49531 ( \49874 , \1293 , RI986fc28_68);
and \U$49532 ( \49875 , RI986fe08_72, \1291 );
nor \U$49533 ( \49876 , \49874 , \49875 );
not \U$49534 ( \49877 , \49876 );
or \U$49535 ( \49878 , \49873 , \49877 );
or \U$49536 ( \49879 , \49876 , \1301 );
nand \U$49537 ( \49880 , \49878 , \49879 );
and \U$49538 ( \49881 , \49872 , \49880 );
and \U$49539 ( \49882 , \49864 , \49871 );
or \U$49540 ( \49883 , \49881 , \49882 );
xor \U$49541 ( \49884 , \49857 , \49883 );
not \U$49542 ( \49885 , \1462 );
and \U$49543 ( \49886 , \2042 , RI98701c8_80);
and \U$49544 ( \49887 , RI9870fd8_110, \2040 );
nor \U$49545 ( \49888 , \49886 , \49887 );
not \U$49546 ( \49889 , \49888 );
or \U$49547 ( \49890 , \49885 , \49889 );
or \U$49548 ( \49891 , \49888 , \2034 );
nand \U$49549 ( \49892 , \49890 , \49891 );
and \U$49550 ( \49893 , \1311 , RI986fef8_74);
and \U$49551 ( \49894 , RI98700d8_78, \1309 );
nor \U$49552 ( \49895 , \49893 , \49894 );
and \U$49553 ( \49896 , \49895 , \1458 );
not \U$49554 ( \49897 , \49895 );
and \U$49555 ( \49898 , \49897 , \1315 );
nor \U$49556 ( \49899 , \49896 , \49898 );
xor \U$49557 ( \49900 , \49892 , \49899 );
and \U$49558 ( \49901 , \2274 , RI9870b28_100);
and \U$49559 ( \49902 , RI9870df8_106, \2272 );
nor \U$49560 ( \49903 , \49901 , \49902 );
and \U$49561 ( \49904 , \49903 , \2030 );
not \U$49562 ( \49905 , \49903 );
and \U$49563 ( \49906 , \49905 , \2031 );
nor \U$49564 ( \49907 , \49904 , \49906 );
and \U$49565 ( \49908 , \49900 , \49907 );
and \U$49566 ( \49909 , \49892 , \49899 );
or \U$49567 ( \49910 , \49908 , \49909 );
and \U$49568 ( \49911 , \49884 , \49910 );
and \U$49569 ( \49912 , \49857 , \49883 );
or \U$49570 ( \49913 , \49911 , \49912 );
and \U$49571 ( \49914 , \9505 , RI986f1d8_46);
and \U$49572 ( \49915 , RI986e5a8_20, \9503 );
nor \U$49573 ( \49916 , \49914 , \49915 );
and \U$49574 ( \49917 , \49916 , \9510 );
not \U$49575 ( \49918 , \49916 );
and \U$49576 ( \49919 , \49918 , \9513 );
nor \U$49577 ( \49920 , \49917 , \49919 );
and \U$49578 ( \49921 , \10424 , RI986e4b8_18);
and \U$49579 ( \49922 , RI986e788_24, \10422 );
nor \U$49580 ( \49923 , \49921 , \49922 );
and \U$49581 ( \49924 , \49923 , \9840 );
not \U$49582 ( \49925 , \49923 );
and \U$49583 ( \49926 , \49925 , \10428 );
nor \U$49584 ( \49927 , \49924 , \49926 );
xor \U$49585 ( \49928 , \49920 , \49927 );
and \U$49586 ( \49929 , \11696 , RI986e698_22);
and \U$49587 ( \49930 , RI986f868_60, \11694 );
nor \U$49588 ( \49931 , \49929 , \49930 );
and \U$49589 ( \49932 , \49931 , \10965 );
not \U$49590 ( \49933 , \49931 );
and \U$49591 ( \49934 , \49933 , \11702 );
nor \U$49592 ( \49935 , \49932 , \49934 );
and \U$49593 ( \49936 , \49928 , \49935 );
and \U$49594 ( \49937 , \49920 , \49927 );
or \U$49595 ( \49938 , \49936 , \49937 );
not \U$49596 ( \49939 , RI9873558_190);
and \U$49597 ( \49940 , \15780 , RI986df18_6);
and \U$49598 ( \49941 , RI986de28_4, RI9873648_192);
nor \U$49599 ( \49942 , \49940 , \49941 );
not \U$49600 ( \49943 , \49942 );
or \U$49601 ( \49944 , \49939 , \49943 );
or \U$49602 ( \49945 , \49942 , RI9873558_190);
nand \U$49603 ( \49946 , \49944 , \49945 );
xor \U$49604 ( \49947 , \49946 , \487 );
and \U$49605 ( \49948 , \14937 , RI986f688_56);
and \U$49606 ( \49949 , RI986e008_8, \14935 );
nor \U$49607 ( \49950 , \49948 , \49949 );
and \U$49608 ( \49951 , \49950 , \14539 );
not \U$49609 ( \49952 , \49950 );
and \U$49610 ( \49953 , \49952 , \14538 );
nor \U$49611 ( \49954 , \49951 , \49953 );
and \U$49612 ( \49955 , \49947 , \49954 );
and \U$49613 ( \49956 , \49946 , \487 );
or \U$49614 ( \49957 , \49955 , \49956 );
xor \U$49615 ( \49958 , \49938 , \49957 );
and \U$49616 ( \49959 , \13882 , RI986f3b8_50);
and \U$49617 ( \49960 , RI986f598_54, \13880 );
nor \U$49618 ( \49961 , \49959 , \49960 );
and \U$49619 ( \49962 , \49961 , \13358 );
not \U$49620 ( \49963 , \49961 );
and \U$49621 ( \49964 , \49963 , \13359 );
nor \U$49622 ( \49965 , \49962 , \49964 );
and \U$49623 ( \49966 , \12293 , RI986f778_58);
and \U$49624 ( \49967 , RI986fa48_64, \12291 );
nor \U$49625 ( \49968 , \49966 , \49967 );
and \U$49626 ( \49969 , \49968 , \11687 );
not \U$49627 ( \49970 , \49968 );
and \U$49628 ( \49971 , \49970 , \11686 );
nor \U$49629 ( \49972 , \49969 , \49971 );
xor \U$49630 ( \49973 , \49965 , \49972 );
and \U$49631 ( \49974 , \13045 , RI986f958_62);
and \U$49632 ( \49975 , RI986f4a8_52, \13043 );
nor \U$49633 ( \49976 , \49974 , \49975 );
and \U$49634 ( \49977 , \49976 , \13047 );
not \U$49635 ( \49978 , \49976 );
and \U$49636 ( \49979 , \49978 , \12619 );
nor \U$49637 ( \49980 , \49977 , \49979 );
and \U$49638 ( \49981 , \49973 , \49980 );
and \U$49639 ( \49982 , \49965 , \49972 );
or \U$49640 ( \49983 , \49981 , \49982 );
and \U$49641 ( \49984 , \49958 , \49983 );
and \U$49642 ( \49985 , \49938 , \49957 );
or \U$49643 ( \49986 , \49984 , \49985 );
xor \U$49644 ( \49987 , \49913 , \49986 );
and \U$49645 ( \49988 , \4203 , RI98711b8_114);
and \U$49646 ( \49989 , RI9871398_118, \4201 );
nor \U$49647 ( \49990 , \49988 , \49989 );
and \U$49648 ( \49991 , \49990 , \3923 );
not \U$49649 ( \49992 , \49990 );
and \U$49650 ( \49993 , \49992 , \4207 );
nor \U$49651 ( \49994 , \49991 , \49993 );
not \U$49652 ( \49995 , \49994 );
and \U$49653 ( \49996 , \4710 , RI9871488_120);
and \U$49654 ( \49997 , RI9871758_126, \4708 );
nor \U$49655 ( \49998 , \49996 , \49997 );
not \U$49656 ( \49999 , \49998 );
not \U$49657 ( \50000 , \4521 );
and \U$49658 ( \50001 , \49999 , \50000 );
and \U$49659 ( \50002 , \49998 , \4519 );
nor \U$49660 ( \50003 , \50001 , \50002 );
not \U$49661 ( \50004 , \50003 );
and \U$49662 ( \50005 , \49995 , \50004 );
and \U$49663 ( \50006 , \50003 , \49994 );
and \U$49664 ( \50007 , \5318 , RI9871848_128);
and \U$49665 ( \50008 , RI9871578_122, \5316 );
nor \U$49666 ( \50009 , \50007 , \50008 );
and \U$49667 ( \50010 , \50009 , \5322 );
not \U$49668 ( \50011 , \50009 );
and \U$49669 ( \50012 , \50011 , \5052 );
nor \U$49670 ( \50013 , \50010 , \50012 );
nor \U$49671 ( \50014 , \50006 , \50013 );
nor \U$49672 ( \50015 , \50005 , \50014 );
and \U$49673 ( \50016 , \7729 , RI986ee18_38);
and \U$49674 ( \50017 , RI986ec38_34, \7727 );
nor \U$49675 ( \50018 , \50016 , \50017 );
and \U$49676 ( \50019 , \50018 , \7733 );
not \U$49677 ( \50020 , \50018 );
and \U$49678 ( \50021 , \50020 , \7480 );
nor \U$49679 ( \50022 , \50019 , \50021 );
not \U$49680 ( \50023 , \50022 );
and \U$49681 ( \50024 , \8486 , RI986ed28_36);
and \U$49682 ( \50025 , RI986f0e8_44, \8484 );
nor \U$49683 ( \50026 , \50024 , \50025 );
and \U$49684 ( \50027 , \50026 , \8051 );
not \U$49685 ( \50028 , \50026 );
and \U$49686 ( \50029 , \50028 , \8050 );
nor \U$49687 ( \50030 , \50027 , \50029 );
not \U$49688 ( \50031 , \50030 );
and \U$49689 ( \50032 , \50023 , \50031 );
and \U$49690 ( \50033 , \50030 , \50022 );
and \U$49691 ( \50034 , \9237 , RI986eff8_42);
and \U$49692 ( \50035 , RI986f2c8_48, \9235 );
nor \U$49693 ( \50036 , \50034 , \50035 );
and \U$49694 ( \50037 , \50036 , \8836 );
not \U$49695 ( \50038 , \50036 );
and \U$49696 ( \50039 , \50038 , \9241 );
nor \U$49697 ( \50040 , \50037 , \50039 );
nor \U$49698 ( \50041 , \50033 , \50040 );
nor \U$49699 ( \50042 , \50032 , \50041 );
or \U$49700 ( \50043 , \50015 , \50042 );
not \U$49701 ( \50044 , \50015 );
not \U$49702 ( \50045 , \50042 );
or \U$49703 ( \50046 , \50044 , \50045 );
and \U$49704 ( \50047 , \6453 , RI986ea58_30);
and \U$49705 ( \50048 , RI986e968_28, \6451 );
nor \U$49706 ( \50049 , \50047 , \50048 );
and \U$49707 ( \50050 , \50049 , \6190 );
not \U$49708 ( \50051 , \50049 );
and \U$49709 ( \50052 , \50051 , \6705 );
nor \U$49710 ( \50053 , \50050 , \50052 );
and \U$49711 ( \50054 , \5881 , RI9871668_124);
and \U$49712 ( \50055 , RI986eb48_32, \5879 );
nor \U$49713 ( \50056 , \50054 , \50055 );
and \U$49714 ( \50057 , \50056 , \5594 );
not \U$49715 ( \50058 , \50056 );
and \U$49716 ( \50059 , \50058 , \5885 );
nor \U$49717 ( \50060 , \50057 , \50059 );
xor \U$49718 ( \50061 , \50053 , \50060 );
and \U$49719 ( \50062 , \7079 , RI986e878_26);
and \U$49720 ( \50063 , RI986ef08_40, \7077 );
nor \U$49721 ( \50064 , \50062 , \50063 );
and \U$49722 ( \50065 , \50064 , \6710 );
not \U$49723 ( \50066 , \50064 );
and \U$49724 ( \50067 , \50066 , \6709 );
nor \U$49725 ( \50068 , \50065 , \50067 );
and \U$49726 ( \50069 , \50061 , \50068 );
and \U$49727 ( \50070 , \50053 , \50060 );
or \U$49728 ( \50071 , \50069 , \50070 );
nand \U$49729 ( \50072 , \50046 , \50071 );
nand \U$49730 ( \50073 , \50043 , \50072 );
and \U$49731 ( \50074 , \49987 , \50073 );
and \U$49732 ( \50075 , \49913 , \49986 );
or \U$49733 ( \50076 , \50074 , \50075 );
xor \U$49734 ( \50077 , \49830 , \50076 );
xor \U$49735 ( \50078 , \49192 , \49199 );
xor \U$49736 ( \50079 , \50078 , \49207 );
xor \U$49737 ( \50080 , \49393 , \49398 );
xor \U$49738 ( \50081 , \50079 , \50080 );
xor \U$49739 ( \50082 , \49347 , \49349 );
xor \U$49740 ( \50083 , \50082 , \49352 );
and \U$49741 ( \50084 , \50081 , \50083 );
xor \U$49742 ( \50085 , \49111 , \49118 );
xor \U$49743 ( \50086 , \50085 , \49126 );
xor \U$49744 ( \50087 , \49656 , \49661 );
xor \U$49745 ( \50088 , \50086 , \50087 );
xor \U$49746 ( \50089 , \49347 , \49349 );
xor \U$49747 ( \50090 , \50089 , \49352 );
and \U$49748 ( \50091 , \50088 , \50090 );
and \U$49749 ( \50092 , \50081 , \50088 );
or \U$49750 ( \50093 , \50084 , \50091 , \50092 );
and \U$49751 ( \50094 , \50077 , \50093 );
and \U$49752 ( \50095 , \49830 , \50076 );
or \U$49753 ( \50096 , \50094 , \50095 );
xor \U$49754 ( \50097 , \49767 , \50096 );
xor \U$49755 ( \50098 , \49487 , \49569 );
xor \U$49756 ( \50099 , \50098 , \49650 );
xor \U$49757 ( \50100 , \49666 , \49668 );
xor \U$49758 ( \50101 , \50100 , \49673 );
and \U$49759 ( \50102 , \50099 , \50101 );
xor \U$49760 ( \50103 , \49355 , \49390 );
xor \U$49761 ( \50104 , \50103 , \49403 );
xor \U$49762 ( \50105 , \49666 , \49668 );
xor \U$49763 ( \50106 , \50105 , \49673 );
and \U$49764 ( \50107 , \50104 , \50106 );
and \U$49765 ( \50108 , \50099 , \50104 );
or \U$49766 ( \50109 , \50102 , \50107 , \50108 );
and \U$49767 ( \50110 , \50097 , \50109 );
and \U$49768 ( \50111 , \49767 , \50096 );
or \U$49769 ( \50112 , \50110 , \50111 );
xor \U$49770 ( \50113 , \49059 , \49132 );
xor \U$49771 ( \50114 , \50113 , \49213 );
xor \U$49772 ( \50115 , \48906 , \48960 );
xor \U$49773 ( \50116 , \50115 , \48973 );
and \U$49774 ( \50117 , \50114 , \50116 );
xor \U$49775 ( \50118 , \49253 , \49255 );
xor \U$49776 ( \50119 , \50118 , \49258 );
xor \U$49777 ( \50120 , \49682 , \49689 );
xor \U$49778 ( \50121 , \50119 , \50120 );
xor \U$49779 ( \50122 , \48906 , \48960 );
xor \U$49780 ( \50123 , \50122 , \48973 );
and \U$49781 ( \50124 , \50121 , \50123 );
and \U$49782 ( \50125 , \50114 , \50121 );
or \U$49783 ( \50126 , \50117 , \50124 , \50125 );
xor \U$49784 ( \50127 , \50112 , \50126 );
xor \U$49785 ( \50128 , \48888 , \48890 );
xor \U$49786 ( \50129 , \50128 , \48893 );
xor \U$49787 ( \50130 , \49700 , \49705 );
xor \U$49788 ( \50131 , \50129 , \50130 );
and \U$49789 ( \50132 , \50127 , \50131 );
and \U$49790 ( \50133 , \50112 , \50126 );
or \U$49791 ( \50134 , \50132 , \50133 );
xor \U$49792 ( \50135 , \49743 , \50134 );
xor \U$49793 ( \50136 , \49313 , \49697 );
xor \U$49794 ( \50137 , \50136 , \49710 );
and \U$49795 ( \50138 , \50135 , \50137 );
and \U$49796 ( \50139 , \49743 , \50134 );
or \U$49797 ( \50140 , \50138 , \50139 );
not \U$49798 ( \50141 , \49300 );
not \U$49799 ( \50142 , \49303 );
or \U$49800 ( \50143 , \50141 , \50142 );
or \U$49801 ( \50144 , \49303 , \49300 );
nand \U$49802 ( \50145 , \50143 , \50144 );
xor \U$49803 ( \50146 , \50140 , \50145 );
not \U$49804 ( \50147 , \49716 );
xor \U$49805 ( \50148 , \49729 , \49713 );
not \U$49806 ( \50149 , \50148 );
or \U$49807 ( \50150 , \50147 , \50149 );
or \U$49808 ( \50151 , \50148 , \49716 );
nand \U$49809 ( \50152 , \50150 , \50151 );
and \U$49810 ( \50153 , \50146 , \50152 );
and \U$49811 ( \50154 , \50140 , \50145 );
or \U$49812 ( \50155 , \50153 , \50154 );
and \U$49813 ( \50156 , \49741 , \50155 );
xor \U$49814 ( \50157 , \50155 , \49741 );
xor \U$49815 ( \50158 , \49345 , \49679 );
xor \U$49816 ( \50159 , \50158 , \49694 );
xor \U$49817 ( \50160 , \48906 , \48960 );
xor \U$49818 ( \50161 , \50160 , \48973 );
xor \U$49819 ( \50162 , \50114 , \50121 );
xor \U$49820 ( \50163 , \50161 , \50162 );
xor \U$49821 ( \50164 , \49406 , \49653 );
xor \U$49822 ( \50165 , \50164 , \49676 );
xor \U$49823 ( \50166 , \50163 , \50165 );
xor \U$49824 ( \50167 , \49767 , \50096 );
xor \U$49825 ( \50168 , \50167 , \50109 );
and \U$49826 ( \50169 , \50166 , \50168 );
and \U$49827 ( \50170 , \50163 , \50165 );
or \U$49828 ( \50171 , \50169 , \50170 );
xor \U$49829 ( \50172 , \50159 , \50171 );
xor \U$49830 ( \50173 , \49913 , \49986 );
xor \U$49831 ( \50174 , \50173 , \50073 );
xor \U$49832 ( \50175 , \49779 , \49814 );
xor \U$49833 ( \50176 , \50175 , \49827 );
and \U$49834 ( \50177 , \50174 , \50176 );
xor \U$49835 ( \50178 , \49347 , \49349 );
xor \U$49836 ( \50179 , \50178 , \49352 );
xor \U$49837 ( \50180 , \50081 , \50088 );
xor \U$49838 ( \50181 , \50179 , \50180 );
xor \U$49839 ( \50182 , \49779 , \49814 );
xor \U$49840 ( \50183 , \50182 , \49827 );
and \U$49841 ( \50184 , \50181 , \50183 );
and \U$49842 ( \50185 , \50174 , \50181 );
or \U$49843 ( \50186 , \50177 , \50184 , \50185 );
and \U$49844 ( \50187 , \6453 , RI986eb48_32);
and \U$49845 ( \50188 , RI986ea58_30, \6451 );
nor \U$49846 ( \50189 , \50187 , \50188 );
and \U$49847 ( \50190 , \50189 , \6190 );
not \U$49848 ( \50191 , \50189 );
and \U$49849 ( \50192 , \50191 , \6705 );
nor \U$49850 ( \50193 , \50190 , \50192 );
and \U$49851 ( \50194 , \5318 , RI9871758_126);
and \U$49852 ( \50195 , RI9871848_128, \5316 );
nor \U$49853 ( \50196 , \50194 , \50195 );
and \U$49854 ( \50197 , \50196 , \5052 );
not \U$49855 ( \50198 , \50196 );
and \U$49856 ( \50199 , \50198 , \5322 );
nor \U$49857 ( \50200 , \50197 , \50199 );
xor \U$49858 ( \50201 , \50193 , \50200 );
and \U$49859 ( \50202 , \5881 , RI9871578_122);
and \U$49860 ( \50203 , RI9871668_124, \5879 );
nor \U$49861 ( \50204 , \50202 , \50203 );
and \U$49862 ( \50205 , \50204 , \5594 );
not \U$49863 ( \50206 , \50204 );
and \U$49864 ( \50207 , \50206 , \5885 );
nor \U$49865 ( \50208 , \50205 , \50207 );
and \U$49866 ( \50209 , \50201 , \50208 );
and \U$49867 ( \50210 , \50193 , \50200 );
or \U$49868 ( \50211 , \50209 , \50210 );
not \U$49869 ( \50212 , \50211 );
and \U$49870 ( \50213 , \7079 , RI986e968_28);
and \U$49871 ( \50214 , RI986e878_26, \7077 );
nor \U$49872 ( \50215 , \50213 , \50214 );
and \U$49873 ( \50216 , \50215 , \6709 );
not \U$49874 ( \50217 , \50215 );
and \U$49875 ( \50218 , \50217 , \6710 );
nor \U$49876 ( \50219 , \50216 , \50218 );
not \U$49877 ( \50220 , \50219 );
and \U$49878 ( \50221 , \7729 , RI986ef08_40);
and \U$49879 ( \50222 , RI986ee18_38, \7727 );
nor \U$49880 ( \50223 , \50221 , \50222 );
and \U$49881 ( \50224 , \50223 , \7733 );
not \U$49882 ( \50225 , \50223 );
and \U$49883 ( \50226 , \50225 , \7480 );
nor \U$49884 ( \50227 , \50224 , \50226 );
not \U$49885 ( \50228 , \50227 );
and \U$49886 ( \50229 , \50220 , \50228 );
and \U$49887 ( \50230 , \50227 , \50219 );
and \U$49888 ( \50231 , \8486 , RI986ec38_34);
and \U$49889 ( \50232 , RI986ed28_36, \8484 );
nor \U$49890 ( \50233 , \50231 , \50232 );
and \U$49891 ( \50234 , \50233 , \8051 );
not \U$49892 ( \50235 , \50233 );
and \U$49893 ( \50236 , \50235 , \8050 );
nor \U$49894 ( \50237 , \50234 , \50236 );
nor \U$49895 ( \50238 , \50230 , \50237 );
nor \U$49896 ( \50239 , \50229 , \50238 );
or \U$49897 ( \50240 , \50212 , \50239 );
and \U$49898 ( \50241 , \50212 , \50239 );
and \U$49899 ( \50242 , \4203 , RI98712a8_116);
and \U$49900 ( \50243 , RI98711b8_114, \4201 );
nor \U$49901 ( \50244 , \50242 , \50243 );
and \U$49902 ( \50245 , \50244 , \4207 );
not \U$49903 ( \50246 , \50244 );
and \U$49904 ( \50247 , \50246 , \3923 );
nor \U$49905 ( \50248 , \50245 , \50247 );
not \U$49906 ( \50249 , \4519 );
and \U$49907 ( \50250 , \4710 , RI9871398_118);
and \U$49908 ( \50251 , RI9871488_120, \4708 );
nor \U$49909 ( \50252 , \50250 , \50251 );
not \U$49910 ( \50253 , \50252 );
or \U$49911 ( \50254 , \50249 , \50253 );
or \U$49912 ( \50255 , \50252 , \4521 );
nand \U$49913 ( \50256 , \50254 , \50255 );
xor \U$49914 ( \50257 , \50248 , \50256 );
not \U$49915 ( \50258 , \3918 );
and \U$49916 ( \50259 , \3683 , RI98710c8_112);
and \U$49917 ( \50260 , RI9870d08_104, \3681 );
nor \U$49918 ( \50261 , \50259 , \50260 );
not \U$49919 ( \50262 , \50261 );
or \U$49920 ( \50263 , \50258 , \50262 );
or \U$49921 ( \50264 , \50261 , \3412 );
nand \U$49922 ( \50265 , \50263 , \50264 );
and \U$49923 ( \50266 , \50257 , \50265 );
and \U$49924 ( \50267 , \50248 , \50256 );
nor \U$49925 ( \50268 , \50266 , \50267 );
nor \U$49926 ( \50269 , \50241 , \50268 );
not \U$49927 ( \50270 , \50269 );
nand \U$49928 ( \50271 , \50240 , \50270 );
and \U$49929 ( \50272 , \776 , RI9870948_96);
and \U$49930 ( \50273 , RI9870858_94, \774 );
nor \U$49931 ( \50274 , \50272 , \50273 );
and \U$49932 ( \50275 , \50274 , \451 );
not \U$49933 ( \50276 , \50274 );
and \U$49934 ( \50277 , \50276 , \474 );
nor \U$49935 ( \50278 , \50275 , \50277 );
not \U$49936 ( \50279 , \50278 );
and \U$49937 ( \50280 , \438 , RI9870768_92);
and \U$49938 ( \50281 , RI9870678_90, \436 );
nor \U$49939 ( \50282 , \50280 , \50281 );
and \U$49940 ( \50283 , \50282 , \443 );
not \U$49941 ( \50284 , \50282 );
and \U$49942 ( \50285 , \50284 , \444 );
nor \U$49943 ( \50286 , \50283 , \50285 );
not \U$49944 ( \50287 , \50286 );
and \U$49945 ( \50288 , \50279 , \50287 );
and \U$49946 ( \50289 , \50286 , \50278 );
and \U$49947 ( \50290 , \1293 , RI986fb38_66);
and \U$49948 ( \50291 , RI986fc28_68, \1291 );
nor \U$49949 ( \50292 , \50290 , \50291 );
not \U$49950 ( \50293 , \50292 );
not \U$49951 ( \50294 , \1301 );
and \U$49952 ( \50295 , \50293 , \50294 );
and \U$49953 ( \50296 , \50292 , \1128 );
nor \U$49954 ( \50297 , \50295 , \50296 );
nor \U$49955 ( \50298 , \50289 , \50297 );
nor \U$49956 ( \50299 , \50288 , \50298 );
and \U$49957 ( \50300 , \2464 , RI9870df8_106);
and \U$49958 ( \50301 , RI9870a38_98, \2462 );
nor \U$49959 ( \50302 , \50300 , \50301 );
and \U$49960 ( \50303 , \50302 , \2468 );
not \U$49961 ( \50304 , \50302 );
and \U$49962 ( \50305 , \50304 , \2263 );
nor \U$49963 ( \50306 , \50303 , \50305 );
not \U$49964 ( \50307 , \2935 );
and \U$49965 ( \50308 , \3254 , RI9870ee8_108);
and \U$49966 ( \50309 , RI9870c18_102, \3252 );
nor \U$49967 ( \50310 , \50308 , \50309 );
not \U$49968 ( \50311 , \50310 );
or \U$49969 ( \50312 , \50307 , \50311 );
or \U$49970 ( \50313 , \50310 , \2935 );
nand \U$49971 ( \50314 , \50312 , \50313 );
xor \U$49972 ( \50315 , \50306 , \50314 );
and \U$49973 ( \50316 , \2274 , RI9870fd8_110);
and \U$49974 ( \50317 , RI9870b28_100, \2272 );
nor \U$49975 ( \50318 , \50316 , \50317 );
and \U$49976 ( \50319 , \50318 , \2030 );
not \U$49977 ( \50320 , \50318 );
and \U$49978 ( \50321 , \50320 , \2031 );
nor \U$49979 ( \50322 , \50319 , \50321 );
and \U$49980 ( \50323 , \50315 , \50322 );
and \U$49981 ( \50324 , \50306 , \50314 );
nor \U$49982 ( \50325 , \50323 , \50324 );
or \U$49983 ( \50326 , \50299 , \50325 );
not \U$49984 ( \50327 , \50299 );
not \U$49985 ( \50328 , \50325 );
or \U$49986 ( \50329 , \50327 , \50328 );
and \U$49987 ( \50330 , \1329 , RI986fe08_72);
and \U$49988 ( \50331 , RI986fd18_70, \1327 );
nor \U$49989 ( \50332 , \50330 , \50331 );
and \U$49990 ( \50333 , \50332 , \1336 );
not \U$49991 ( \50334 , \50332 );
and \U$49992 ( \50335 , \50334 , \1337 );
nor \U$49993 ( \50336 , \50333 , \50335 );
and \U$49994 ( \50337 , \1311 , RI986ffe8_76);
and \U$49995 ( \50338 , RI986fef8_74, \1309 );
nor \U$49996 ( \50339 , \50337 , \50338 );
and \U$49997 ( \50340 , \50339 , \1458 );
not \U$49998 ( \50341 , \50339 );
and \U$49999 ( \50342 , \50341 , \1315 );
nor \U$50000 ( \50343 , \50340 , \50342 );
xor \U$50001 ( \50344 , \50336 , \50343 );
not \U$50002 ( \50345 , \1462 );
and \U$50003 ( \50346 , \2042 , RI98700d8_78);
and \U$50004 ( \50347 , RI98701c8_80, \2040 );
nor \U$50005 ( \50348 , \50346 , \50347 );
not \U$50006 ( \50349 , \50348 );
or \U$50007 ( \50350 , \50345 , \50349 );
or \U$50008 ( \50351 , \50348 , \1462 );
nand \U$50009 ( \50352 , \50350 , \50351 );
and \U$50010 ( \50353 , \50344 , \50352 );
and \U$50011 ( \50354 , \50336 , \50343 );
or \U$50012 ( \50355 , \50353 , \50354 );
nand \U$50013 ( \50356 , \50329 , \50355 );
nand \U$50014 ( \50357 , \50326 , \50356 );
xor \U$50015 ( \50358 , \50271 , \50357 );
and \U$50016 ( \50359 , \9505 , RI986f2c8_48);
and \U$50017 ( \50360 , RI986f1d8_46, \9503 );
nor \U$50018 ( \50361 , \50359 , \50360 );
and \U$50019 ( \50362 , \50361 , \9510 );
not \U$50020 ( \50363 , \50361 );
and \U$50021 ( \50364 , \50363 , \9513 );
nor \U$50022 ( \50365 , \50362 , \50364 );
and \U$50023 ( \50366 , \10424 , RI986e5a8_20);
and \U$50024 ( \50367 , RI986e4b8_18, \10422 );
nor \U$50025 ( \50368 , \50366 , \50367 );
and \U$50026 ( \50369 , \50368 , \9840 );
not \U$50027 ( \50370 , \50368 );
and \U$50028 ( \50371 , \50370 , \10428 );
nor \U$50029 ( \50372 , \50369 , \50371 );
xor \U$50030 ( \50373 , \50365 , \50372 );
and \U$50031 ( \50374 , \9237 , RI986f0e8_44);
and \U$50032 ( \50375 , RI986eff8_42, \9235 );
nor \U$50033 ( \50376 , \50374 , \50375 );
and \U$50034 ( \50377 , \50376 , \9241 );
not \U$50035 ( \50378 , \50376 );
and \U$50036 ( \50379 , \50378 , \8836 );
nor \U$50037 ( \50380 , \50377 , \50379 );
and \U$50038 ( \50381 , \50373 , \50380 );
and \U$50039 ( \50382 , \50365 , \50372 );
nor \U$50040 ( \50383 , \50381 , \50382 );
and \U$50041 ( \50384 , \11696 , RI986e788_24);
and \U$50042 ( \50385 , RI986e698_22, \11694 );
nor \U$50043 ( \50386 , \50384 , \50385 );
and \U$50044 ( \50387 , \50386 , \11702 );
not \U$50045 ( \50388 , \50386 );
and \U$50046 ( \50389 , \50388 , \10965 );
nor \U$50047 ( \50390 , \50387 , \50389 );
not \U$50048 ( \50391 , \50390 );
and \U$50049 ( \50392 , \13045 , RI986fa48_64);
and \U$50050 ( \50393 , RI986f958_62, \13043 );
nor \U$50051 ( \50394 , \50392 , \50393 );
and \U$50052 ( \50395 , \50394 , \12619 );
not \U$50053 ( \50396 , \50394 );
and \U$50054 ( \50397 , \50396 , \13047 );
nor \U$50055 ( \50398 , \50395 , \50397 );
not \U$50056 ( \50399 , \50398 );
and \U$50057 ( \50400 , \50391 , \50399 );
and \U$50058 ( \50401 , \50398 , \50390 );
and \U$50059 ( \50402 , \12293 , RI986f868_60);
and \U$50060 ( \50403 , RI986f778_58, \12291 );
nor \U$50061 ( \50404 , \50402 , \50403 );
and \U$50062 ( \50405 , \50404 , \11686 );
not \U$50063 ( \50406 , \50404 );
and \U$50064 ( \50407 , \50406 , \11687 );
nor \U$50065 ( \50408 , \50405 , \50407 );
nor \U$50066 ( \50409 , \50401 , \50408 );
nor \U$50067 ( \50410 , \50400 , \50409 );
or \U$50068 ( \50411 , \50383 , \50410 );
not \U$50069 ( \50412 , \50383 );
not \U$50070 ( \50413 , \50410 );
or \U$50071 ( \50414 , \50412 , \50413 );
and \U$50072 ( \50415 , \14937 , RI986f598_54);
and \U$50073 ( \50416 , RI986f688_56, \14935 );
nor \U$50074 ( \50417 , \50415 , \50416 );
and \U$50075 ( \50418 , \50417 , \14539 );
not \U$50076 ( \50419 , \50417 );
and \U$50077 ( \50420 , \50419 , \14538 );
nor \U$50078 ( \50421 , \50418 , \50420 );
not \U$50079 ( \50422 , RI9873558_190);
and \U$50080 ( \50423 , \15780 , RI986e008_8);
and \U$50081 ( \50424 , RI986df18_6, RI9873648_192);
nor \U$50082 ( \50425 , \50423 , \50424 );
not \U$50083 ( \50426 , \50425 );
or \U$50084 ( \50427 , \50422 , \50426 );
or \U$50085 ( \50428 , \50425 , RI9873558_190);
nand \U$50086 ( \50429 , \50427 , \50428 );
xor \U$50087 ( \50430 , \50421 , \50429 );
and \U$50088 ( \50431 , \13882 , RI986f4a8_52);
and \U$50089 ( \50432 , RI986f3b8_50, \13880 );
nor \U$50090 ( \50433 , \50431 , \50432 );
and \U$50091 ( \50434 , \50433 , \13358 );
not \U$50092 ( \50435 , \50433 );
and \U$50093 ( \50436 , \50435 , \13359 );
nor \U$50094 ( \50437 , \50434 , \50436 );
and \U$50095 ( \50438 , \50430 , \50437 );
and \U$50096 ( \50439 , \50421 , \50429 );
or \U$50097 ( \50440 , \50438 , \50439 );
nand \U$50098 ( \50441 , \50414 , \50440 );
nand \U$50099 ( \50442 , \50411 , \50441 );
and \U$50100 ( \50443 , \50358 , \50442 );
and \U$50101 ( \50444 , \50271 , \50357 );
or \U$50102 ( \50445 , \50443 , \50444 );
xor \U$50103 ( \50446 , \49629 , \49636 );
xor \U$50104 ( \50447 , \50446 , \49644 );
xor \U$50105 ( \50448 , \49602 , \49610 );
xor \U$50106 ( \50449 , \50448 , \49618 );
xor \U$50107 ( \50450 , \50447 , \50449 );
xor \U$50108 ( \50451 , \49413 , \49420 );
xor \U$50109 ( \50452 , \50451 , \49428 );
xor \U$50110 ( \50453 , \49769 , \49774 );
xor \U$50111 ( \50454 , \50452 , \50453 );
and \U$50112 ( \50455 , \50450 , \50454 );
and \U$50113 ( \50456 , \50447 , \50449 );
or \U$50114 ( \50457 , \50455 , \50456 );
xor \U$50115 ( \50458 , \50445 , \50457 );
xor \U$50116 ( \50459 , \49892 , \49899 );
xor \U$50117 ( \50460 , \50459 , \49907 );
xor \U$50118 ( \50461 , \49838 , \49845 );
xor \U$50119 ( \50462 , \50461 , \49854 );
and \U$50120 ( \50463 , \50460 , \50462 );
not \U$50121 ( \50464 , \49994 );
xor \U$50122 ( \50465 , \50003 , \50013 );
not \U$50123 ( \50466 , \50465 );
or \U$50124 ( \50467 , \50464 , \50466 );
or \U$50125 ( \50468 , \50465 , \49994 );
nand \U$50126 ( \50469 , \50467 , \50468 );
xor \U$50127 ( \50470 , \49838 , \49845 );
xor \U$50128 ( \50471 , \50470 , \49854 );
and \U$50129 ( \50472 , \50469 , \50471 );
and \U$50130 ( \50473 , \50460 , \50469 );
or \U$50131 ( \50474 , \50463 , \50472 , \50473 );
nand \U$50132 ( \50475 , RI9870498_86, \393 );
not \U$50133 ( \50476 , \50475 );
not \U$50134 ( \50477 , \386 );
or \U$50135 ( \50478 , \50476 , \50477 );
or \U$50136 ( \50479 , \386 , \50475 );
nand \U$50137 ( \50480 , \50478 , \50479 );
xor \U$50138 ( \50481 , \49864 , \49871 );
xor \U$50139 ( \50482 , \50481 , \49880 );
and \U$50140 ( \50483 , \50480 , \50482 );
xor \U$50141 ( \50484 , \49789 , \49796 );
xor \U$50142 ( \50485 , \50484 , \49805 );
xor \U$50143 ( \50486 , \49864 , \49871 );
xor \U$50144 ( \50487 , \50486 , \49880 );
and \U$50145 ( \50488 , \50485 , \50487 );
and \U$50146 ( \50489 , \50480 , \50485 );
or \U$50147 ( \50490 , \50483 , \50488 , \50489 );
xor \U$50148 ( \50491 , \50474 , \50490 );
not \U$50149 ( \50492 , \50022 );
xor \U$50150 ( \50493 , \50030 , \50040 );
not \U$50151 ( \50494 , \50493 );
or \U$50152 ( \50495 , \50492 , \50494 );
or \U$50153 ( \50496 , \50493 , \50022 );
nand \U$50154 ( \50497 , \50495 , \50496 );
xor \U$50155 ( \50498 , \50053 , \50060 );
xor \U$50156 ( \50499 , \50498 , \50068 );
xor \U$50157 ( \50500 , \50497 , \50499 );
xor \U$50158 ( \50501 , \49920 , \49927 );
xor \U$50159 ( \50502 , \50501 , \49935 );
and \U$50160 ( \50503 , \50500 , \50502 );
and \U$50161 ( \50504 , \50497 , \50499 );
or \U$50162 ( \50505 , \50503 , \50504 );
and \U$50163 ( \50506 , \50491 , \50505 );
and \U$50164 ( \50507 , \50474 , \50490 );
or \U$50165 ( \50508 , \50506 , \50507 );
and \U$50166 ( \50509 , \50458 , \50508 );
and \U$50167 ( \50510 , \50445 , \50457 );
or \U$50168 ( \50511 , \50509 , \50510 );
xor \U$50169 ( \50512 , \50186 , \50511 );
xor \U$50170 ( \50513 , \49857 , \49883 );
xor \U$50171 ( \50514 , \50513 , \49910 );
xor \U$50172 ( \50515 , \49781 , \49808 );
xor \U$50173 ( \50516 , \50515 , \49811 );
and \U$50174 ( \50517 , \50514 , \50516 );
xor \U$50175 ( \50518 , \49494 , \49501 );
xor \U$50176 ( \50519 , \50518 , \49510 );
xor \U$50177 ( \50520 , \49817 , \49822 );
xor \U$50178 ( \50521 , \50519 , \50520 );
xor \U$50179 ( \50522 , \49781 , \49808 );
xor \U$50180 ( \50523 , \50522 , \49811 );
and \U$50181 ( \50524 , \50521 , \50523 );
and \U$50182 ( \50525 , \50514 , \50521 );
or \U$50183 ( \50526 , \50517 , \50524 , \50525 );
xor \U$50184 ( \50527 , \49595 , \49621 );
xor \U$50185 ( \50528 , \50527 , \49647 );
xor \U$50186 ( \50529 , \50526 , \50528 );
xor \U$50187 ( \50530 , \49431 , \49458 );
xor \U$50188 ( \50531 , \50530 , \49484 );
xor \U$50189 ( \50532 , \49749 , \49754 );
xor \U$50190 ( \50533 , \50531 , \50532 );
and \U$50191 ( \50534 , \50529 , \50533 );
and \U$50192 ( \50535 , \50526 , \50528 );
or \U$50193 ( \50536 , \50534 , \50535 );
and \U$50194 ( \50537 , \50512 , \50536 );
and \U$50195 ( \50538 , \50186 , \50511 );
or \U$50196 ( \50539 , \50537 , \50538 );
xor \U$50197 ( \50540 , \49325 , \49327 );
xor \U$50198 ( \50541 , \50540 , \49342 );
xor \U$50199 ( \50542 , \50539 , \50541 );
xor \U$50200 ( \50543 , \49830 , \50076 );
xor \U$50201 ( \50544 , \50543 , \50093 );
xor \U$50202 ( \50545 , \49747 , \49759 );
xor \U$50203 ( \50546 , \50545 , \49764 );
and \U$50204 ( \50547 , \50544 , \50546 );
xor \U$50205 ( \50548 , \49666 , \49668 );
xor \U$50206 ( \50549 , \50548 , \49673 );
xor \U$50207 ( \50550 , \50099 , \50104 );
xor \U$50208 ( \50551 , \50549 , \50550 );
xor \U$50209 ( \50552 , \49747 , \49759 );
xor \U$50210 ( \50553 , \50552 , \49764 );
and \U$50211 ( \50554 , \50551 , \50553 );
and \U$50212 ( \50555 , \50544 , \50551 );
or \U$50213 ( \50556 , \50547 , \50554 , \50555 );
and \U$50214 ( \50557 , \50542 , \50556 );
and \U$50215 ( \50558 , \50539 , \50541 );
or \U$50216 ( \50559 , \50557 , \50558 );
and \U$50217 ( \50560 , \50172 , \50559 );
and \U$50218 ( \50561 , \50159 , \50171 );
nor \U$50219 ( \50562 , \50560 , \50561 );
not \U$50220 ( \50563 , \50562 );
xor \U$50221 ( \50564 , \49743 , \50134 );
xor \U$50222 ( \50565 , \50564 , \50137 );
not \U$50223 ( \50566 , \50565 );
or \U$50224 ( \50567 , \50563 , \50566 );
or \U$50225 ( \50568 , \50565 , \50562 );
nand \U$50226 ( \50569 , \50567 , \50568 );
xor \U$50227 ( \50570 , \50445 , \50457 );
xor \U$50228 ( \50571 , \50570 , \50508 );
xor \U$50229 ( \50572 , \50526 , \50528 );
xor \U$50230 ( \50573 , \50572 , \50533 );
and \U$50231 ( \50574 , \50571 , \50573 );
xor \U$50232 ( \50575 , \49779 , \49814 );
xor \U$50233 ( \50576 , \50575 , \49827 );
xor \U$50234 ( \50577 , \50174 , \50181 );
xor \U$50235 ( \50578 , \50576 , \50577 );
xor \U$50236 ( \50579 , \50526 , \50528 );
xor \U$50237 ( \50580 , \50579 , \50533 );
and \U$50238 ( \50581 , \50578 , \50580 );
and \U$50239 ( \50582 , \50571 , \50578 );
or \U$50240 ( \50583 , \50574 , \50581 , \50582 );
xor \U$50241 ( \50584 , \49938 , \49957 );
xor \U$50242 ( \50585 , \50584 , \49983 );
xor \U$50243 ( \50586 , \50447 , \50449 );
xor \U$50244 ( \50587 , \50586 , \50454 );
and \U$50245 ( \50588 , \50585 , \50587 );
xor \U$50246 ( \50589 , \49781 , \49808 );
xor \U$50247 ( \50590 , \50589 , \49811 );
xor \U$50248 ( \50591 , \50514 , \50521 );
xor \U$50249 ( \50592 , \50590 , \50591 );
xor \U$50250 ( \50593 , \50447 , \50449 );
xor \U$50251 ( \50594 , \50593 , \50454 );
and \U$50252 ( \50595 , \50592 , \50594 );
and \U$50253 ( \50596 , \50585 , \50592 );
or \U$50254 ( \50597 , \50588 , \50595 , \50596 );
not \U$50255 ( \50598 , \50597 );
not \U$50256 ( \50599 , \50440 );
not \U$50257 ( \50600 , \50410 );
or \U$50258 ( \50601 , \50599 , \50600 );
or \U$50259 ( \50602 , \50410 , \50440 );
nand \U$50260 ( \50603 , \50601 , \50602 );
not \U$50261 ( \50604 , \50603 );
not \U$50262 ( \50605 , \50383 );
and \U$50263 ( \50606 , \50604 , \50605 );
and \U$50264 ( \50607 , \50603 , \50383 );
nor \U$50265 ( \50608 , \50606 , \50607 );
not \U$50266 ( \50609 , \50608 );
not \U$50267 ( \50610 , \50355 );
not \U$50268 ( \50611 , \50299 );
or \U$50269 ( \50612 , \50610 , \50611 );
or \U$50270 ( \50613 , \50299 , \50355 );
nand \U$50271 ( \50614 , \50612 , \50613 );
not \U$50272 ( \50615 , \50614 );
not \U$50273 ( \50616 , \50325 );
and \U$50274 ( \50617 , \50615 , \50616 );
and \U$50275 ( \50618 , \50614 , \50325 );
nor \U$50276 ( \50619 , \50617 , \50618 );
not \U$50277 ( \50620 , \50619 );
and \U$50278 ( \50621 , \50609 , \50620 );
and \U$50279 ( \50622 , \50608 , \50619 );
not \U$50280 ( \50623 , \50211 );
not \U$50281 ( \50624 , \50268 );
or \U$50282 ( \50625 , \50623 , \50624 );
or \U$50283 ( \50626 , \50268 , \50211 );
nand \U$50284 ( \50627 , \50625 , \50626 );
not \U$50285 ( \50628 , \50627 );
not \U$50286 ( \50629 , \50239 );
and \U$50287 ( \50630 , \50628 , \50629 );
and \U$50288 ( \50631 , \50627 , \50239 );
nor \U$50289 ( \50632 , \50630 , \50631 );
nor \U$50290 ( \50633 , \50622 , \50632 );
nor \U$50291 ( \50634 , \50621 , \50633 );
not \U$50292 ( \50635 , \50071 );
not \U$50293 ( \50636 , \50015 );
or \U$50294 ( \50637 , \50635 , \50636 );
or \U$50295 ( \50638 , \50015 , \50071 );
nand \U$50296 ( \50639 , \50637 , \50638 );
not \U$50297 ( \50640 , \50639 );
not \U$50298 ( \50641 , \50042 );
and \U$50299 ( \50642 , \50640 , \50641 );
and \U$50300 ( \50643 , \50639 , \50042 );
nor \U$50301 ( \50644 , \50642 , \50643 );
or \U$50302 ( \50645 , \50634 , \50644 );
not \U$50303 ( \50646 , \50644 );
not \U$50304 ( \50647 , \50634 );
or \U$50305 ( \50648 , \50646 , \50647 );
xor \U$50306 ( \50649 , \49864 , \49871 );
xor \U$50307 ( \50650 , \50649 , \49880 );
xor \U$50308 ( \50651 , \50480 , \50485 );
xor \U$50309 ( \50652 , \50650 , \50651 );
xor \U$50310 ( \50653 , \50497 , \50499 );
xor \U$50311 ( \50654 , \50653 , \50502 );
and \U$50312 ( \50655 , \50652 , \50654 );
xor \U$50313 ( \50656 , \49838 , \49845 );
xor \U$50314 ( \50657 , \50656 , \49854 );
xor \U$50315 ( \50658 , \50460 , \50469 );
xor \U$50316 ( \50659 , \50657 , \50658 );
xor \U$50317 ( \50660 , \50497 , \50499 );
xor \U$50318 ( \50661 , \50660 , \50502 );
and \U$50319 ( \50662 , \50659 , \50661 );
and \U$50320 ( \50663 , \50652 , \50659 );
or \U$50321 ( \50664 , \50655 , \50662 , \50663 );
nand \U$50322 ( \50665 , \50648 , \50664 );
nand \U$50323 ( \50666 , \50645 , \50665 );
not \U$50324 ( \50667 , \50666 );
or \U$50325 ( \50668 , \50598 , \50667 );
or \U$50326 ( \50669 , \50666 , \50597 );
and \U$50327 ( \50670 , \8486 , RI986ee18_38);
and \U$50328 ( \50671 , RI986ec38_34, \8484 );
nor \U$50329 ( \50672 , \50670 , \50671 );
and \U$50330 ( \50673 , \50672 , \8050 );
not \U$50331 ( \50674 , \50672 );
and \U$50332 ( \50675 , \50674 , \8051 );
nor \U$50333 ( \50676 , \50673 , \50675 );
and \U$50334 ( \50677 , \7729 , RI986e878_26);
and \U$50335 ( \50678 , RI986ef08_40, \7727 );
nor \U$50336 ( \50679 , \50677 , \50678 );
and \U$50337 ( \50680 , \50679 , \7480 );
not \U$50338 ( \50681 , \50679 );
and \U$50339 ( \50682 , \50681 , \7733 );
nor \U$50340 ( \50683 , \50680 , \50682 );
xor \U$50341 ( \50684 , \50676 , \50683 );
and \U$50342 ( \50685 , \9237 , RI986ed28_36);
and \U$50343 ( \50686 , RI986f0e8_44, \9235 );
nor \U$50344 ( \50687 , \50685 , \50686 );
and \U$50345 ( \50688 , \50687 , \9241 );
not \U$50346 ( \50689 , \50687 );
and \U$50347 ( \50690 , \50689 , \8836 );
nor \U$50348 ( \50691 , \50688 , \50690 );
and \U$50349 ( \50692 , \50684 , \50691 );
and \U$50350 ( \50693 , \50676 , \50683 );
or \U$50351 ( \50694 , \50692 , \50693 );
and \U$50352 ( \50695 , \5318 , RI9871488_120);
and \U$50353 ( \50696 , RI9871758_126, \5316 );
nor \U$50354 ( \50697 , \50695 , \50696 );
and \U$50355 ( \50698 , \50697 , \5052 );
not \U$50356 ( \50699 , \50697 );
and \U$50357 ( \50700 , \50699 , \5322 );
nor \U$50358 ( \50701 , \50698 , \50700 );
and \U$50359 ( \50702 , \4203 , RI9870d08_104);
and \U$50360 ( \50703 , RI98712a8_116, \4201 );
nor \U$50361 ( \50704 , \50702 , \50703 );
and \U$50362 ( \50705 , \50704 , \4207 );
not \U$50363 ( \50706 , \50704 );
and \U$50364 ( \50707 , \50706 , \3922 );
nor \U$50365 ( \50708 , \50705 , \50707 );
xor \U$50366 ( \50709 , \50701 , \50708 );
not \U$50367 ( \50710 , \4519 );
and \U$50368 ( \50711 , \4710 , RI98711b8_114);
and \U$50369 ( \50712 , RI9871398_118, \4708 );
nor \U$50370 ( \50713 , \50711 , \50712 );
not \U$50371 ( \50714 , \50713 );
or \U$50372 ( \50715 , \50710 , \50714 );
or \U$50373 ( \50716 , \50713 , \4519 );
nand \U$50374 ( \50717 , \50715 , \50716 );
and \U$50375 ( \50718 , \50709 , \50717 );
and \U$50376 ( \50719 , \50701 , \50708 );
or \U$50377 ( \50720 , \50718 , \50719 );
xor \U$50378 ( \50721 , \50694 , \50720 );
and \U$50379 ( \50722 , \7079 , RI986ea58_30);
and \U$50380 ( \50723 , RI986e968_28, \7077 );
nor \U$50381 ( \50724 , \50722 , \50723 );
and \U$50382 ( \50725 , \50724 , \6710 );
not \U$50383 ( \50726 , \50724 );
and \U$50384 ( \50727 , \50726 , \6709 );
nor \U$50385 ( \50728 , \50725 , \50727 );
and \U$50386 ( \50729 , \5881 , RI9871848_128);
and \U$50387 ( \50730 , RI9871578_122, \5879 );
nor \U$50388 ( \50731 , \50729 , \50730 );
and \U$50389 ( \50732 , \50731 , \5594 );
not \U$50390 ( \50733 , \50731 );
and \U$50391 ( \50734 , \50733 , \5885 );
nor \U$50392 ( \50735 , \50732 , \50734 );
xor \U$50393 ( \50736 , \50728 , \50735 );
and \U$50394 ( \50737 , \6453 , RI9871668_124);
and \U$50395 ( \50738 , RI986eb48_32, \6451 );
nor \U$50396 ( \50739 , \50737 , \50738 );
and \U$50397 ( \50740 , \50739 , \6190 );
not \U$50398 ( \50741 , \50739 );
and \U$50399 ( \50742 , \50741 , \6705 );
nor \U$50400 ( \50743 , \50740 , \50742 );
and \U$50401 ( \50744 , \50736 , \50743 );
and \U$50402 ( \50745 , \50728 , \50735 );
or \U$50403 ( \50746 , \50744 , \50745 );
and \U$50404 ( \50747 , \50721 , \50746 );
and \U$50405 ( \50748 , \50694 , \50720 );
or \U$50406 ( \50749 , \50747 , \50748 );
and \U$50407 ( \50750 , \13045 , RI986f778_58);
and \U$50408 ( \50751 , RI986fa48_64, \13043 );
nor \U$50409 ( \50752 , \50750 , \50751 );
and \U$50410 ( \50753 , \50752 , \13047 );
not \U$50411 ( \50754 , \50752 );
and \U$50412 ( \50755 , \50754 , \12619 );
nor \U$50413 ( \50756 , \50753 , \50755 );
and \U$50414 ( \50757 , \12293 , RI986e698_22);
and \U$50415 ( \50758 , RI986f868_60, \12291 );
nor \U$50416 ( \50759 , \50757 , \50758 );
and \U$50417 ( \50760 , \50759 , \11687 );
not \U$50418 ( \50761 , \50759 );
and \U$50419 ( \50762 , \50761 , \11686 );
nor \U$50420 ( \50763 , \50760 , \50762 );
xor \U$50421 ( \50764 , \50756 , \50763 );
and \U$50422 ( \50765 , \13882 , RI986f958_62);
and \U$50423 ( \50766 , RI986f4a8_52, \13880 );
nor \U$50424 ( \50767 , \50765 , \50766 );
and \U$50425 ( \50768 , \50767 , \13358 );
not \U$50426 ( \50769 , \50767 );
and \U$50427 ( \50770 , \50769 , \13359 );
nor \U$50428 ( \50771 , \50768 , \50770 );
and \U$50429 ( \50772 , \50764 , \50771 );
and \U$50430 ( \50773 , \50756 , \50763 );
or \U$50431 ( \50774 , \50772 , \50773 );
not \U$50432 ( \50775 , RI9873558_190);
and \U$50433 ( \50776 , \15780 , RI986f688_56);
and \U$50434 ( \50777 , RI986e008_8, RI9873648_192);
nor \U$50435 ( \50778 , \50776 , \50777 );
not \U$50436 ( \50779 , \50778 );
or \U$50437 ( \50780 , \50775 , \50779 );
or \U$50438 ( \50781 , \50778 , RI9873558_190);
nand \U$50439 ( \50782 , \50780 , \50781 );
xor \U$50440 ( \50783 , \50782 , \367 );
and \U$50441 ( \50784 , \14937 , RI986f3b8_50);
and \U$50442 ( \50785 , RI986f598_54, \14935 );
nor \U$50443 ( \50786 , \50784 , \50785 );
and \U$50444 ( \50787 , \50786 , \14539 );
not \U$50445 ( \50788 , \50786 );
and \U$50446 ( \50789 , \50788 , \14538 );
nor \U$50447 ( \50790 , \50787 , \50789 );
and \U$50448 ( \50791 , \50783 , \50790 );
and \U$50449 ( \50792 , \50782 , \367 );
or \U$50450 ( \50793 , \50791 , \50792 );
xor \U$50451 ( \50794 , \50774 , \50793 );
and \U$50452 ( \50795 , \9505 , RI986eff8_42);
and \U$50453 ( \50796 , RI986f2c8_48, \9503 );
nor \U$50454 ( \50797 , \50795 , \50796 );
and \U$50455 ( \50798 , \50797 , \9510 );
not \U$50456 ( \50799 , \50797 );
and \U$50457 ( \50800 , \50799 , \9513 );
nor \U$50458 ( \50801 , \50798 , \50800 );
and \U$50459 ( \50802 , \10424 , RI986f1d8_46);
and \U$50460 ( \50803 , RI986e5a8_20, \10422 );
nor \U$50461 ( \50804 , \50802 , \50803 );
and \U$50462 ( \50805 , \50804 , \9840 );
not \U$50463 ( \50806 , \50804 );
and \U$50464 ( \50807 , \50806 , \10428 );
nor \U$50465 ( \50808 , \50805 , \50807 );
xor \U$50466 ( \50809 , \50801 , \50808 );
and \U$50467 ( \50810 , \11696 , RI986e4b8_18);
and \U$50468 ( \50811 , RI986e788_24, \11694 );
nor \U$50469 ( \50812 , \50810 , \50811 );
and \U$50470 ( \50813 , \50812 , \10965 );
not \U$50471 ( \50814 , \50812 );
and \U$50472 ( \50815 , \50814 , \11702 );
nor \U$50473 ( \50816 , \50813 , \50815 );
and \U$50474 ( \50817 , \50809 , \50816 );
and \U$50475 ( \50818 , \50801 , \50808 );
or \U$50476 ( \50819 , \50817 , \50818 );
and \U$50477 ( \50820 , \50794 , \50819 );
and \U$50478 ( \50821 , \50774 , \50793 );
or \U$50479 ( \50822 , \50820 , \50821 );
xor \U$50480 ( \50823 , \50749 , \50822 );
not \U$50481 ( \50824 , \3406 );
and \U$50482 ( \50825 , \3254 , RI9870a38_98);
and \U$50483 ( \50826 , RI9870ee8_108, \3252 );
nor \U$50484 ( \50827 , \50825 , \50826 );
not \U$50485 ( \50828 , \50827 );
or \U$50486 ( \50829 , \50824 , \50828 );
or \U$50487 ( \50830 , \50827 , \3406 );
nand \U$50488 ( \50831 , \50829 , \50830 );
and \U$50489 ( \50832 , \2464 , RI9870b28_100);
and \U$50490 ( \50833 , RI9870df8_106, \2462 );
nor \U$50491 ( \50834 , \50832 , \50833 );
and \U$50492 ( \50835 , \50834 , \2468 );
not \U$50493 ( \50836 , \50834 );
and \U$50494 ( \50837 , \50836 , \2263 );
nor \U$50495 ( \50838 , \50835 , \50837 );
xor \U$50496 ( \50839 , \50831 , \50838 );
not \U$50497 ( \50840 , \3918 );
and \U$50498 ( \50841 , \3683 , RI9870c18_102);
and \U$50499 ( \50842 , RI98710c8_112, \3681 );
nor \U$50500 ( \50843 , \50841 , \50842 );
not \U$50501 ( \50844 , \50843 );
or \U$50502 ( \50845 , \50840 , \50844 );
or \U$50503 ( \50846 , \50843 , \3412 );
nand \U$50504 ( \50847 , \50845 , \50846 );
and \U$50505 ( \50848 , \50839 , \50847 );
and \U$50506 ( \50849 , \50831 , \50838 );
or \U$50507 ( \50850 , \50848 , \50849 );
and \U$50508 ( \50851 , \776 , RI9870678_90);
and \U$50509 ( \50852 , RI9870948_96, \774 );
nor \U$50510 ( \50853 , \50851 , \50852 );
and \U$50511 ( \50854 , \50853 , \474 );
not \U$50512 ( \50855 , \50853 );
and \U$50513 ( \50856 , \50855 , \451 );
nor \U$50514 ( \50857 , \50854 , \50856 );
not \U$50515 ( \50858 , \1128 );
and \U$50516 ( \50859 , \1293 , RI9870858_94);
and \U$50517 ( \50860 , RI986fb38_66, \1291 );
nor \U$50518 ( \50861 , \50859 , \50860 );
not \U$50519 ( \50862 , \50861 );
or \U$50520 ( \50863 , \50858 , \50862 );
or \U$50521 ( \50864 , \50861 , \1301 );
nand \U$50522 ( \50865 , \50863 , \50864 );
xor \U$50523 ( \50866 , \50857 , \50865 );
and \U$50524 ( \50867 , \1329 , RI986fc28_68);
and \U$50525 ( \50868 , RI986fe08_72, \1327 );
nor \U$50526 ( \50869 , \50867 , \50868 );
and \U$50527 ( \50870 , \50869 , \1336 );
not \U$50528 ( \50871 , \50869 );
and \U$50529 ( \50872 , \50871 , \1337 );
nor \U$50530 ( \50873 , \50870 , \50872 );
and \U$50531 ( \50874 , \50866 , \50873 );
and \U$50532 ( \50875 , \50857 , \50865 );
or \U$50533 ( \50876 , \50874 , \50875 );
xor \U$50534 ( \50877 , \50850 , \50876 );
and \U$50535 ( \50878 , \2274 , RI98701c8_80);
and \U$50536 ( \50879 , RI9870fd8_110, \2272 );
nor \U$50537 ( \50880 , \50878 , \50879 );
and \U$50538 ( \50881 , \50880 , \2030 );
not \U$50539 ( \50882 , \50880 );
and \U$50540 ( \50883 , \50882 , \2031 );
nor \U$50541 ( \50884 , \50881 , \50883 );
and \U$50542 ( \50885 , \1311 , RI986fd18_70);
and \U$50543 ( \50886 , RI986ffe8_76, \1309 );
nor \U$50544 ( \50887 , \50885 , \50886 );
and \U$50545 ( \50888 , \50887 , \1458 );
not \U$50546 ( \50889 , \50887 );
and \U$50547 ( \50890 , \50889 , \1318 );
nor \U$50548 ( \50891 , \50888 , \50890 );
xor \U$50549 ( \50892 , \50884 , \50891 );
not \U$50550 ( \50893 , \2034 );
and \U$50551 ( \50894 , \2042 , RI986fef8_74);
and \U$50552 ( \50895 , RI98700d8_78, \2040 );
nor \U$50553 ( \50896 , \50894 , \50895 );
not \U$50554 ( \50897 , \50896 );
or \U$50555 ( \50898 , \50893 , \50897 );
or \U$50556 ( \50899 , \50896 , \1462 );
nand \U$50557 ( \50900 , \50898 , \50899 );
and \U$50558 ( \50901 , \50892 , \50900 );
and \U$50559 ( \50902 , \50884 , \50891 );
or \U$50560 ( \50903 , \50901 , \50902 );
and \U$50561 ( \50904 , \50877 , \50903 );
and \U$50562 ( \50905 , \50850 , \50876 );
or \U$50563 ( \50906 , \50904 , \50905 );
and \U$50564 ( \50907 , \50823 , \50906 );
and \U$50565 ( \50908 , \50749 , \50822 );
or \U$50566 ( \50909 , \50907 , \50908 );
xor \U$50567 ( \50910 , \49946 , \487 );
xor \U$50568 ( \50911 , \50910 , \49954 );
xor \U$50569 ( \50912 , \49965 , \49972 );
xor \U$50570 ( \50913 , \50912 , \49980 );
and \U$50571 ( \50914 , \50911 , \50913 );
xor \U$50572 ( \50915 , \50365 , \50372 );
xor \U$50573 ( \50916 , \50915 , \50380 );
xor \U$50574 ( \50917 , \50421 , \50429 );
xor \U$50575 ( \50918 , \50917 , \50437 );
xor \U$50576 ( \50919 , \50916 , \50918 );
not \U$50577 ( \50920 , \50390 );
xor \U$50578 ( \50921 , \50408 , \50398 );
not \U$50579 ( \50922 , \50921 );
or \U$50580 ( \50923 , \50920 , \50922 );
or \U$50581 ( \50924 , \50921 , \50390 );
nand \U$50582 ( \50925 , \50923 , \50924 );
and \U$50583 ( \50926 , \50919 , \50925 );
and \U$50584 ( \50927 , \50916 , \50918 );
or \U$50585 ( \50928 , \50926 , \50927 );
xor \U$50586 ( \50929 , \49965 , \49972 );
xor \U$50587 ( \50930 , \50929 , \49980 );
and \U$50588 ( \50931 , \50928 , \50930 );
and \U$50589 ( \50932 , \50911 , \50928 );
or \U$50590 ( \50933 , \50914 , \50931 , \50932 );
xor \U$50591 ( \50934 , \50909 , \50933 );
not \U$50592 ( \50935 , \50219 );
xor \U$50593 ( \50936 , \50227 , \50237 );
not \U$50594 ( \50937 , \50936 );
or \U$50595 ( \50938 , \50935 , \50937 );
or \U$50596 ( \50939 , \50936 , \50219 );
nand \U$50597 ( \50940 , \50938 , \50939 );
xor \U$50598 ( \50941 , \50248 , \50256 );
xor \U$50599 ( \50942 , \50941 , \50265 );
xor \U$50600 ( \50943 , \50940 , \50942 );
xor \U$50601 ( \50944 , \50193 , \50200 );
xor \U$50602 ( \50945 , \50944 , \50208 );
and \U$50603 ( \50946 , \50943 , \50945 );
and \U$50604 ( \50947 , \50940 , \50942 );
or \U$50605 ( \50948 , \50946 , \50947 );
not \U$50606 ( \50949 , \367 );
and \U$50607 ( \50950 , \376 , RI9870498_86);
and \U$50608 ( \50951 , RI9870588_88, \374 );
nor \U$50609 ( \50952 , \50950 , \50951 );
not \U$50610 ( \50953 , \50952 );
or \U$50611 ( \50954 , \50949 , \50953 );
or \U$50612 ( \50955 , \50952 , \365 );
nand \U$50613 ( \50956 , \50954 , \50955 );
not \U$50614 ( \50957 , \454 );
and \U$50615 ( \50958 , \465 , RI98703a8_84);
and \U$50616 ( \50959 , RI98702b8_82, \463 );
nor \U$50617 ( \50960 , \50958 , \50959 );
not \U$50618 ( \50961 , \50960 );
or \U$50619 ( \50962 , \50957 , \50961 );
or \U$50620 ( \50963 , \50960 , \454 );
nand \U$50621 ( \50964 , \50962 , \50963 );
xor \U$50622 ( \50965 , \50956 , \50964 );
not \U$50623 ( \50966 , \456 );
and \U$50624 ( \50967 , \465 , RI9870588_88);
and \U$50625 ( \50968 , RI98703a8_84, \463 );
nor \U$50626 ( \50969 , \50967 , \50968 );
not \U$50627 ( \50970 , \50969 );
or \U$50628 ( \50971 , \50966 , \50970 );
or \U$50629 ( \50972 , \50969 , \454 );
nand \U$50630 ( \50973 , \50971 , \50972 );
nand \U$50631 ( \50974 , RI9870498_86, \374 );
not \U$50632 ( \50975 , \50974 );
not \U$50633 ( \50976 , \365 );
or \U$50634 ( \50977 , \50975 , \50976 );
or \U$50635 ( \50978 , \365 , \50974 );
nand \U$50636 ( \50979 , \50977 , \50978 );
xor \U$50637 ( \50980 , \50973 , \50979 );
and \U$50638 ( \50981 , \438 , RI98702b8_82);
and \U$50639 ( \50982 , RI9870768_92, \436 );
nor \U$50640 ( \50983 , \50981 , \50982 );
and \U$50641 ( \50984 , \50983 , \444 );
not \U$50642 ( \50985 , \50983 );
and \U$50643 ( \50986 , \50985 , \443 );
nor \U$50644 ( \50987 , \50984 , \50986 );
and \U$50645 ( \50988 , \50980 , \50987 );
and \U$50646 ( \50989 , \50973 , \50979 );
or \U$50647 ( \50990 , \50988 , \50989 );
and \U$50648 ( \50991 , \50965 , \50990 );
and \U$50649 ( \50992 , \50956 , \50964 );
or \U$50650 ( \50993 , \50991 , \50992 );
xor \U$50651 ( \50994 , \50948 , \50993 );
not \U$50652 ( \50995 , \50286 );
xor \U$50653 ( \50996 , \50278 , \50297 );
not \U$50654 ( \50997 , \50996 );
or \U$50655 ( \50998 , \50995 , \50997 );
or \U$50656 ( \50999 , \50996 , \50286 );
nand \U$50657 ( \51000 , \50998 , \50999 );
xor \U$50658 ( \51001 , \50336 , \50343 );
xor \U$50659 ( \51002 , \51001 , \50352 );
xor \U$50660 ( \51003 , \51000 , \51002 );
xor \U$50661 ( \51004 , \50306 , \50314 );
xor \U$50662 ( \51005 , \51004 , \50322 );
and \U$50663 ( \51006 , \51003 , \51005 );
and \U$50664 ( \51007 , \51000 , \51002 );
or \U$50665 ( \51008 , \51006 , \51007 );
and \U$50666 ( \51009 , \50994 , \51008 );
and \U$50667 ( \51010 , \50948 , \50993 );
or \U$50668 ( \51011 , \51009 , \51010 );
and \U$50669 ( \51012 , \50934 , \51011 );
and \U$50670 ( \51013 , \50909 , \50933 );
or \U$50671 ( \51014 , \51012 , \51013 );
nand \U$50672 ( \51015 , \50669 , \51014 );
nand \U$50673 ( \51016 , \50668 , \51015 );
xor \U$50674 ( \51017 , \50583 , \51016 );
xor \U$50675 ( \51018 , \49747 , \49759 );
xor \U$50676 ( \51019 , \51018 , \49764 );
xor \U$50677 ( \51020 , \50544 , \50551 );
xor \U$50678 ( \51021 , \51019 , \51020 );
and \U$50679 ( \51022 , \51017 , \51021 );
and \U$50680 ( \51023 , \50583 , \51016 );
or \U$50681 ( \51024 , \51022 , \51023 );
xor \U$50682 ( \51025 , \50163 , \50165 );
xor \U$50683 ( \51026 , \51025 , \50168 );
and \U$50684 ( \51027 , \51024 , \51026 );
xor \U$50685 ( \51028 , \50539 , \50541 );
xor \U$50686 ( \51029 , \51028 , \50556 );
xor \U$50687 ( \51030 , \50163 , \50165 );
xor \U$50688 ( \51031 , \51030 , \50168 );
and \U$50689 ( \51032 , \51029 , \51031 );
and \U$50690 ( \51033 , \51024 , \51029 );
or \U$50691 ( \51034 , \51027 , \51032 , \51033 );
xor \U$50692 ( \51035 , \50112 , \50126 );
xor \U$50693 ( \51036 , \51035 , \50131 );
xor \U$50694 ( \51037 , \51034 , \51036 );
xor \U$50695 ( \51038 , \50159 , \50171 );
xor \U$50696 ( \51039 , \51038 , \50559 );
and \U$50697 ( \51040 , \51037 , \51039 );
and \U$50698 ( \51041 , \51034 , \51036 );
or \U$50699 ( \51042 , \51040 , \51041 );
and \U$50700 ( \51043 , \50569 , \51042 );
xor \U$50701 ( \51044 , \51042 , \50569 );
xor \U$50702 ( \51045 , \50474 , \50490 );
xor \U$50703 ( \51046 , \51045 , \50505 );
xor \U$50704 ( \51047 , \50271 , \50357 );
xor \U$50705 ( \51048 , \51047 , \50442 );
xor \U$50706 ( \51049 , \50447 , \50449 );
xor \U$50707 ( \51050 , \51049 , \50454 );
xor \U$50708 ( \51051 , \50585 , \50592 );
xor \U$50709 ( \51052 , \51050 , \51051 );
xor \U$50710 ( \51053 , \51048 , \51052 );
xor \U$50711 ( \51054 , \51046 , \51053 );
xor \U$50712 ( \51055 , \50909 , \50933 );
xor \U$50713 ( \51056 , \51055 , \51011 );
and \U$50714 ( \51057 , \51054 , \51056 );
not \U$50715 ( \51058 , \51054 );
not \U$50716 ( \51059 , \51056 );
and \U$50717 ( \51060 , \51058 , \51059 );
xor \U$50718 ( \51061 , \50801 , \50808 );
xor \U$50719 ( \51062 , \51061 , \50816 );
xor \U$50720 ( \51063 , \50676 , \50683 );
xor \U$50721 ( \51064 , \51063 , \50691 );
and \U$50722 ( \51065 , \51062 , \51064 );
xor \U$50723 ( \51066 , \50756 , \50763 );
xor \U$50724 ( \51067 , \51066 , \50771 );
xor \U$50725 ( \51068 , \50676 , \50683 );
xor \U$50726 ( \51069 , \51068 , \50691 );
and \U$50727 ( \51070 , \51067 , \51069 );
and \U$50728 ( \51071 , \51062 , \51067 );
or \U$50729 ( \51072 , \51065 , \51070 , \51071 );
xor \U$50730 ( \51073 , \50728 , \50735 );
xor \U$50731 ( \51074 , \51073 , \50743 );
xor \U$50732 ( \51075 , \50831 , \50838 );
xor \U$50733 ( \51076 , \51075 , \50847 );
xor \U$50734 ( \51077 , \51074 , \51076 );
xor \U$50735 ( \51078 , \50701 , \50708 );
xor \U$50736 ( \51079 , \51078 , \50717 );
and \U$50737 ( \51080 , \51077 , \51079 );
and \U$50738 ( \51081 , \51074 , \51076 );
or \U$50739 ( \51082 , \51080 , \51081 );
xor \U$50740 ( \51083 , \51072 , \51082 );
xor \U$50741 ( \51084 , \50857 , \50865 );
xor \U$50742 ( \51085 , \51084 , \50873 );
xor \U$50743 ( \51086 , \50973 , \50979 );
xor \U$50744 ( \51087 , \51086 , \50987 );
and \U$50745 ( \51088 , \51085 , \51087 );
xor \U$50746 ( \51089 , \50884 , \50891 );
xor \U$50747 ( \51090 , \51089 , \50900 );
xor \U$50748 ( \51091 , \50973 , \50979 );
xor \U$50749 ( \51092 , \51091 , \50987 );
and \U$50750 ( \51093 , \51090 , \51092 );
and \U$50751 ( \51094 , \51085 , \51090 );
or \U$50752 ( \51095 , \51088 , \51093 , \51094 );
and \U$50753 ( \51096 , \51083 , \51095 );
and \U$50754 ( \51097 , \51072 , \51082 );
or \U$50755 ( \51098 , \51096 , \51097 );
and \U$50756 ( \51099 , \1311 , RI986fe08_72);
and \U$50757 ( \51100 , RI986fd18_70, \1309 );
nor \U$50758 ( \51101 , \51099 , \51100 );
and \U$50759 ( \51102 , \51101 , \1315 );
not \U$50760 ( \51103 , \51101 );
and \U$50761 ( \51104 , \51103 , \1319 );
nor \U$50762 ( \51105 , \51102 , \51104 );
and \U$50763 ( \51106 , \2042 , RI986ffe8_76);
and \U$50764 ( \51107 , RI986fef8_74, \2040 );
nor \U$50765 ( \51108 , \51106 , \51107 );
not \U$50766 ( \51109 , \51108 );
not \U$50767 ( \51110 , \2034 );
and \U$50768 ( \51111 , \51109 , \51110 );
and \U$50769 ( \51112 , \51108 , \1462 );
nor \U$50770 ( \51113 , \51111 , \51112 );
xor \U$50771 ( \51114 , \51105 , \51113 );
and \U$50772 ( \51115 , \1329 , RI986fb38_66);
and \U$50773 ( \51116 , RI986fc28_68, \1327 );
nor \U$50774 ( \51117 , \51115 , \51116 );
and \U$50775 ( \51118 , \51117 , \1337 );
not \U$50776 ( \51119 , \51117 );
and \U$50777 ( \51120 , \51119 , \1336 );
nor \U$50778 ( \51121 , \51118 , \51120 );
and \U$50779 ( \51122 , \51114 , \51121 );
and \U$50780 ( \51123 , \51105 , \51113 );
nor \U$50781 ( \51124 , \51122 , \51123 );
not \U$50782 ( \51125 , \1301 );
and \U$50783 ( \51126 , \1293 , RI9870948_96);
and \U$50784 ( \51127 , RI9870858_94, \1291 );
nor \U$50785 ( \51128 , \51126 , \51127 );
not \U$50786 ( \51129 , \51128 );
or \U$50787 ( \51130 , \51125 , \51129 );
or \U$50788 ( \51131 , \51128 , \1128 );
nand \U$50789 ( \51132 , \51130 , \51131 );
and \U$50790 ( \51133 , \776 , RI9870768_92);
and \U$50791 ( \51134 , RI9870678_90, \774 );
nor \U$50792 ( \51135 , \51133 , \51134 );
and \U$50793 ( \51136 , \51135 , \474 );
not \U$50794 ( \51137 , \51135 );
and \U$50795 ( \51138 , \51137 , \451 );
nor \U$50796 ( \51139 , \51136 , \51138 );
xor \U$50797 ( \51140 , \51132 , \51139 );
and \U$50798 ( \51141 , \438 , RI98703a8_84);
and \U$50799 ( \51142 , RI98702b8_82, \436 );
nor \U$50800 ( \51143 , \51141 , \51142 );
and \U$50801 ( \51144 , \51143 , \444 );
not \U$50802 ( \51145 , \51143 );
and \U$50803 ( \51146 , \51145 , \443 );
nor \U$50804 ( \51147 , \51144 , \51146 );
and \U$50805 ( \51148 , \51140 , \51147 );
and \U$50806 ( \51149 , \51132 , \51139 );
or \U$50807 ( \51150 , \51148 , \51149 );
xor \U$50808 ( \51151 , \51124 , \51150 );
and \U$50809 ( \51152 , \2464 , RI9870fd8_110);
and \U$50810 ( \51153 , RI9870b28_100, \2462 );
nor \U$50811 ( \51154 , \51152 , \51153 );
and \U$50812 ( \51155 , \51154 , \2468 );
not \U$50813 ( \51156 , \51154 );
and \U$50814 ( \51157 , \51156 , \2263 );
nor \U$50815 ( \51158 , \51155 , \51157 );
and \U$50816 ( \51159 , \2274 , RI98700d8_78);
and \U$50817 ( \51160 , RI98701c8_80, \2272 );
nor \U$50818 ( \51161 , \51159 , \51160 );
and \U$50819 ( \51162 , \51161 , \2030 );
not \U$50820 ( \51163 , \51161 );
and \U$50821 ( \51164 , \51163 , \2031 );
nor \U$50822 ( \51165 , \51162 , \51164 );
xor \U$50823 ( \51166 , \51158 , \51165 );
not \U$50824 ( \51167 , \2935 );
and \U$50825 ( \51168 , \3254 , RI9870df8_106);
and \U$50826 ( \51169 , RI9870a38_98, \3252 );
nor \U$50827 ( \51170 , \51168 , \51169 );
not \U$50828 ( \51171 , \51170 );
or \U$50829 ( \51172 , \51167 , \51171 );
or \U$50830 ( \51173 , \51170 , \2935 );
nand \U$50831 ( \51174 , \51172 , \51173 );
and \U$50832 ( \51175 , \51166 , \51174 );
and \U$50833 ( \51176 , \51158 , \51165 );
or \U$50834 ( \51177 , \51175 , \51176 );
and \U$50835 ( \51178 , \51151 , \51177 );
and \U$50836 ( \51179 , \51124 , \51150 );
or \U$50837 ( \51180 , \51178 , \51179 );
and \U$50838 ( \51181 , \9237 , RI986ec38_34);
and \U$50839 ( \51182 , RI986ed28_36, \9235 );
nor \U$50840 ( \51183 , \51181 , \51182 );
and \U$50841 ( \51184 , \51183 , \8836 );
not \U$50842 ( \51185 , \51183 );
and \U$50843 ( \51186 , \51185 , \9241 );
nor \U$50844 ( \51187 , \51184 , \51186 );
and \U$50845 ( \51188 , \9505 , RI986f0e8_44);
and \U$50846 ( \51189 , RI986eff8_42, \9503 );
nor \U$50847 ( \51190 , \51188 , \51189 );
and \U$50848 ( \51191 , \51190 , \9513 );
not \U$50849 ( \51192 , \51190 );
and \U$50850 ( \51193 , \51192 , \9510 );
nor \U$50851 ( \51194 , \51191 , \51193 );
or \U$50852 ( \51195 , \51187 , \51194 );
not \U$50853 ( \51196 , \51194 );
not \U$50854 ( \51197 , \51187 );
or \U$50855 ( \51198 , \51196 , \51197 );
and \U$50856 ( \51199 , \10424 , RI986f2c8_48);
and \U$50857 ( \51200 , RI986f1d8_46, \10422 );
nor \U$50858 ( \51201 , \51199 , \51200 );
and \U$50859 ( \51202 , \51201 , \9840 );
not \U$50860 ( \51203 , \51201 );
and \U$50861 ( \51204 , \51203 , \10428 );
nor \U$50862 ( \51205 , \51202 , \51204 );
nand \U$50863 ( \51206 , \51198 , \51205 );
nand \U$50864 ( \51207 , \51195 , \51206 );
and \U$50865 ( \51208 , \15780 , RI986f598_54);
and \U$50866 ( \51209 , RI986f688_56, RI9873648_192);
nor \U$50867 ( \51210 , \51208 , \51209 );
not \U$50868 ( \51211 , \51210 );
not \U$50869 ( \51212 , RI9873558_190);
and \U$50870 ( \51213 , \51211 , \51212 );
and \U$50871 ( \51214 , \51210 , RI9873558_190);
nor \U$50872 ( \51215 , \51213 , \51214 );
and \U$50873 ( \51216 , \14937 , RI986f4a8_52);
and \U$50874 ( \51217 , RI986f3b8_50, \14935 );
nor \U$50875 ( \51218 , \51216 , \51217 );
and \U$50876 ( \51219 , \51218 , \14538 );
not \U$50877 ( \51220 , \51218 );
and \U$50878 ( \51221 , \51220 , \14539 );
nor \U$50879 ( \51222 , \51219 , \51221 );
xor \U$50880 ( \51223 , \51215 , \51222 );
and \U$50881 ( \51224 , \13882 , RI986fa48_64);
and \U$50882 ( \51225 , RI986f958_62, \13880 );
nor \U$50883 ( \51226 , \51224 , \51225 );
and \U$50884 ( \51227 , \51226 , \13359 );
not \U$50885 ( \51228 , \51226 );
and \U$50886 ( \51229 , \51228 , \13358 );
nor \U$50887 ( \51230 , \51227 , \51229 );
and \U$50888 ( \51231 , \51223 , \51230 );
and \U$50889 ( \51232 , \51215 , \51222 );
nor \U$50890 ( \51233 , \51231 , \51232 );
xor \U$50891 ( \51234 , \51207 , \51233 );
and \U$50892 ( \51235 , \12293 , RI986e788_24);
and \U$50893 ( \51236 , RI986e698_22, \12291 );
nor \U$50894 ( \51237 , \51235 , \51236 );
and \U$50895 ( \51238 , \51237 , \11686 );
not \U$50896 ( \51239 , \51237 );
and \U$50897 ( \51240 , \51239 , \11687 );
nor \U$50898 ( \51241 , \51238 , \51240 );
and \U$50899 ( \51242 , \13045 , RI986f868_60);
and \U$50900 ( \51243 , RI986f778_58, \13043 );
nor \U$50901 ( \51244 , \51242 , \51243 );
and \U$50902 ( \51245 , \51244 , \12619 );
not \U$50903 ( \51246 , \51244 );
and \U$50904 ( \51247 , \51246 , \13047 );
nor \U$50905 ( \51248 , \51245 , \51247 );
xor \U$50906 ( \51249 , \51241 , \51248 );
and \U$50907 ( \51250 , \11696 , RI986e5a8_20);
and \U$50908 ( \51251 , RI986e4b8_18, \11694 );
nor \U$50909 ( \51252 , \51250 , \51251 );
and \U$50910 ( \51253 , \51252 , \11702 );
not \U$50911 ( \51254 , \51252 );
and \U$50912 ( \51255 , \51254 , \10965 );
nor \U$50913 ( \51256 , \51253 , \51255 );
and \U$50914 ( \51257 , \51249 , \51256 );
and \U$50915 ( \51258 , \51241 , \51248 );
nor \U$50916 ( \51259 , \51257 , \51258 );
and \U$50917 ( \51260 , \51234 , \51259 );
and \U$50918 ( \51261 , \51207 , \51233 );
or \U$50919 ( \51262 , \51260 , \51261 );
xor \U$50920 ( \51263 , \51180 , \51262 );
and \U$50921 ( \51264 , \7729 , RI986e968_28);
and \U$50922 ( \51265 , RI986e878_26, \7727 );
nor \U$50923 ( \51266 , \51264 , \51265 );
and \U$50924 ( \51267 , \51266 , \7733 );
not \U$50925 ( \51268 , \51266 );
and \U$50926 ( \51269 , \51268 , \7480 );
nor \U$50927 ( \51270 , \51267 , \51269 );
and \U$50928 ( \51271 , \8486 , RI986ef08_40);
and \U$50929 ( \51272 , RI986ee18_38, \8484 );
nor \U$50930 ( \51273 , \51271 , \51272 );
and \U$50931 ( \51274 , \51273 , \8051 );
not \U$50932 ( \51275 , \51273 );
and \U$50933 ( \51276 , \51275 , \8050 );
nor \U$50934 ( \51277 , \51274 , \51276 );
xor \U$50935 ( \51278 , \51270 , \51277 );
and \U$50936 ( \51279 , \7079 , RI986eb48_32);
and \U$50937 ( \51280 , RI986ea58_30, \7077 );
nor \U$50938 ( \51281 , \51279 , \51280 );
and \U$50939 ( \51282 , \51281 , \6709 );
not \U$50940 ( \51283 , \51281 );
and \U$50941 ( \51284 , \51283 , \6710 );
nor \U$50942 ( \51285 , \51282 , \51284 );
and \U$50943 ( \51286 , \51278 , \51285 );
and \U$50944 ( \51287 , \51270 , \51277 );
nor \U$50945 ( \51288 , \51286 , \51287 );
and \U$50946 ( \51289 , \4203 , RI98710c8_112);
and \U$50947 ( \51290 , RI9870d08_104, \4201 );
nor \U$50948 ( \51291 , \51289 , \51290 );
and \U$50949 ( \51292 , \51291 , \4207 );
not \U$50950 ( \51293 , \51291 );
and \U$50951 ( \51294 , \51293 , \3923 );
nor \U$50952 ( \51295 , \51292 , \51294 );
not \U$50953 ( \51296 , \3918 );
and \U$50954 ( \51297 , \3683 , RI9870ee8_108);
and \U$50955 ( \51298 , RI9870c18_102, \3681 );
nor \U$50956 ( \51299 , \51297 , \51298 );
not \U$50957 ( \51300 , \51299 );
or \U$50958 ( \51301 , \51296 , \51300 );
or \U$50959 ( \51302 , \51299 , \3918 );
nand \U$50960 ( \51303 , \51301 , \51302 );
xor \U$50961 ( \51304 , \51295 , \51303 );
not \U$50962 ( \51305 , \4521 );
and \U$50963 ( \51306 , \4710 , RI98712a8_116);
and \U$50964 ( \51307 , RI98711b8_114, \4708 );
nor \U$50965 ( \51308 , \51306 , \51307 );
not \U$50966 ( \51309 , \51308 );
or \U$50967 ( \51310 , \51305 , \51309 );
or \U$50968 ( \51311 , \51308 , \4521 );
nand \U$50969 ( \51312 , \51310 , \51311 );
and \U$50970 ( \51313 , \51304 , \51312 );
and \U$50971 ( \51314 , \51295 , \51303 );
or \U$50972 ( \51315 , \51313 , \51314 );
xor \U$50973 ( \51316 , \51288 , \51315 );
and \U$50974 ( \51317 , \5318 , RI9871398_118);
and \U$50975 ( \51318 , RI9871488_120, \5316 );
nor \U$50976 ( \51319 , \51317 , \51318 );
and \U$50977 ( \51320 , \51319 , \5052 );
not \U$50978 ( \51321 , \51319 );
and \U$50979 ( \51322 , \51321 , \5322 );
nor \U$50980 ( \51323 , \51320 , \51322 );
and \U$50981 ( \51324 , \5881 , RI9871758_126);
and \U$50982 ( \51325 , RI9871848_128, \5879 );
nor \U$50983 ( \51326 , \51324 , \51325 );
and \U$50984 ( \51327 , \51326 , \5594 );
not \U$50985 ( \51328 , \51326 );
and \U$50986 ( \51329 , \51328 , \5885 );
nor \U$50987 ( \51330 , \51327 , \51329 );
xor \U$50988 ( \51331 , \51323 , \51330 );
and \U$50989 ( \51332 , \6453 , RI9871578_122);
and \U$50990 ( \51333 , RI9871668_124, \6451 );
nor \U$50991 ( \51334 , \51332 , \51333 );
and \U$50992 ( \51335 , \51334 , \6190 );
not \U$50993 ( \51336 , \51334 );
and \U$50994 ( \51337 , \51336 , \6705 );
nor \U$50995 ( \51338 , \51335 , \51337 );
and \U$50996 ( \51339 , \51331 , \51338 );
and \U$50997 ( \51340 , \51323 , \51330 );
or \U$50998 ( \51341 , \51339 , \51340 );
and \U$50999 ( \51342 , \51316 , \51341 );
and \U$51000 ( \51343 , \51288 , \51315 );
or \U$51001 ( \51344 , \51342 , \51343 );
and \U$51002 ( \51345 , \51263 , \51344 );
and \U$51003 ( \51346 , \51180 , \51262 );
or \U$51004 ( \51347 , \51345 , \51346 );
xor \U$51005 ( \51348 , \51098 , \51347 );
xor \U$51006 ( \51349 , \51000 , \51002 );
xor \U$51007 ( \51350 , \51349 , \51005 );
xor \U$51008 ( \51351 , \50940 , \50942 );
xor \U$51009 ( \51352 , \51351 , \50945 );
and \U$51010 ( \51353 , \51350 , \51352 );
xor \U$51011 ( \51354 , \50916 , \50918 );
xor \U$51012 ( \51355 , \51354 , \50925 );
xor \U$51013 ( \51356 , \50940 , \50942 );
xor \U$51014 ( \51357 , \51356 , \50945 );
and \U$51015 ( \51358 , \51355 , \51357 );
and \U$51016 ( \51359 , \51350 , \51355 );
or \U$51017 ( \51360 , \51353 , \51358 , \51359 );
and \U$51018 ( \51361 , \51348 , \51360 );
and \U$51019 ( \51362 , \51098 , \51347 );
nor \U$51020 ( \51363 , \51361 , \51362 );
not \U$51021 ( \51364 , \51363 );
xor \U$51022 ( \51365 , \50749 , \50822 );
xor \U$51023 ( \51366 , \51365 , \50906 );
xor \U$51024 ( \51367 , \50948 , \50993 );
xor \U$51025 ( \51368 , \51367 , \51008 );
and \U$51026 ( \51369 , \51366 , \51368 );
xor \U$51027 ( \51370 , \49965 , \49972 );
xor \U$51028 ( \51371 , \51370 , \49980 );
xor \U$51029 ( \51372 , \50911 , \50928 );
xor \U$51030 ( \51373 , \51371 , \51372 );
xor \U$51031 ( \51374 , \50948 , \50993 );
xor \U$51032 ( \51375 , \51374 , \51008 );
and \U$51033 ( \51376 , \51373 , \51375 );
and \U$51034 ( \51377 , \51366 , \51373 );
or \U$51035 ( \51378 , \51369 , \51376 , \51377 );
not \U$51036 ( \51379 , \51378 );
or \U$51037 ( \51380 , \51364 , \51379 );
or \U$51038 ( \51381 , \51378 , \51363 );
nand \U$51039 ( \51382 , \51380 , \51381 );
not \U$51040 ( \51383 , \51382 );
not \U$51041 ( \51384 , \50608 );
xor \U$51042 ( \51385 , \50619 , \50632 );
not \U$51043 ( \51386 , \51385 );
or \U$51044 ( \51387 , \51384 , \51386 );
or \U$51045 ( \51388 , \51385 , \50608 );
nand \U$51046 ( \51389 , \51387 , \51388 );
xor \U$51047 ( \51390 , \50956 , \50964 );
xor \U$51048 ( \51391 , \51390 , \50990 );
xor \U$51049 ( \51392 , \50694 , \50720 );
xor \U$51050 ( \51393 , \51392 , \50746 );
and \U$51051 ( \51394 , \51391 , \51393 );
xor \U$51052 ( \51395 , \50850 , \50876 );
xor \U$51053 ( \51396 , \51395 , \50903 );
xor \U$51054 ( \51397 , \50694 , \50720 );
xor \U$51055 ( \51398 , \51397 , \50746 );
and \U$51056 ( \51399 , \51396 , \51398 );
and \U$51057 ( \51400 , \51391 , \51396 );
or \U$51058 ( \51401 , \51394 , \51399 , \51400 );
xor \U$51059 ( \51402 , \51389 , \51401 );
xor \U$51060 ( \51403 , \50497 , \50499 );
xor \U$51061 ( \51404 , \51403 , \50502 );
xor \U$51062 ( \51405 , \50652 , \50659 );
xor \U$51063 ( \51406 , \51404 , \51405 );
and \U$51064 ( \51407 , \51402 , \51406 );
and \U$51065 ( \51408 , \51389 , \51401 );
nor \U$51066 ( \51409 , \51407 , \51408 );
not \U$51067 ( \51410 , \51409 );
and \U$51068 ( \51411 , \51383 , \51410 );
and \U$51069 ( \51412 , \51382 , \51409 );
nor \U$51070 ( \51413 , \51411 , \51412 );
nor \U$51071 ( \51414 , \51060 , \51413 );
nor \U$51072 ( \51415 , \51057 , \51414 );
xnor \U$51073 ( \51416 , \51014 , \50666 );
not \U$51074 ( \51417 , \51416 );
not \U$51075 ( \51418 , \50597 );
and \U$51076 ( \51419 , \51417 , \51418 );
and \U$51077 ( \51420 , \51416 , \50597 );
nor \U$51078 ( \51421 , \51419 , \51420 );
xor \U$51079 ( \51422 , \51415 , \51421 );
xor \U$51080 ( \51423 , \51124 , \51150 );
xor \U$51081 ( \51424 , \51423 , \51177 );
xor \U$51082 ( \51425 , \51288 , \51315 );
xor \U$51083 ( \51426 , \51425 , \51341 );
and \U$51084 ( \51427 , \51424 , \51426 );
xor \U$51085 ( \51428 , \50973 , \50979 );
xor \U$51086 ( \51429 , \51428 , \50987 );
xor \U$51087 ( \51430 , \51085 , \51090 );
xor \U$51088 ( \51431 , \51429 , \51430 );
xor \U$51089 ( \51432 , \51288 , \51315 );
xor \U$51090 ( \51433 , \51432 , \51341 );
and \U$51091 ( \51434 , \51431 , \51433 );
and \U$51092 ( \51435 , \51424 , \51431 );
or \U$51093 ( \51436 , \51427 , \51434 , \51435 );
xor \U$51094 ( \51437 , \50774 , \50793 );
xor \U$51095 ( \51438 , \51437 , \50819 );
xor \U$51096 ( \51439 , \51436 , \51438 );
xor \U$51097 ( \51440 , \50694 , \50720 );
xor \U$51098 ( \51441 , \51440 , \50746 );
xor \U$51099 ( \51442 , \51391 , \51396 );
xor \U$51100 ( \51443 , \51441 , \51442 );
and \U$51101 ( \51444 , \51439 , \51443 );
and \U$51102 ( \51445 , \51436 , \51438 );
or \U$51103 ( \51446 , \51444 , \51445 );
xor \U$51104 ( \51447 , \51158 , \51165 );
xor \U$51105 ( \51448 , \51447 , \51174 );
xor \U$51106 ( \51449 , \51323 , \51330 );
xor \U$51107 ( \51450 , \51449 , \51338 );
and \U$51108 ( \51451 , \51448 , \51450 );
xor \U$51109 ( \51452 , \51295 , \51303 );
xor \U$51110 ( \51453 , \51452 , \51312 );
xor \U$51111 ( \51454 , \51323 , \51330 );
xor \U$51112 ( \51455 , \51454 , \51338 );
and \U$51113 ( \51456 , \51453 , \51455 );
and \U$51114 ( \51457 , \51448 , \51453 );
or \U$51115 ( \51458 , \51451 , \51456 , \51457 );
xor \U$51116 ( \51459 , \51105 , \51113 );
xor \U$51117 ( \51460 , \51459 , \51121 );
and \U$51118 ( \51461 , \465 , RI9870498_86);
and \U$51119 ( \51462 , RI9870588_88, \463 );
nor \U$51120 ( \51463 , \51461 , \51462 );
not \U$51121 ( \51464 , \51463 );
not \U$51122 ( \51465 , \456 );
and \U$51123 ( \51466 , \51464 , \51465 );
and \U$51124 ( \51467 , \51463 , \454 );
nor \U$51125 ( \51468 , \51466 , \51467 );
or \U$51126 ( \51469 , \51460 , \51468 );
not \U$51127 ( \51470 , \51468 );
not \U$51128 ( \51471 , \51460 );
or \U$51129 ( \51472 , \51470 , \51471 );
xor \U$51130 ( \51473 , \51132 , \51139 );
xor \U$51131 ( \51474 , \51473 , \51147 );
nand \U$51132 ( \51475 , \51472 , \51474 );
nand \U$51133 ( \51476 , \51469 , \51475 );
xor \U$51134 ( \51477 , \51458 , \51476 );
xor \U$51135 ( \51478 , \51270 , \51277 );
xor \U$51136 ( \51479 , \51478 , \51285 );
not \U$51137 ( \51480 , \51194 );
not \U$51138 ( \51481 , \51205 );
or \U$51139 ( \51482 , \51480 , \51481 );
or \U$51140 ( \51483 , \51194 , \51205 );
nand \U$51141 ( \51484 , \51482 , \51483 );
not \U$51142 ( \51485 , \51484 );
not \U$51143 ( \51486 , \51187 );
and \U$51144 ( \51487 , \51485 , \51486 );
and \U$51145 ( \51488 , \51484 , \51187 );
nor \U$51146 ( \51489 , \51487 , \51488 );
xor \U$51147 ( \51490 , \51479 , \51489 );
xor \U$51148 ( \51491 , \51241 , \51248 );
xor \U$51149 ( \51492 , \51491 , \51256 );
and \U$51150 ( \51493 , \51490 , \51492 );
and \U$51151 ( \51494 , \51479 , \51489 );
nor \U$51152 ( \51495 , \51493 , \51494 );
and \U$51153 ( \51496 , \51477 , \51495 );
and \U$51154 ( \51497 , \51458 , \51476 );
or \U$51155 ( \51498 , \51496 , \51497 );
and \U$51156 ( \51499 , \776 , RI98702b8_82);
and \U$51157 ( \51500 , RI9870768_92, \774 );
nor \U$51158 ( \51501 , \51499 , \51500 );
and \U$51159 ( \51502 , \51501 , \451 );
not \U$51160 ( \51503 , \51501 );
and \U$51161 ( \51504 , \51503 , \474 );
nor \U$51162 ( \51505 , \51502 , \51504 );
not \U$51163 ( \51506 , \51505 );
and \U$51164 ( \51507 , \1329 , RI9870858_94);
and \U$51165 ( \51508 , RI986fb38_66, \1327 );
nor \U$51166 ( \51509 , \51507 , \51508 );
and \U$51167 ( \51510 , \51509 , \1337 );
not \U$51168 ( \51511 , \51509 );
and \U$51169 ( \51512 , \51511 , \1336 );
nor \U$51170 ( \51513 , \51510 , \51512 );
not \U$51171 ( \51514 , \51513 );
and \U$51172 ( \51515 , \51506 , \51514 );
and \U$51173 ( \51516 , \51513 , \51505 );
and \U$51174 ( \51517 , \1293 , RI9870678_90);
and \U$51175 ( \51518 , RI9870948_96, \1291 );
nor \U$51176 ( \51519 , \51517 , \51518 );
not \U$51177 ( \51520 , \51519 );
not \U$51178 ( \51521 , \1301 );
and \U$51179 ( \51522 , \51520 , \51521 );
and \U$51180 ( \51523 , \51519 , \1301 );
nor \U$51181 ( \51524 , \51522 , \51523 );
nor \U$51182 ( \51525 , \51516 , \51524 );
nor \U$51183 ( \51526 , \51515 , \51525 );
and \U$51184 ( \51527 , \3683 , RI9870a38_98);
and \U$51185 ( \51528 , RI9870ee8_108, \3681 );
nor \U$51186 ( \51529 , \51527 , \51528 );
not \U$51187 ( \51530 , \51529 );
not \U$51188 ( \51531 , \3412 );
and \U$51189 ( \51532 , \51530 , \51531 );
and \U$51190 ( \51533 , \51529 , \3412 );
nor \U$51191 ( \51534 , \51532 , \51533 );
and \U$51192 ( \51535 , \2464 , RI98701c8_80);
and \U$51193 ( \51536 , RI9870fd8_110, \2462 );
nor \U$51194 ( \51537 , \51535 , \51536 );
and \U$51195 ( \51538 , \51537 , \2263 );
not \U$51196 ( \51539 , \51537 );
and \U$51197 ( \51540 , \51539 , \2468 );
nor \U$51198 ( \51541 , \51538 , \51540 );
xor \U$51199 ( \51542 , \51534 , \51541 );
and \U$51200 ( \51543 , \3254 , RI9870b28_100);
and \U$51201 ( \51544 , RI9870df8_106, \3252 );
nor \U$51202 ( \51545 , \51543 , \51544 );
not \U$51203 ( \51546 , \51545 );
not \U$51204 ( \51547 , \2935 );
and \U$51205 ( \51548 , \51546 , \51547 );
and \U$51206 ( \51549 , \51545 , \3406 );
nor \U$51207 ( \51550 , \51548 , \51549 );
and \U$51208 ( \51551 , \51542 , \51550 );
and \U$51209 ( \51552 , \51534 , \51541 );
or \U$51210 ( \51553 , \51551 , \51552 );
xor \U$51211 ( \51554 , \51526 , \51553 );
and \U$51212 ( \51555 , \1311 , RI986fc28_68);
and \U$51213 ( \51556 , RI986fe08_72, \1309 );
nor \U$51214 ( \51557 , \51555 , \51556 );
and \U$51215 ( \51558 , \51557 , \1315 );
not \U$51216 ( \51559 , \51557 );
and \U$51217 ( \51560 , \51559 , \1319 );
nor \U$51218 ( \51561 , \51558 , \51560 );
and \U$51219 ( \51562 , \2042 , RI986fd18_70);
and \U$51220 ( \51563 , RI986ffe8_76, \2040 );
nor \U$51221 ( \51564 , \51562 , \51563 );
not \U$51222 ( \51565 , \51564 );
not \U$51223 ( \51566 , \1462 );
and \U$51224 ( \51567 , \51565 , \51566 );
and \U$51225 ( \51568 , \51564 , \2034 );
nor \U$51226 ( \51569 , \51567 , \51568 );
xor \U$51227 ( \51570 , \51561 , \51569 );
and \U$51228 ( \51571 , \2274 , RI986fef8_74);
and \U$51229 ( \51572 , RI98700d8_78, \2272 );
nor \U$51230 ( \51573 , \51571 , \51572 );
and \U$51231 ( \51574 , \51573 , \2031 );
not \U$51232 ( \51575 , \51573 );
and \U$51233 ( \51576 , \51575 , \2030 );
nor \U$51234 ( \51577 , \51574 , \51576 );
and \U$51235 ( \51578 , \51570 , \51577 );
and \U$51236 ( \51579 , \51561 , \51569 );
or \U$51237 ( \51580 , \51578 , \51579 );
and \U$51238 ( \51581 , \51554 , \51580 );
and \U$51239 ( \51582 , \51526 , \51553 );
nor \U$51240 ( \51583 , \51581 , \51582 );
and \U$51241 ( \51584 , \10424 , RI986eff8_42);
and \U$51242 ( \51585 , RI986f2c8_48, \10422 );
nor \U$51243 ( \51586 , \51584 , \51585 );
and \U$51244 ( \51587 , \51586 , \10428 );
not \U$51245 ( \51588 , \51586 );
and \U$51246 ( \51589 , \51588 , \9840 );
nor \U$51247 ( \51590 , \51587 , \51589 );
and \U$51248 ( \51591 , \11696 , RI986f1d8_46);
and \U$51249 ( \51592 , RI986e5a8_20, \11694 );
nor \U$51250 ( \51593 , \51591 , \51592 );
and \U$51251 ( \51594 , \51593 , \11702 );
not \U$51252 ( \51595 , \51593 );
and \U$51253 ( \51596 , \51595 , \10965 );
nor \U$51254 ( \51597 , \51594 , \51596 );
xor \U$51255 ( \51598 , \51590 , \51597 );
and \U$51256 ( \51599 , \9505 , RI986ed28_36);
and \U$51257 ( \51600 , RI986f0e8_44, \9503 );
nor \U$51258 ( \51601 , \51599 , \51600 );
and \U$51259 ( \51602 , \51601 , \9513 );
not \U$51260 ( \51603 , \51601 );
and \U$51261 ( \51604 , \51603 , \9510 );
nor \U$51262 ( \51605 , \51602 , \51604 );
and \U$51263 ( \51606 , \51598 , \51605 );
and \U$51264 ( \51607 , \51590 , \51597 );
nor \U$51265 ( \51608 , \51606 , \51607 );
not \U$51266 ( \51609 , RI9873558_190);
and \U$51267 ( \51610 , \15780 , RI986f3b8_50);
and \U$51268 ( \51611 , RI986f598_54, RI9873648_192);
nor \U$51269 ( \51612 , \51610 , \51611 );
not \U$51270 ( \51613 , \51612 );
or \U$51271 ( \51614 , \51609 , \51613 );
or \U$51272 ( \51615 , \51612 , RI9873558_190);
nand \U$51273 ( \51616 , \51614 , \51615 );
xor \U$51274 ( \51617 , \51616 , \456 );
and \U$51275 ( \51618 , \14937 , RI986f958_62);
and \U$51276 ( \51619 , RI986f4a8_52, \14935 );
nor \U$51277 ( \51620 , \51618 , \51619 );
and \U$51278 ( \51621 , \51620 , \14539 );
not \U$51279 ( \51622 , \51620 );
and \U$51280 ( \51623 , \51622 , \14538 );
nor \U$51281 ( \51624 , \51621 , \51623 );
and \U$51282 ( \51625 , \51617 , \51624 );
and \U$51283 ( \51626 , \51616 , \456 );
or \U$51284 ( \51627 , \51625 , \51626 );
xor \U$51285 ( \51628 , \51608 , \51627 );
and \U$51286 ( \51629 , \13882 , RI986f778_58);
and \U$51287 ( \51630 , RI986fa48_64, \13880 );
nor \U$51288 ( \51631 , \51629 , \51630 );
and \U$51289 ( \51632 , \51631 , \13358 );
not \U$51290 ( \51633 , \51631 );
and \U$51291 ( \51634 , \51633 , \13359 );
nor \U$51292 ( \51635 , \51632 , \51634 );
and \U$51293 ( \51636 , \12293 , RI986e4b8_18);
and \U$51294 ( \51637 , RI986e788_24, \12291 );
nor \U$51295 ( \51638 , \51636 , \51637 );
and \U$51296 ( \51639 , \51638 , \11687 );
not \U$51297 ( \51640 , \51638 );
and \U$51298 ( \51641 , \51640 , \11686 );
nor \U$51299 ( \51642 , \51639 , \51641 );
xor \U$51300 ( \51643 , \51635 , \51642 );
and \U$51301 ( \51644 , \13045 , RI986e698_22);
and \U$51302 ( \51645 , RI986f868_60, \13043 );
nor \U$51303 ( \51646 , \51644 , \51645 );
and \U$51304 ( \51647 , \51646 , \13047 );
not \U$51305 ( \51648 , \51646 );
and \U$51306 ( \51649 , \51648 , \12619 );
nor \U$51307 ( \51650 , \51647 , \51649 );
and \U$51308 ( \51651 , \51643 , \51650 );
and \U$51309 ( \51652 , \51635 , \51642 );
or \U$51310 ( \51653 , \51651 , \51652 );
and \U$51311 ( \51654 , \51628 , \51653 );
and \U$51312 ( \51655 , \51608 , \51627 );
or \U$51313 ( \51656 , \51654 , \51655 );
xor \U$51314 ( \51657 , \51583 , \51656 );
and \U$51315 ( \51658 , \5881 , RI9871488_120);
and \U$51316 ( \51659 , RI9871758_126, \5879 );
nor \U$51317 ( \51660 , \51658 , \51659 );
and \U$51318 ( \51661 , \51660 , \5885 );
not \U$51319 ( \51662 , \51660 );
and \U$51320 ( \51663 , \51662 , \5594 );
nor \U$51321 ( \51664 , \51661 , \51663 );
and \U$51322 ( \51665 , \6453 , RI9871848_128);
and \U$51323 ( \51666 , RI9871578_122, \6451 );
nor \U$51324 ( \51667 , \51665 , \51666 );
and \U$51325 ( \51668 , \51667 , \6180 );
not \U$51326 ( \51669 , \51667 );
and \U$51327 ( \51670 , \51669 , \6190 );
nor \U$51328 ( \51671 , \51668 , \51670 );
xor \U$51329 ( \51672 , \51664 , \51671 );
and \U$51330 ( \51673 , \7079 , RI9871668_124);
and \U$51331 ( \51674 , RI986eb48_32, \7077 );
nor \U$51332 ( \51675 , \51673 , \51674 );
and \U$51333 ( \51676 , \51675 , \6709 );
not \U$51334 ( \51677 , \51675 );
and \U$51335 ( \51678 , \51677 , \6710 );
nor \U$51336 ( \51679 , \51676 , \51678 );
and \U$51337 ( \51680 , \51672 , \51679 );
and \U$51338 ( \51681 , \51664 , \51671 );
or \U$51339 ( \51682 , \51680 , \51681 );
and \U$51340 ( \51683 , \7729 , RI986ea58_30);
and \U$51341 ( \51684 , RI986e968_28, \7727 );
nor \U$51342 ( \51685 , \51683 , \51684 );
and \U$51343 ( \51686 , \51685 , \7733 );
not \U$51344 ( \51687 , \51685 );
and \U$51345 ( \51688 , \51687 , \7480 );
nor \U$51346 ( \51689 , \51686 , \51688 );
and \U$51347 ( \51690 , \8486 , RI986e878_26);
and \U$51348 ( \51691 , RI986ef08_40, \8484 );
nor \U$51349 ( \51692 , \51690 , \51691 );
and \U$51350 ( \51693 , \51692 , \8051 );
not \U$51351 ( \51694 , \51692 );
and \U$51352 ( \51695 , \51694 , \8050 );
nor \U$51353 ( \51696 , \51693 , \51695 );
xor \U$51354 ( \51697 , \51689 , \51696 );
and \U$51355 ( \51698 , \9237 , RI986ee18_38);
and \U$51356 ( \51699 , RI986ec38_34, \9235 );
nor \U$51357 ( \51700 , \51698 , \51699 );
and \U$51358 ( \51701 , \51700 , \8836 );
not \U$51359 ( \51702 , \51700 );
and \U$51360 ( \51703 , \51702 , \9241 );
nor \U$51361 ( \51704 , \51701 , \51703 );
and \U$51362 ( \51705 , \51697 , \51704 );
and \U$51363 ( \51706 , \51689 , \51696 );
or \U$51364 ( \51707 , \51705 , \51706 );
or \U$51365 ( \51708 , \51682 , \51707 );
not \U$51366 ( \51709 , \51682 );
not \U$51367 ( \51710 , \51707 );
or \U$51368 ( \51711 , \51709 , \51710 );
and \U$51369 ( \51712 , \4710 , RI9870d08_104);
and \U$51370 ( \51713 , RI98712a8_116, \4708 );
nor \U$51371 ( \51714 , \51712 , \51713 );
not \U$51372 ( \51715 , \51714 );
not \U$51373 ( \51716 , \4519 );
and \U$51374 ( \51717 , \51715 , \51716 );
and \U$51375 ( \51718 , \51714 , \4519 );
nor \U$51376 ( \51719 , \51717 , \51718 );
and \U$51377 ( \51720 , \5318 , RI98711b8_114);
and \U$51378 ( \51721 , RI9871398_118, \5316 );
nor \U$51379 ( \51722 , \51720 , \51721 );
and \U$51380 ( \51723 , \51722 , \5322 );
not \U$51381 ( \51724 , \51722 );
and \U$51382 ( \51725 , \51724 , \5052 );
nor \U$51383 ( \51726 , \51723 , \51725 );
xor \U$51384 ( \51727 , \51719 , \51726 );
and \U$51385 ( \51728 , \4203 , RI9870c18_102);
and \U$51386 ( \51729 , RI98710c8_112, \4201 );
nor \U$51387 ( \51730 , \51728 , \51729 );
and \U$51388 ( \51731 , \51730 , \3923 );
not \U$51389 ( \51732 , \51730 );
and \U$51390 ( \51733 , \51732 , \4207 );
nor \U$51391 ( \51734 , \51731 , \51733 );
and \U$51392 ( \51735 , \51727 , \51734 );
and \U$51393 ( \51736 , \51719 , \51726 );
nor \U$51394 ( \51737 , \51735 , \51736 );
nand \U$51395 ( \51738 , \51711 , \51737 );
nand \U$51396 ( \51739 , \51708 , \51738 );
and \U$51397 ( \51740 , \51657 , \51739 );
and \U$51398 ( \51741 , \51583 , \51656 );
or \U$51399 ( \51742 , \51740 , \51741 );
xor \U$51400 ( \51743 , \51498 , \51742 );
xor \U$51401 ( \51744 , \50782 , \367 );
xor \U$51402 ( \51745 , \51744 , \50790 );
xor \U$51403 ( \51746 , \51074 , \51076 );
xor \U$51404 ( \51747 , \51746 , \51079 );
and \U$51405 ( \51748 , \51745 , \51747 );
xor \U$51406 ( \51749 , \50676 , \50683 );
xor \U$51407 ( \51750 , \51749 , \50691 );
xor \U$51408 ( \51751 , \51062 , \51067 );
xor \U$51409 ( \51752 , \51750 , \51751 );
xor \U$51410 ( \51753 , \51074 , \51076 );
xor \U$51411 ( \51754 , \51753 , \51079 );
and \U$51412 ( \51755 , \51752 , \51754 );
and \U$51413 ( \51756 , \51745 , \51752 );
or \U$51414 ( \51757 , \51748 , \51755 , \51756 );
and \U$51415 ( \51758 , \51743 , \51757 );
and \U$51416 ( \51759 , \51498 , \51742 );
or \U$51417 ( \51760 , \51758 , \51759 );
xor \U$51418 ( \51761 , \51446 , \51760 );
xor \U$51419 ( \51762 , \51180 , \51262 );
xor \U$51420 ( \51763 , \51762 , \51344 );
xor \U$51421 ( \51764 , \51072 , \51082 );
xor \U$51422 ( \51765 , \51764 , \51095 );
and \U$51423 ( \51766 , \51763 , \51765 );
xor \U$51424 ( \51767 , \50940 , \50942 );
xor \U$51425 ( \51768 , \51767 , \50945 );
xor \U$51426 ( \51769 , \51350 , \51355 );
xor \U$51427 ( \51770 , \51768 , \51769 );
xor \U$51428 ( \51771 , \51072 , \51082 );
xor \U$51429 ( \51772 , \51771 , \51095 );
and \U$51430 ( \51773 , \51770 , \51772 );
and \U$51431 ( \51774 , \51763 , \51770 );
or \U$51432 ( \51775 , \51766 , \51773 , \51774 );
and \U$51433 ( \51776 , \51761 , \51775 );
and \U$51434 ( \51777 , \51446 , \51760 );
nor \U$51435 ( \51778 , \51776 , \51777 );
not \U$51436 ( \51779 , \50664 );
not \U$51437 ( \51780 , \50634 );
or \U$51438 ( \51781 , \51779 , \51780 );
or \U$51439 ( \51782 , \50634 , \50664 );
nand \U$51440 ( \51783 , \51781 , \51782 );
not \U$51441 ( \51784 , \51783 );
not \U$51442 ( \51785 , \50644 );
and \U$51443 ( \51786 , \51784 , \51785 );
and \U$51444 ( \51787 , \51783 , \50644 );
nor \U$51445 ( \51788 , \51786 , \51787 );
xor \U$51446 ( \51789 , \51778 , \51788 );
xor \U$51447 ( \51790 , \50948 , \50993 );
xor \U$51448 ( \51791 , \51790 , \51008 );
xor \U$51449 ( \51792 , \51366 , \51373 );
xor \U$51450 ( \51793 , \51791 , \51792 );
xor \U$51451 ( \51794 , \51098 , \51347 );
xor \U$51452 ( \51795 , \51794 , \51360 );
and \U$51453 ( \51796 , \51793 , \51795 );
xor \U$51454 ( \51797 , \51389 , \51401 );
xor \U$51455 ( \51798 , \51797 , \51406 );
or \U$51456 ( \51799 , \51793 , \51795 );
and \U$51457 ( \51800 , \51798 , \51799 );
nor \U$51458 ( \51801 , \51796 , \51800 );
and \U$51459 ( \51802 , \51789 , \51801 );
and \U$51460 ( \51803 , \51778 , \51788 );
or \U$51461 ( \51804 , \51802 , \51803 );
and \U$51462 ( \51805 , \51422 , \51804 );
and \U$51463 ( \51806 , \51415 , \51421 );
or \U$51464 ( \51807 , \51805 , \51806 );
not \U$51465 ( \51808 , \51807 );
xor \U$51466 ( \51809 , \50583 , \51016 );
xor \U$51467 ( \51810 , \51809 , \51021 );
xor \U$51468 ( \51811 , \50186 , \50511 );
xor \U$51469 ( \51812 , \51811 , \50536 );
xor \U$51470 ( \51813 , \51810 , \51812 );
not \U$51471 ( \51814 , \51378 );
or \U$51472 ( \51815 , \51409 , \51814 );
and \U$51473 ( \51816 , \51409 , \51814 );
nor \U$51474 ( \51817 , \51816 , \51363 );
not \U$51475 ( \51818 , \51817 );
nand \U$51476 ( \51819 , \51815 , \51818 );
xor \U$51477 ( \51820 , \50474 , \50490 );
xor \U$51478 ( \51821 , \51820 , \50505 );
and \U$51479 ( \51822 , \51048 , \51821 );
xor \U$51480 ( \51823 , \50474 , \50490 );
xor \U$51481 ( \51824 , \51823 , \50505 );
and \U$51482 ( \51825 , \51052 , \51824 );
and \U$51483 ( \51826 , \51048 , \51052 );
or \U$51484 ( \51827 , \51822 , \51825 , \51826 );
xor \U$51485 ( \51828 , \51819 , \51827 );
xor \U$51486 ( \51829 , \50526 , \50528 );
xor \U$51487 ( \51830 , \51829 , \50533 );
xor \U$51488 ( \51831 , \50571 , \50578 );
xor \U$51489 ( \51832 , \51830 , \51831 );
and \U$51490 ( \51833 , \51828 , \51832 );
and \U$51491 ( \51834 , \51819 , \51827 );
or \U$51492 ( \51835 , \51833 , \51834 );
xor \U$51493 ( \51836 , \51813 , \51835 );
nand \U$51494 ( \51837 , \51808 , \51836 );
xor \U$51495 ( \51838 , \50163 , \50165 );
xor \U$51496 ( \51839 , \51838 , \50168 );
xor \U$51497 ( \51840 , \51024 , \51029 );
xor \U$51498 ( \51841 , \51839 , \51840 );
not \U$51499 ( \51842 , \51841 );
xor \U$51500 ( \51843 , \51810 , \51812 );
and \U$51501 ( \51844 , \51843 , \51835 );
and \U$51502 ( \51845 , \51810 , \51812 );
nor \U$51503 ( \51846 , \51844 , \51845 );
not \U$51504 ( \51847 , \51846 );
and \U$51505 ( \51848 , \51842 , \51847 );
and \U$51506 ( \51849 , \51841 , \51846 );
nor \U$51507 ( \51850 , \51848 , \51849 );
xor \U$51508 ( \51851 , \51837 , \51850 );
xor \U$51509 ( \51852 , \51415 , \51421 );
xor \U$51510 ( \51853 , \51852 , \51804 );
xor \U$51511 ( \51854 , \51819 , \51827 );
xor \U$51512 ( \51855 , \51854 , \51832 );
not \U$51513 ( \51856 , \51855 );
or \U$51514 ( \51857 , \51853 , \51856 );
not \U$51515 ( \51858 , \51856 );
not \U$51516 ( \51859 , \51853 );
or \U$51517 ( \51860 , \51858 , \51859 );
not \U$51518 ( \51861 , \51054 );
not \U$51519 ( \51862 , \51413 );
not \U$51520 ( \51863 , \51056 );
and \U$51521 ( \51864 , \51862 , \51863 );
and \U$51522 ( \51865 , \51413 , \51056 );
nor \U$51523 ( \51866 , \51864 , \51865 );
not \U$51524 ( \51867 , \51866 );
or \U$51525 ( \51868 , \51861 , \51867 );
or \U$51526 ( \51869 , \51866 , \51054 );
nand \U$51527 ( \51870 , \51868 , \51869 );
not \U$51528 ( \51871 , \51870 );
xor \U$51529 ( \51872 , \51778 , \51788 );
xor \U$51530 ( \51873 , \51872 , \51801 );
or \U$51531 ( \51874 , \51871 , \51873 );
not \U$51532 ( \51875 , \51873 );
not \U$51533 ( \51876 , \51871 );
or \U$51534 ( \51877 , \51875 , \51876 );
xor \U$51535 ( \51878 , \51498 , \51742 );
xor \U$51536 ( \51879 , \51878 , \51757 );
xor \U$51537 ( \51880 , \51436 , \51438 );
xor \U$51538 ( \51881 , \51880 , \51443 );
and \U$51539 ( \51882 , \51879 , \51881 );
xor \U$51540 ( \51883 , \51072 , \51082 );
xor \U$51541 ( \51884 , \51883 , \51095 );
xor \U$51542 ( \51885 , \51763 , \51770 );
xor \U$51543 ( \51886 , \51884 , \51885 );
xor \U$51544 ( \51887 , \51436 , \51438 );
xor \U$51545 ( \51888 , \51887 , \51443 );
and \U$51546 ( \51889 , \51886 , \51888 );
and \U$51547 ( \51890 , \51879 , \51886 );
or \U$51548 ( \51891 , \51882 , \51889 , \51890 );
xor \U$51549 ( \51892 , \51526 , \51553 );
xor \U$51550 ( \51893 , \51892 , \51580 );
not \U$51551 ( \51894 , \51737 );
not \U$51552 ( \51895 , \51682 );
or \U$51553 ( \51896 , \51894 , \51895 );
or \U$51554 ( \51897 , \51682 , \51737 );
nand \U$51555 ( \51898 , \51896 , \51897 );
not \U$51556 ( \51899 , \51898 );
not \U$51557 ( \51900 , \51707 );
and \U$51558 ( \51901 , \51899 , \51900 );
and \U$51559 ( \51902 , \51898 , \51707 );
nor \U$51560 ( \51903 , \51901 , \51902 );
xor \U$51561 ( \51904 , \51893 , \51903 );
not \U$51562 ( \51905 , \51468 );
not \U$51563 ( \51906 , \51474 );
or \U$51564 ( \51907 , \51905 , \51906 );
or \U$51565 ( \51908 , \51474 , \51468 );
nand \U$51566 ( \51909 , \51907 , \51908 );
not \U$51567 ( \51910 , \51909 );
not \U$51568 ( \51911 , \51460 );
and \U$51569 ( \51912 , \51910 , \51911 );
and \U$51570 ( \51913 , \51909 , \51460 );
nor \U$51571 ( \51914 , \51912 , \51913 );
and \U$51572 ( \51915 , \51904 , \51914 );
and \U$51573 ( \51916 , \51893 , \51903 );
nor \U$51574 ( \51917 , \51915 , \51916 );
xor \U$51575 ( \51918 , \51207 , \51233 );
xor \U$51576 ( \51919 , \51918 , \51259 );
xor \U$51577 ( \51920 , \51917 , \51919 );
xor \U$51578 ( \51921 , \51288 , \51315 );
xor \U$51579 ( \51922 , \51921 , \51341 );
xor \U$51580 ( \51923 , \51424 , \51431 );
xor \U$51581 ( \51924 , \51922 , \51923 );
and \U$51582 ( \51925 , \51920 , \51924 );
and \U$51583 ( \51926 , \51917 , \51919 );
or \U$51584 ( \51927 , \51925 , \51926 );
nand \U$51585 ( \51928 , RI9870498_86, \463 );
not \U$51586 ( \51929 , \51928 );
not \U$51587 ( \51930 , \454 );
or \U$51588 ( \51931 , \51929 , \51930 );
or \U$51589 ( \51932 , \454 , \51928 );
nand \U$51590 ( \51933 , \51931 , \51932 );
and \U$51591 ( \51934 , \438 , RI9870588_88);
and \U$51592 ( \51935 , RI98703a8_84, \436 );
nor \U$51593 ( \51936 , \51934 , \51935 );
and \U$51594 ( \51937 , \51936 , \444 );
not \U$51595 ( \51938 , \51936 );
and \U$51596 ( \51939 , \51938 , \443 );
nor \U$51597 ( \51940 , \51937 , \51939 );
xor \U$51598 ( \51941 , \51933 , \51940 );
not \U$51599 ( \51942 , \51505 );
xor \U$51600 ( \51943 , \51524 , \51513 );
not \U$51601 ( \51944 , \51943 );
or \U$51602 ( \51945 , \51942 , \51944 );
or \U$51603 ( \51946 , \51943 , \51505 );
nand \U$51604 ( \51947 , \51945 , \51946 );
and \U$51605 ( \51948 , \51941 , \51947 );
and \U$51606 ( \51949 , \51933 , \51940 );
nor \U$51607 ( \51950 , \51948 , \51949 );
xor \U$51608 ( \51951 , \51561 , \51569 );
xor \U$51609 ( \51952 , \51951 , \51577 );
not \U$51610 ( \51953 , \51952 );
xor \U$51611 ( \51954 , \51719 , \51726 );
xor \U$51612 ( \51955 , \51954 , \51734 );
not \U$51613 ( \51956 , \51955 );
and \U$51614 ( \51957 , \51953 , \51956 );
and \U$51615 ( \51958 , \51955 , \51952 );
xor \U$51616 ( \51959 , \51534 , \51541 );
xor \U$51617 ( \51960 , \51959 , \51550 );
nor \U$51618 ( \51961 , \51958 , \51960 );
nor \U$51619 ( \51962 , \51957 , \51961 );
xor \U$51620 ( \51963 , \51950 , \51962 );
xor \U$51621 ( \51964 , \51689 , \51696 );
xor \U$51622 ( \51965 , \51964 , \51704 );
not \U$51623 ( \51966 , \51965 );
xor \U$51624 ( \51967 , \51590 , \51597 );
xor \U$51625 ( \51968 , \51967 , \51605 );
not \U$51626 ( \51969 , \51968 );
and \U$51627 ( \51970 , \51966 , \51969 );
and \U$51628 ( \51971 , \51968 , \51965 );
xor \U$51629 ( \51972 , \51664 , \51671 );
xor \U$51630 ( \51973 , \51972 , \51679 );
nor \U$51631 ( \51974 , \51971 , \51973 );
nor \U$51632 ( \51975 , \51970 , \51974 );
and \U$51633 ( \51976 , \51963 , \51975 );
and \U$51634 ( \51977 , \51950 , \51962 );
nor \U$51635 ( \51978 , \51976 , \51977 );
and \U$51636 ( \51979 , \13882 , RI986f868_60);
and \U$51637 ( \51980 , RI986f778_58, \13880 );
nor \U$51638 ( \51981 , \51979 , \51980 );
and \U$51639 ( \51982 , \51981 , \13359 );
not \U$51640 ( \51983 , \51981 );
and \U$51641 ( \51984 , \51983 , \13358 );
nor \U$51642 ( \51985 , \51982 , \51984 );
and \U$51643 ( \51986 , \15780 , RI986f4a8_52);
and \U$51644 ( \51987 , RI986f3b8_50, RI9873648_192);
nor \U$51645 ( \51988 , \51986 , \51987 );
not \U$51646 ( \51989 , \51988 );
not \U$51647 ( \51990 , RI9873558_190);
and \U$51648 ( \51991 , \51989 , \51990 );
and \U$51649 ( \51992 , \51988 , RI9873558_190);
nor \U$51650 ( \51993 , \51991 , \51992 );
xor \U$51651 ( \51994 , \51985 , \51993 );
and \U$51652 ( \51995 , \14937 , RI986fa48_64);
and \U$51653 ( \51996 , RI986f958_62, \14935 );
nor \U$51654 ( \51997 , \51995 , \51996 );
and \U$51655 ( \51998 , \51997 , \14538 );
not \U$51656 ( \51999 , \51997 );
and \U$51657 ( \52000 , \51999 , \14539 );
nor \U$51658 ( \52001 , \51998 , \52000 );
and \U$51659 ( \52002 , \51994 , \52001 );
and \U$51660 ( \52003 , \51985 , \51993 );
or \U$51661 ( \52004 , \52002 , \52003 );
not \U$51662 ( \52005 , \52004 );
and \U$51663 ( \52006 , \11696 , RI986f2c8_48);
and \U$51664 ( \52007 , RI986f1d8_46, \11694 );
nor \U$51665 ( \52008 , \52006 , \52007 );
and \U$51666 ( \52009 , \52008 , \11702 );
not \U$51667 ( \52010 , \52008 );
and \U$51668 ( \52011 , \52010 , \10965 );
nor \U$51669 ( \52012 , \52009 , \52011 );
and \U$51670 ( \52013 , \12293 , RI986e5a8_20);
and \U$51671 ( \52014 , RI986e4b8_18, \12291 );
nor \U$51672 ( \52015 , \52013 , \52014 );
and \U$51673 ( \52016 , \52015 , \11686 );
not \U$51674 ( \52017 , \52015 );
and \U$51675 ( \52018 , \52017 , \11687 );
nor \U$51676 ( \52019 , \52016 , \52018 );
xor \U$51677 ( \52020 , \52012 , \52019 );
and \U$51678 ( \52021 , \13045 , RI986e788_24);
and \U$51679 ( \52022 , RI986e698_22, \13043 );
nor \U$51680 ( \52023 , \52021 , \52022 );
and \U$51681 ( \52024 , \52023 , \12619 );
not \U$51682 ( \52025 , \52023 );
and \U$51683 ( \52026 , \52025 , \13047 );
nor \U$51684 ( \52027 , \52024 , \52026 );
and \U$51685 ( \52028 , \52020 , \52027 );
and \U$51686 ( \52029 , \52012 , \52019 );
or \U$51687 ( \52030 , \52028 , \52029 );
not \U$51688 ( \52031 , \52030 );
and \U$51689 ( \52032 , \52005 , \52031 );
and \U$51690 ( \52033 , \52030 , \52004 );
and \U$51691 ( \52034 , \9505 , RI986ec38_34);
and \U$51692 ( \52035 , RI986ed28_36, \9503 );
nor \U$51693 ( \52036 , \52034 , \52035 );
and \U$51694 ( \52037 , \52036 , \9513 );
not \U$51695 ( \52038 , \52036 );
and \U$51696 ( \52039 , \52038 , \9510 );
nor \U$51697 ( \52040 , \52037 , \52039 );
and \U$51698 ( \52041 , \9237 , RI986ef08_40);
and \U$51699 ( \52042 , RI986ee18_38, \9235 );
nor \U$51700 ( \52043 , \52041 , \52042 );
and \U$51701 ( \52044 , \52043 , \8836 );
not \U$51702 ( \52045 , \52043 );
and \U$51703 ( \52046 , \52045 , \9241 );
nor \U$51704 ( \52047 , \52044 , \52046 );
xor \U$51705 ( \52048 , \52040 , \52047 );
and \U$51706 ( \52049 , \10424 , RI986f0e8_44);
and \U$51707 ( \52050 , RI986eff8_42, \10422 );
nor \U$51708 ( \52051 , \52049 , \52050 );
and \U$51709 ( \52052 , \52051 , \10428 );
not \U$51710 ( \52053 , \52051 );
and \U$51711 ( \52054 , \52053 , \9840 );
nor \U$51712 ( \52055 , \52052 , \52054 );
and \U$51713 ( \52056 , \52048 , \52055 );
and \U$51714 ( \52057 , \52040 , \52047 );
or \U$51715 ( \52058 , \52056 , \52057 );
nor \U$51716 ( \52059 , \52033 , \52058 );
nor \U$51717 ( \52060 , \52032 , \52059 );
and \U$51718 ( \52061 , \5881 , RI9871398_118);
and \U$51719 ( \52062 , RI9871488_120, \5879 );
nor \U$51720 ( \52063 , \52061 , \52062 );
and \U$51721 ( \52064 , \52063 , \5885 );
not \U$51722 ( \52065 , \52063 );
and \U$51723 ( \52066 , \52065 , \5594 );
nor \U$51724 ( \52067 , \52064 , \52066 );
and \U$51725 ( \52068 , \6453 , RI9871758_126);
and \U$51726 ( \52069 , RI9871848_128, \6451 );
nor \U$51727 ( \52070 , \52068 , \52069 );
and \U$51728 ( \52071 , \52070 , \6180 );
not \U$51729 ( \52072 , \52070 );
and \U$51730 ( \52073 , \52072 , \6190 );
nor \U$51731 ( \52074 , \52071 , \52073 );
xor \U$51732 ( \52075 , \52067 , \52074 );
and \U$51733 ( \52076 , \5318 , RI98712a8_116);
and \U$51734 ( \52077 , RI98711b8_114, \5316 );
nor \U$51735 ( \52078 , \52076 , \52077 );
and \U$51736 ( \52079 , \52078 , \5322 );
not \U$51737 ( \52080 , \52078 );
and \U$51738 ( \52081 , \52080 , \5052 );
nor \U$51739 ( \52082 , \52079 , \52081 );
and \U$51740 ( \52083 , \52075 , \52082 );
and \U$51741 ( \52084 , \52067 , \52074 );
nor \U$51742 ( \52085 , \52083 , \52084 );
and \U$51743 ( \52086 , \4203 , RI9870ee8_108);
and \U$51744 ( \52087 , RI9870c18_102, \4201 );
nor \U$51745 ( \52088 , \52086 , \52087 );
and \U$51746 ( \52089 , \52088 , \3922 );
not \U$51747 ( \52090 , \52088 );
and \U$51748 ( \52091 , \52090 , \4207 );
nor \U$51749 ( \52092 , \52089 , \52091 );
and \U$51750 ( \52093 , \4710 , RI98710c8_112);
and \U$51751 ( \52094 , RI9870d08_104, \4708 );
nor \U$51752 ( \52095 , \52093 , \52094 );
not \U$51753 ( \52096 , \52095 );
not \U$51754 ( \52097 , \4519 );
and \U$51755 ( \52098 , \52096 , \52097 );
and \U$51756 ( \52099 , \52095 , \4519 );
nor \U$51757 ( \52100 , \52098 , \52099 );
xor \U$51758 ( \52101 , \52092 , \52100 );
and \U$51759 ( \52102 , \3683 , RI9870df8_106);
and \U$51760 ( \52103 , RI9870a38_98, \3681 );
nor \U$51761 ( \52104 , \52102 , \52103 );
not \U$51762 ( \52105 , \52104 );
not \U$51763 ( \52106 , \3918 );
and \U$51764 ( \52107 , \52105 , \52106 );
and \U$51765 ( \52108 , \52104 , \3918 );
nor \U$51766 ( \52109 , \52107 , \52108 );
and \U$51767 ( \52110 , \52101 , \52109 );
and \U$51768 ( \52111 , \52092 , \52100 );
nor \U$51769 ( \52112 , \52110 , \52111 );
xor \U$51770 ( \52113 , \52085 , \52112 );
and \U$51771 ( \52114 , \7729 , RI986eb48_32);
and \U$51772 ( \52115 , RI986ea58_30, \7727 );
nor \U$51773 ( \52116 , \52114 , \52115 );
and \U$51774 ( \52117 , \52116 , \7733 );
not \U$51775 ( \52118 , \52116 );
and \U$51776 ( \52119 , \52118 , \7480 );
nor \U$51777 ( \52120 , \52117 , \52119 );
and \U$51778 ( \52121 , \8486 , RI986e968_28);
and \U$51779 ( \52122 , RI986e878_26, \8484 );
nor \U$51780 ( \52123 , \52121 , \52122 );
and \U$51781 ( \52124 , \52123 , \8051 );
not \U$51782 ( \52125 , \52123 );
and \U$51783 ( \52126 , \52125 , \8050 );
nor \U$51784 ( \52127 , \52124 , \52126 );
xor \U$51785 ( \52128 , \52120 , \52127 );
and \U$51786 ( \52129 , \7079 , RI9871578_122);
and \U$51787 ( \52130 , RI9871668_124, \7077 );
nor \U$51788 ( \52131 , \52129 , \52130 );
and \U$51789 ( \52132 , \52131 , \6709 );
not \U$51790 ( \52133 , \52131 );
and \U$51791 ( \52134 , \52133 , \6710 );
nor \U$51792 ( \52135 , \52132 , \52134 );
and \U$51793 ( \52136 , \52128 , \52135 );
and \U$51794 ( \52137 , \52120 , \52127 );
nor \U$51795 ( \52138 , \52136 , \52137 );
and \U$51796 ( \52139 , \52113 , \52138 );
and \U$51797 ( \52140 , \52085 , \52112 );
nor \U$51798 ( \52141 , \52139 , \52140 );
or \U$51799 ( \52142 , \52060 , \52141 );
not \U$51800 ( \52143 , \52060 );
not \U$51801 ( \52144 , \52141 );
or \U$51802 ( \52145 , \52143 , \52144 );
and \U$51803 ( \52146 , \2464 , RI98700d8_78);
and \U$51804 ( \52147 , RI98701c8_80, \2462 );
nor \U$51805 ( \52148 , \52146 , \52147 );
and \U$51806 ( \52149 , \52148 , \2263 );
not \U$51807 ( \52150 , \52148 );
and \U$51808 ( \52151 , \52150 , \2468 );
nor \U$51809 ( \52152 , \52149 , \52151 );
and \U$51810 ( \52153 , \3254 , RI9870fd8_110);
and \U$51811 ( \52154 , RI9870b28_100, \3252 );
nor \U$51812 ( \52155 , \52153 , \52154 );
not \U$51813 ( \52156 , \52155 );
not \U$51814 ( \52157 , \3406 );
and \U$51815 ( \52158 , \52156 , \52157 );
and \U$51816 ( \52159 , \52155 , \2935 );
nor \U$51817 ( \52160 , \52158 , \52159 );
xor \U$51818 ( \52161 , \52152 , \52160 );
and \U$51819 ( \52162 , \2274 , RI986ffe8_76);
and \U$51820 ( \52163 , RI986fef8_74, \2272 );
nor \U$51821 ( \52164 , \52162 , \52163 );
and \U$51822 ( \52165 , \52164 , \2031 );
not \U$51823 ( \52166 , \52164 );
and \U$51824 ( \52167 , \52166 , \2030 );
nor \U$51825 ( \52168 , \52165 , \52167 );
and \U$51826 ( \52169 , \52161 , \52168 );
and \U$51827 ( \52170 , \52152 , \52160 );
nor \U$51828 ( \52171 , \52169 , \52170 );
and \U$51829 ( \52172 , \438 , RI9870498_86);
and \U$51830 ( \52173 , RI9870588_88, \436 );
nor \U$51831 ( \52174 , \52172 , \52173 );
and \U$51832 ( \52175 , \52174 , \444 );
not \U$51833 ( \52176 , \52174 );
and \U$51834 ( \52177 , \52176 , \443 );
nor \U$51835 ( \52178 , \52175 , \52177 );
and \U$51836 ( \52179 , \776 , RI98703a8_84);
and \U$51837 ( \52180 , RI98702b8_82, \774 );
nor \U$51838 ( \52181 , \52179 , \52180 );
and \U$51839 ( \52182 , \52181 , \474 );
not \U$51840 ( \52183 , \52181 );
and \U$51841 ( \52184 , \52183 , \451 );
nor \U$51842 ( \52185 , \52182 , \52184 );
xor \U$51843 ( \52186 , \52178 , \52185 );
not \U$51844 ( \52187 , \1301 );
and \U$51845 ( \52188 , \1293 , RI9870768_92);
and \U$51846 ( \52189 , RI9870678_90, \1291 );
nor \U$51847 ( \52190 , \52188 , \52189 );
not \U$51848 ( \52191 , \52190 );
or \U$51849 ( \52192 , \52187 , \52191 );
or \U$51850 ( \52193 , \52190 , \1301 );
nand \U$51851 ( \52194 , \52192 , \52193 );
and \U$51852 ( \52195 , \52186 , \52194 );
and \U$51853 ( \52196 , \52178 , \52185 );
or \U$51854 ( \52197 , \52195 , \52196 );
xor \U$51855 ( \52198 , \52171 , \52197 );
and \U$51856 ( \52199 , \1329 , RI9870948_96);
and \U$51857 ( \52200 , RI9870858_94, \1327 );
nor \U$51858 ( \52201 , \52199 , \52200 );
and \U$51859 ( \52202 , \52201 , \1337 );
not \U$51860 ( \52203 , \52201 );
and \U$51861 ( \52204 , \52203 , \1336 );
nor \U$51862 ( \52205 , \52202 , \52204 );
and \U$51863 ( \52206 , \2042 , RI986fe08_72);
and \U$51864 ( \52207 , RI986fd18_70, \2040 );
nor \U$51865 ( \52208 , \52206 , \52207 );
not \U$51866 ( \52209 , \52208 );
not \U$51867 ( \52210 , \1462 );
and \U$51868 ( \52211 , \52209 , \52210 );
and \U$51869 ( \52212 , \52208 , \1462 );
nor \U$51870 ( \52213 , \52211 , \52212 );
or \U$51871 ( \52214 , \52205 , \52213 );
not \U$51872 ( \52215 , \52213 );
not \U$51873 ( \52216 , \52205 );
or \U$51874 ( \52217 , \52215 , \52216 );
and \U$51875 ( \52218 , \1311 , RI986fb38_66);
and \U$51876 ( \52219 , RI986fc28_68, \1309 );
nor \U$51877 ( \52220 , \52218 , \52219 );
and \U$51878 ( \52221 , \52220 , \1458 );
not \U$51879 ( \52222 , \52220 );
and \U$51880 ( \52223 , \52222 , \1318 );
nor \U$51881 ( \52224 , \52221 , \52223 );
nand \U$51882 ( \52225 , \52217 , \52224 );
nand \U$51883 ( \52226 , \52214 , \52225 );
and \U$51884 ( \52227 , \52198 , \52226 );
and \U$51885 ( \52228 , \52171 , \52197 );
or \U$51886 ( \52229 , \52227 , \52228 );
nand \U$51887 ( \52230 , \52145 , \52229 );
nand \U$51888 ( \52231 , \52142 , \52230 );
xor \U$51889 ( \52232 , \51978 , \52231 );
xor \U$51890 ( \52233 , \51479 , \51489 );
xor \U$51891 ( \52234 , \52233 , \51492 );
xor \U$51892 ( \52235 , \51215 , \51222 );
xor \U$51893 ( \52236 , \52235 , \51230 );
or \U$51894 ( \52237 , \52234 , \52236 );
not \U$51895 ( \52238 , \52236 );
not \U$51896 ( \52239 , \52234 );
or \U$51897 ( \52240 , \52238 , \52239 );
xor \U$51898 ( \52241 , \51323 , \51330 );
xor \U$51899 ( \52242 , \52241 , \51338 );
xor \U$51900 ( \52243 , \51448 , \51453 );
xor \U$51901 ( \52244 , \52242 , \52243 );
nand \U$51902 ( \52245 , \52240 , \52244 );
nand \U$51903 ( \52246 , \52237 , \52245 );
and \U$51904 ( \52247 , \52232 , \52246 );
and \U$51905 ( \52248 , \51978 , \52231 );
or \U$51906 ( \52249 , \52247 , \52248 );
xor \U$51907 ( \52250 , \51927 , \52249 );
xor \U$51908 ( \52251 , \51583 , \51656 );
xor \U$51909 ( \52252 , \52251 , \51739 );
xor \U$51910 ( \52253 , \51458 , \51476 );
xor \U$51911 ( \52254 , \52253 , \51495 );
and \U$51912 ( \52255 , \52252 , \52254 );
xor \U$51913 ( \52256 , \51074 , \51076 );
xor \U$51914 ( \52257 , \52256 , \51079 );
xor \U$51915 ( \52258 , \51745 , \51752 );
xor \U$51916 ( \52259 , \52257 , \52258 );
xor \U$51917 ( \52260 , \51458 , \51476 );
xor \U$51918 ( \52261 , \52260 , \51495 );
and \U$51919 ( \52262 , \52259 , \52261 );
and \U$51920 ( \52263 , \52252 , \52259 );
or \U$51921 ( \52264 , \52255 , \52262 , \52263 );
and \U$51922 ( \52265 , \52250 , \52264 );
and \U$51923 ( \52266 , \51927 , \52249 );
or \U$51924 ( \52267 , \52265 , \52266 );
xor \U$51925 ( \52268 , \51891 , \52267 );
not \U$51926 ( \52269 , \51798 );
xnor \U$51927 ( \52270 , \51795 , \51793 );
not \U$51928 ( \52271 , \52270 );
or \U$51929 ( \52272 , \52269 , \52271 );
or \U$51930 ( \52273 , \52270 , \51798 );
nand \U$51931 ( \52274 , \52272 , \52273 );
and \U$51932 ( \52275 , \52268 , \52274 );
and \U$51933 ( \52276 , \51891 , \52267 );
or \U$51934 ( \52277 , \52275 , \52276 );
nand \U$51935 ( \52278 , \51877 , \52277 );
nand \U$51936 ( \52279 , \51874 , \52278 );
nand \U$51937 ( \52280 , \51860 , \52279 );
nand \U$51938 ( \52281 , \51857 , \52280 );
not \U$51939 ( \52282 , \51807 );
not \U$51940 ( \52283 , \51836 );
or \U$51941 ( \52284 , \52282 , \52283 );
or \U$51942 ( \52285 , \51836 , \51807 );
nand \U$51943 ( \52286 , \52284 , \52285 );
and \U$51944 ( \52287 , \52281 , \52286 );
xor \U$51945 ( \52288 , \52286 , \52281 );
not \U$51946 ( \52289 , \51853 );
not \U$51947 ( \52290 , \52279 );
and \U$51948 ( \52291 , \52289 , \52290 );
and \U$51949 ( \52292 , \52279 , \51853 );
nor \U$51950 ( \52293 , \52291 , \52292 );
not \U$51951 ( \52294 , \52293 );
not \U$51952 ( \52295 , \51855 );
and \U$51953 ( \52296 , \52294 , \52295 );
and \U$51954 ( \52297 , \52293 , \51855 );
nor \U$51955 ( \52298 , \52296 , \52297 );
not \U$51956 ( \52299 , \51873 );
not \U$51957 ( \52300 , \52277 );
and \U$51958 ( \52301 , \52299 , \52300 );
and \U$51959 ( \52302 , \51873 , \52277 );
nor \U$51960 ( \52303 , \52301 , \52302 );
not \U$51961 ( \52304 , \52303 );
not \U$51962 ( \52305 , \51870 );
and \U$51963 ( \52306 , \52304 , \52305 );
and \U$51964 ( \52307 , \52303 , \51870 );
nor \U$51965 ( \52308 , \52306 , \52307 );
not \U$51966 ( \52309 , \52308 );
xor \U$51967 ( \52310 , \51978 , \52231 );
xor \U$51968 ( \52311 , \52310 , \52246 );
xor \U$51969 ( \52312 , \51917 , \51919 );
xor \U$51970 ( \52313 , \52312 , \51924 );
and \U$51971 ( \52314 , \52311 , \52313 );
xor \U$51972 ( \52315 , \51458 , \51476 );
xor \U$51973 ( \52316 , \52315 , \51495 );
xor \U$51974 ( \52317 , \52252 , \52259 );
xor \U$51975 ( \52318 , \52316 , \52317 );
xor \U$51976 ( \52319 , \51917 , \51919 );
xor \U$51977 ( \52320 , \52319 , \51924 );
and \U$51978 ( \52321 , \52318 , \52320 );
and \U$51979 ( \52322 , \52311 , \52318 );
or \U$51980 ( \52323 , \52314 , \52321 , \52322 );
xor \U$51981 ( \52324 , \51616 , \456 );
xor \U$51982 ( \52325 , \52324 , \51624 );
xor \U$51983 ( \52326 , \51635 , \51642 );
xor \U$51984 ( \52327 , \52326 , \51650 );
and \U$51985 ( \52328 , \52325 , \52327 );
not \U$51986 ( \52329 , \51965 );
xor \U$51987 ( \52330 , \51973 , \51968 );
not \U$51988 ( \52331 , \52330 );
or \U$51989 ( \52332 , \52329 , \52331 );
or \U$51990 ( \52333 , \52330 , \51965 );
nand \U$51991 ( \52334 , \52332 , \52333 );
xor \U$51992 ( \52335 , \51635 , \51642 );
xor \U$51993 ( \52336 , \52335 , \51650 );
and \U$51994 ( \52337 , \52334 , \52336 );
and \U$51995 ( \52338 , \52325 , \52334 );
or \U$51996 ( \52339 , \52328 , \52337 , \52338 );
and \U$51997 ( \52340 , \776 , RI9870588_88);
and \U$51998 ( \52341 , RI98703a8_84, \774 );
nor \U$51999 ( \52342 , \52340 , \52341 );
and \U$52000 ( \52343 , \52342 , \451 );
not \U$52001 ( \52344 , \52342 );
and \U$52002 ( \52345 , \52344 , \474 );
nor \U$52003 ( \52346 , \52343 , \52345 );
not \U$52004 ( \52347 , \52346 );
and \U$52005 ( \52348 , \1329 , RI9870678_90);
and \U$52006 ( \52349 , RI9870948_96, \1327 );
nor \U$52007 ( \52350 , \52348 , \52349 );
and \U$52008 ( \52351 , \52350 , \1337 );
not \U$52009 ( \52352 , \52350 );
and \U$52010 ( \52353 , \52352 , \1336 );
nor \U$52011 ( \52354 , \52351 , \52353 );
not \U$52012 ( \52355 , \52354 );
and \U$52013 ( \52356 , \52347 , \52355 );
and \U$52014 ( \52357 , \52354 , \52346 );
and \U$52015 ( \52358 , \1293 , RI98702b8_82);
and \U$52016 ( \52359 , RI9870768_92, \1291 );
nor \U$52017 ( \52360 , \52358 , \52359 );
not \U$52018 ( \52361 , \52360 );
not \U$52019 ( \52362 , \1301 );
and \U$52020 ( \52363 , \52361 , \52362 );
and \U$52021 ( \52364 , \52360 , \1128 );
nor \U$52022 ( \52365 , \52363 , \52364 );
nor \U$52023 ( \52366 , \52357 , \52365 );
nor \U$52024 ( \52367 , \52356 , \52366 );
and \U$52025 ( \52368 , \1311 , RI9870858_94);
and \U$52026 ( \52369 , RI986fb38_66, \1309 );
nor \U$52027 ( \52370 , \52368 , \52369 );
and \U$52028 ( \52371 , \52370 , \1315 );
not \U$52029 ( \52372 , \52370 );
and \U$52030 ( \52373 , \52372 , \1458 );
nor \U$52031 ( \52374 , \52371 , \52373 );
not \U$52032 ( \52375 , \52374 );
and \U$52033 ( \52376 , \2274 , RI986fd18_70);
and \U$52034 ( \52377 , RI986ffe8_76, \2272 );
nor \U$52035 ( \52378 , \52376 , \52377 );
and \U$52036 ( \52379 , \52378 , \2031 );
not \U$52037 ( \52380 , \52378 );
and \U$52038 ( \52381 , \52380 , \2030 );
nor \U$52039 ( \52382 , \52379 , \52381 );
not \U$52040 ( \52383 , \52382 );
and \U$52041 ( \52384 , \52375 , \52383 );
and \U$52042 ( \52385 , \52382 , \52374 );
and \U$52043 ( \52386 , \2042 , RI986fc28_68);
and \U$52044 ( \52387 , RI986fe08_72, \2040 );
nor \U$52045 ( \52388 , \52386 , \52387 );
not \U$52046 ( \52389 , \52388 );
not \U$52047 ( \52390 , \2034 );
and \U$52048 ( \52391 , \52389 , \52390 );
and \U$52049 ( \52392 , \52388 , \1462 );
nor \U$52050 ( \52393 , \52391 , \52392 );
nor \U$52051 ( \52394 , \52385 , \52393 );
nor \U$52052 ( \52395 , \52384 , \52394 );
or \U$52053 ( \52396 , \52367 , \52395 );
not \U$52054 ( \52397 , \52367 );
not \U$52055 ( \52398 , \52395 );
or \U$52056 ( \52399 , \52397 , \52398 );
and \U$52057 ( \52400 , \3254 , RI98701c8_80);
and \U$52058 ( \52401 , RI9870fd8_110, \3252 );
nor \U$52059 ( \52402 , \52400 , \52401 );
not \U$52060 ( \52403 , \52402 );
not \U$52061 ( \52404 , \3406 );
and \U$52062 ( \52405 , \52403 , \52404 );
and \U$52063 ( \52406 , \52402 , \2935 );
nor \U$52064 ( \52407 , \52405 , \52406 );
and \U$52065 ( \52408 , \3683 , RI9870b28_100);
and \U$52066 ( \52409 , RI9870df8_106, \3681 );
nor \U$52067 ( \52410 , \52408 , \52409 );
not \U$52068 ( \52411 , \52410 );
not \U$52069 ( \52412 , \3412 );
and \U$52070 ( \52413 , \52411 , \52412 );
and \U$52071 ( \52414 , \52410 , \3918 );
nor \U$52072 ( \52415 , \52413 , \52414 );
xor \U$52073 ( \52416 , \52407 , \52415 );
and \U$52074 ( \52417 , \2464 , RI986fef8_74);
and \U$52075 ( \52418 , RI98700d8_78, \2462 );
nor \U$52076 ( \52419 , \52417 , \52418 );
and \U$52077 ( \52420 , \52419 , \2263 );
not \U$52078 ( \52421 , \52419 );
and \U$52079 ( \52422 , \52421 , \2468 );
nor \U$52080 ( \52423 , \52420 , \52422 );
and \U$52081 ( \52424 , \52416 , \52423 );
and \U$52082 ( \52425 , \52407 , \52415 );
nor \U$52083 ( \52426 , \52424 , \52425 );
nand \U$52084 ( \52427 , \52399 , \52426 );
nand \U$52085 ( \52428 , \52396 , \52427 );
and \U$52086 ( \52429 , \15780 , RI986f958_62);
and \U$52087 ( \52430 , RI986f4a8_52, RI9873648_192);
nor \U$52088 ( \52431 , \52429 , \52430 );
not \U$52089 ( \52432 , \52431 );
not \U$52090 ( \52433 , RI9873558_190);
and \U$52091 ( \52434 , \52432 , \52433 );
and \U$52092 ( \52435 , \52431 , RI9873558_190);
nor \U$52093 ( \52436 , \52434 , \52435 );
not \U$52094 ( \52437 , \52436 );
not \U$52095 ( \52438 , \444 );
and \U$52096 ( \52439 , \52437 , \52438 );
and \U$52097 ( \52440 , \52436 , \444 );
and \U$52098 ( \52441 , \14937 , RI986f778_58);
and \U$52099 ( \52442 , RI986fa48_64, \14935 );
nor \U$52100 ( \52443 , \52441 , \52442 );
and \U$52101 ( \52444 , \52443 , \14538 );
not \U$52102 ( \52445 , \52443 );
and \U$52103 ( \52446 , \52445 , \14539 );
nor \U$52104 ( \52447 , \52444 , \52446 );
nor \U$52105 ( \52448 , \52440 , \52447 );
nor \U$52106 ( \52449 , \52439 , \52448 );
and \U$52107 ( \52450 , \12293 , RI986f1d8_46);
and \U$52108 ( \52451 , RI986e5a8_20, \12291 );
nor \U$52109 ( \52452 , \52450 , \52451 );
and \U$52110 ( \52453 , \52452 , \11686 );
not \U$52111 ( \52454 , \52452 );
and \U$52112 ( \52455 , \52454 , \11687 );
nor \U$52113 ( \52456 , \52453 , \52455 );
not \U$52114 ( \52457 , \52456 );
and \U$52115 ( \52458 , \13882 , RI986e698_22);
and \U$52116 ( \52459 , RI986f868_60, \13880 );
nor \U$52117 ( \52460 , \52458 , \52459 );
and \U$52118 ( \52461 , \52460 , \13359 );
not \U$52119 ( \52462 , \52460 );
and \U$52120 ( \52463 , \52462 , \13358 );
nor \U$52121 ( \52464 , \52461 , \52463 );
not \U$52122 ( \52465 , \52464 );
and \U$52123 ( \52466 , \52457 , \52465 );
and \U$52124 ( \52467 , \52464 , \52456 );
and \U$52125 ( \52468 , \13045 , RI986e4b8_18);
and \U$52126 ( \52469 , RI986e788_24, \13043 );
nor \U$52127 ( \52470 , \52468 , \52469 );
and \U$52128 ( \52471 , \52470 , \12619 );
not \U$52129 ( \52472 , \52470 );
and \U$52130 ( \52473 , \52472 , \13047 );
nor \U$52131 ( \52474 , \52471 , \52473 );
nor \U$52132 ( \52475 , \52467 , \52474 );
nor \U$52133 ( \52476 , \52466 , \52475 );
xor \U$52134 ( \52477 , \52449 , \52476 );
and \U$52135 ( \52478 , \9505 , RI986ee18_38);
and \U$52136 ( \52479 , RI986ec38_34, \9503 );
nor \U$52137 ( \52480 , \52478 , \52479 );
and \U$52138 ( \52481 , \52480 , \9513 );
not \U$52139 ( \52482 , \52480 );
and \U$52140 ( \52483 , \52482 , \9510 );
nor \U$52141 ( \52484 , \52481 , \52483 );
not \U$52142 ( \52485 , \52484 );
and \U$52143 ( \52486 , \11696 , RI986eff8_42);
and \U$52144 ( \52487 , RI986f2c8_48, \11694 );
nor \U$52145 ( \52488 , \52486 , \52487 );
and \U$52146 ( \52489 , \52488 , \11702 );
not \U$52147 ( \52490 , \52488 );
and \U$52148 ( \52491 , \52490 , \10965 );
nor \U$52149 ( \52492 , \52489 , \52491 );
not \U$52150 ( \52493 , \52492 );
and \U$52151 ( \52494 , \52485 , \52493 );
and \U$52152 ( \52495 , \52492 , \52484 );
and \U$52153 ( \52496 , \10424 , RI986ed28_36);
and \U$52154 ( \52497 , RI986f0e8_44, \10422 );
nor \U$52155 ( \52498 , \52496 , \52497 );
and \U$52156 ( \52499 , \52498 , \10428 );
not \U$52157 ( \52500 , \52498 );
and \U$52158 ( \52501 , \52500 , \9840 );
nor \U$52159 ( \52502 , \52499 , \52501 );
nor \U$52160 ( \52503 , \52495 , \52502 );
nor \U$52161 ( \52504 , \52494 , \52503 );
and \U$52162 ( \52505 , \52477 , \52504 );
and \U$52163 ( \52506 , \52449 , \52476 );
nor \U$52164 ( \52507 , \52505 , \52506 );
xor \U$52165 ( \52508 , \52428 , \52507 );
and \U$52166 ( \52509 , \5881 , RI98711b8_114);
and \U$52167 ( \52510 , RI9871398_118, \5879 );
nor \U$52168 ( \52511 , \52509 , \52510 );
and \U$52169 ( \52512 , \52511 , \5885 );
not \U$52170 ( \52513 , \52511 );
and \U$52171 ( \52514 , \52513 , \5594 );
nor \U$52172 ( \52515 , \52512 , \52514 );
and \U$52173 ( \52516 , \7079 , RI9871848_128);
and \U$52174 ( \52517 , RI9871578_122, \7077 );
nor \U$52175 ( \52518 , \52516 , \52517 );
and \U$52176 ( \52519 , \52518 , \6709 );
not \U$52177 ( \52520 , \52518 );
and \U$52178 ( \52521 , \52520 , \6710 );
nor \U$52179 ( \52522 , \52519 , \52521 );
or \U$52180 ( \52523 , \52515 , \52522 );
not \U$52181 ( \52524 , \52522 );
not \U$52182 ( \52525 , \52515 );
or \U$52183 ( \52526 , \52524 , \52525 );
and \U$52184 ( \52527 , \6453 , RI9871488_120);
and \U$52185 ( \52528 , RI9871758_126, \6451 );
nor \U$52186 ( \52529 , \52527 , \52528 );
and \U$52187 ( \52530 , \52529 , \6190 );
not \U$52188 ( \52531 , \52529 );
and \U$52189 ( \52532 , \52531 , \6705 );
nor \U$52190 ( \52533 , \52530 , \52532 );
nand \U$52191 ( \52534 , \52526 , \52533 );
nand \U$52192 ( \52535 , \52523 , \52534 );
and \U$52193 ( \52536 , \4710 , RI9870c18_102);
and \U$52194 ( \52537 , RI98710c8_112, \4708 );
nor \U$52195 ( \52538 , \52536 , \52537 );
not \U$52196 ( \52539 , \52538 );
not \U$52197 ( \52540 , \4521 );
and \U$52198 ( \52541 , \52539 , \52540 );
and \U$52199 ( \52542 , \52538 , \4519 );
nor \U$52200 ( \52543 , \52541 , \52542 );
and \U$52201 ( \52544 , \5318 , RI9870d08_104);
and \U$52202 ( \52545 , RI98712a8_116, \5316 );
nor \U$52203 ( \52546 , \52544 , \52545 );
and \U$52204 ( \52547 , \52546 , \5322 );
not \U$52205 ( \52548 , \52546 );
and \U$52206 ( \52549 , \52548 , \5052 );
nor \U$52207 ( \52550 , \52547 , \52549 );
xor \U$52208 ( \52551 , \52543 , \52550 );
and \U$52209 ( \52552 , \4203 , RI9870a38_98);
and \U$52210 ( \52553 , RI9870ee8_108, \4201 );
nor \U$52211 ( \52554 , \52552 , \52553 );
and \U$52212 ( \52555 , \52554 , \3923 );
not \U$52213 ( \52556 , \52554 );
and \U$52214 ( \52557 , \52556 , \4207 );
nor \U$52215 ( \52558 , \52555 , \52557 );
and \U$52216 ( \52559 , \52551 , \52558 );
and \U$52217 ( \52560 , \52543 , \52550 );
nor \U$52218 ( \52561 , \52559 , \52560 );
xor \U$52219 ( \52562 , \52535 , \52561 );
and \U$52220 ( \52563 , \8486 , RI986ea58_30);
and \U$52221 ( \52564 , RI986e968_28, \8484 );
nor \U$52222 ( \52565 , \52563 , \52564 );
and \U$52223 ( \52566 , \52565 , \8050 );
not \U$52224 ( \52567 , \52565 );
and \U$52225 ( \52568 , \52567 , \8051 );
nor \U$52226 ( \52569 , \52566 , \52568 );
and \U$52227 ( \52570 , \7729 , RI9871668_124);
and \U$52228 ( \52571 , RI986eb48_32, \7727 );
nor \U$52229 ( \52572 , \52570 , \52571 );
and \U$52230 ( \52573 , \52572 , \7480 );
not \U$52231 ( \52574 , \52572 );
and \U$52232 ( \52575 , \52574 , \7733 );
nor \U$52233 ( \52576 , \52573 , \52575 );
xor \U$52234 ( \52577 , \52569 , \52576 );
and \U$52235 ( \52578 , \9237 , RI986e878_26);
and \U$52236 ( \52579 , RI986ef08_40, \9235 );
nor \U$52237 ( \52580 , \52578 , \52579 );
and \U$52238 ( \52581 , \52580 , \9241 );
not \U$52239 ( \52582 , \52580 );
and \U$52240 ( \52583 , \52582 , \8836 );
nor \U$52241 ( \52584 , \52581 , \52583 );
and \U$52242 ( \52585 , \52577 , \52584 );
and \U$52243 ( \52586 , \52569 , \52576 );
or \U$52244 ( \52587 , \52585 , \52586 );
and \U$52245 ( \52588 , \52562 , \52587 );
and \U$52246 ( \52589 , \52535 , \52561 );
or \U$52247 ( \52590 , \52588 , \52589 );
and \U$52248 ( \52591 , \52508 , \52590 );
and \U$52249 ( \52592 , \52428 , \52507 );
or \U$52250 ( \52593 , \52591 , \52592 );
xor \U$52251 ( \52594 , \52339 , \52593 );
xor \U$52252 ( \52595 , \52092 , \52100 );
xor \U$52253 ( \52596 , \52595 , \52109 );
xor \U$52254 ( \52597 , \52067 , \52074 );
xor \U$52255 ( \52598 , \52597 , \52082 );
xor \U$52256 ( \52599 , \52596 , \52598 );
xor \U$52257 ( \52600 , \52120 , \52127 );
xor \U$52258 ( \52601 , \52600 , \52135 );
and \U$52259 ( \52602 , \52599 , \52601 );
and \U$52260 ( \52603 , \52596 , \52598 );
nor \U$52261 ( \52604 , \52602 , \52603 );
not \U$52262 ( \52605 , \52213 );
not \U$52263 ( \52606 , \52224 );
or \U$52264 ( \52607 , \52605 , \52606 );
or \U$52265 ( \52608 , \52213 , \52224 );
nand \U$52266 ( \52609 , \52607 , \52608 );
not \U$52267 ( \52610 , \52609 );
not \U$52268 ( \52611 , \52205 );
and \U$52269 ( \52612 , \52610 , \52611 );
and \U$52270 ( \52613 , \52609 , \52205 );
nor \U$52271 ( \52614 , \52612 , \52613 );
xor \U$52272 ( \52615 , \52152 , \52160 );
xor \U$52273 ( \52616 , \52615 , \52168 );
or \U$52274 ( \52617 , \52614 , \52616 );
not \U$52275 ( \52618 , \52616 );
not \U$52276 ( \52619 , \52614 );
or \U$52277 ( \52620 , \52618 , \52619 );
xor \U$52278 ( \52621 , \52178 , \52185 );
xor \U$52279 ( \52622 , \52621 , \52194 );
nand \U$52280 ( \52623 , \52620 , \52622 );
nand \U$52281 ( \52624 , \52617 , \52623 );
xor \U$52282 ( \52625 , \52604 , \52624 );
xor \U$52283 ( \52626 , \52040 , \52047 );
xor \U$52284 ( \52627 , \52626 , \52055 );
xor \U$52285 ( \52628 , \52012 , \52019 );
xor \U$52286 ( \52629 , \52628 , \52027 );
xor \U$52287 ( \52630 , \52627 , \52629 );
xor \U$52288 ( \52631 , \51985 , \51993 );
xor \U$52289 ( \52632 , \52631 , \52001 );
and \U$52290 ( \52633 , \52630 , \52632 );
and \U$52291 ( \52634 , \52627 , \52629 );
nor \U$52292 ( \52635 , \52633 , \52634 );
and \U$52293 ( \52636 , \52625 , \52635 );
and \U$52294 ( \52637 , \52604 , \52624 );
or \U$52295 ( \52638 , \52636 , \52637 );
and \U$52296 ( \52639 , \52594 , \52638 );
and \U$52297 ( \52640 , \52339 , \52593 );
or \U$52298 ( \52641 , \52639 , \52640 );
xor \U$52299 ( \52642 , \51608 , \51627 );
xor \U$52300 ( \52643 , \52642 , \51653 );
not \U$52301 ( \52644 , \52643 );
xor \U$52302 ( \52645 , \52085 , \52112 );
xor \U$52303 ( \52646 , \52645 , \52138 );
not \U$52304 ( \52647 , \52004 );
xor \U$52305 ( \52648 , \52058 , \52030 );
not \U$52306 ( \52649 , \52648 );
or \U$52307 ( \52650 , \52647 , \52649 );
or \U$52308 ( \52651 , \52648 , \52004 );
nand \U$52309 ( \52652 , \52650 , \52651 );
and \U$52310 ( \52653 , \52646 , \52652 );
not \U$52311 ( \52654 , \52653 );
or \U$52312 ( \52655 , \52644 , \52654 );
or \U$52313 ( \52656 , \52653 , \52643 );
xor \U$52314 ( \52657 , \51933 , \51940 );
xor \U$52315 ( \52658 , \52657 , \51947 );
xor \U$52316 ( \52659 , \52171 , \52197 );
xor \U$52317 ( \52660 , \52659 , \52226 );
and \U$52318 ( \52661 , \52658 , \52660 );
not \U$52319 ( \52662 , \51952 );
xor \U$52320 ( \52663 , \51960 , \51955 );
not \U$52321 ( \52664 , \52663 );
or \U$52322 ( \52665 , \52662 , \52664 );
or \U$52323 ( \52666 , \52663 , \51952 );
nand \U$52324 ( \52667 , \52665 , \52666 );
xor \U$52325 ( \52668 , \52171 , \52197 );
xor \U$52326 ( \52669 , \52668 , \52226 );
and \U$52327 ( \52670 , \52667 , \52669 );
and \U$52328 ( \52671 , \52658 , \52667 );
or \U$52329 ( \52672 , \52661 , \52670 , \52671 );
nand \U$52330 ( \52673 , \52656 , \52672 );
nand \U$52331 ( \52674 , \52655 , \52673 );
xor \U$52332 ( \52675 , \52641 , \52674 );
xor \U$52333 ( \52676 , \51950 , \51962 );
xor \U$52334 ( \52677 , \52676 , \51975 );
xor \U$52335 ( \52678 , \51893 , \51903 );
xor \U$52336 ( \52679 , \52678 , \51914 );
xor \U$52337 ( \52680 , \52677 , \52679 );
not \U$52338 ( \52681 , \52236 );
not \U$52339 ( \52682 , \52244 );
or \U$52340 ( \52683 , \52681 , \52682 );
or \U$52341 ( \52684 , \52244 , \52236 );
nand \U$52342 ( \52685 , \52683 , \52684 );
not \U$52343 ( \52686 , \52685 );
not \U$52344 ( \52687 , \52234 );
and \U$52345 ( \52688 , \52686 , \52687 );
and \U$52346 ( \52689 , \52685 , \52234 );
nor \U$52347 ( \52690 , \52688 , \52689 );
and \U$52348 ( \52691 , \52680 , \52690 );
and \U$52349 ( \52692 , \52677 , \52679 );
nor \U$52350 ( \52693 , \52691 , \52692 );
and \U$52351 ( \52694 , \52675 , \52693 );
and \U$52352 ( \52695 , \52641 , \52674 );
or \U$52353 ( \52696 , \52694 , \52695 );
xor \U$52354 ( \52697 , \52323 , \52696 );
xor \U$52355 ( \52698 , \51436 , \51438 );
xor \U$52356 ( \52699 , \52698 , \51443 );
xor \U$52357 ( \52700 , \51879 , \51886 );
xor \U$52358 ( \52701 , \52699 , \52700 );
and \U$52359 ( \52702 , \52697 , \52701 );
and \U$52360 ( \52703 , \52323 , \52696 );
or \U$52361 ( \52704 , \52702 , \52703 );
xor \U$52362 ( \52705 , \51446 , \51760 );
xor \U$52363 ( \52706 , \52705 , \51775 );
xor \U$52364 ( \52707 , \52704 , \52706 );
xor \U$52365 ( \52708 , \51891 , \52267 );
xor \U$52366 ( \52709 , \52708 , \52274 );
and \U$52367 ( \52710 , \52707 , \52709 );
and \U$52368 ( \52711 , \52704 , \52706 );
or \U$52369 ( \52712 , \52710 , \52711 );
nand \U$52370 ( \52713 , \52309 , \52712 );
or \U$52371 ( \52714 , \52298 , \52713 );
xnor \U$52372 ( \52715 , \52713 , \52298 );
xor \U$52373 ( \52716 , \52641 , \52674 );
xor \U$52374 ( \52717 , \52716 , \52693 );
not \U$52375 ( \52718 , \52717 );
xnor \U$52376 ( \52719 , \52672 , \52653 );
not \U$52377 ( \52720 , \52719 );
not \U$52378 ( \52721 , \52643 );
and \U$52379 ( \52722 , \52720 , \52721 );
and \U$52380 ( \52723 , \52719 , \52643 );
nor \U$52381 ( \52724 , \52722 , \52723 );
not \U$52382 ( \52725 , \52060 );
not \U$52383 ( \52726 , \52229 );
or \U$52384 ( \52727 , \52725 , \52726 );
or \U$52385 ( \52728 , \52229 , \52060 );
nand \U$52386 ( \52729 , \52727 , \52728 );
not \U$52387 ( \52730 , \52729 );
not \U$52388 ( \52731 , \52141 );
and \U$52389 ( \52732 , \52730 , \52731 );
and \U$52390 ( \52733 , \52729 , \52141 );
nor \U$52391 ( \52734 , \52732 , \52733 );
xor \U$52392 ( \52735 , \52724 , \52734 );
xor \U$52393 ( \52736 , \52677 , \52679 );
xor \U$52394 ( \52737 , \52736 , \52690 );
xor \U$52395 ( \52738 , \52735 , \52737 );
not \U$52396 ( \52739 , \52738 );
not \U$52397 ( \52740 , \52426 );
not \U$52398 ( \52741 , \52367 );
or \U$52399 ( \52742 , \52740 , \52741 );
or \U$52400 ( \52743 , \52367 , \52426 );
nand \U$52401 ( \52744 , \52742 , \52743 );
not \U$52402 ( \52745 , \52744 );
not \U$52403 ( \52746 , \52395 );
and \U$52404 ( \52747 , \52745 , \52746 );
and \U$52405 ( \52748 , \52744 , \52395 );
nor \U$52406 ( \52749 , \52747 , \52748 );
xor \U$52407 ( \52750 , \52449 , \52476 );
xor \U$52408 ( \52751 , \52750 , \52504 );
or \U$52409 ( \52752 , \52749 , \52751 );
not \U$52410 ( \52753 , \52751 );
not \U$52411 ( \52754 , \52749 );
or \U$52412 ( \52755 , \52753 , \52754 );
xor \U$52413 ( \52756 , \52535 , \52561 );
xor \U$52414 ( \52757 , \52756 , \52587 );
nand \U$52415 ( \52758 , \52755 , \52757 );
nand \U$52416 ( \52759 , \52752 , \52758 );
xor \U$52417 ( \52760 , \52646 , \52652 );
xor \U$52418 ( \52761 , \52759 , \52760 );
xor \U$52419 ( \52762 , \52171 , \52197 );
xor \U$52420 ( \52763 , \52762 , \52226 );
xor \U$52421 ( \52764 , \52658 , \52667 );
xor \U$52422 ( \52765 , \52763 , \52764 );
and \U$52423 ( \52766 , \52761 , \52765 );
and \U$52424 ( \52767 , \52759 , \52760 );
or \U$52425 ( \52768 , \52766 , \52767 );
not \U$52426 ( \52769 , \52768 );
and \U$52427 ( \52770 , \7729 , RI9871578_122);
and \U$52428 ( \52771 , RI9871668_124, \7727 );
nor \U$52429 ( \52772 , \52770 , \52771 );
and \U$52430 ( \52773 , \52772 , \7733 );
not \U$52431 ( \52774 , \52772 );
and \U$52432 ( \52775 , \52774 , \7480 );
nor \U$52433 ( \52776 , \52773 , \52775 );
and \U$52434 ( \52777 , \8486 , RI986eb48_32);
and \U$52435 ( \52778 , RI986ea58_30, \8484 );
nor \U$52436 ( \52779 , \52777 , \52778 );
and \U$52437 ( \52780 , \52779 , \8051 );
not \U$52438 ( \52781 , \52779 );
and \U$52439 ( \52782 , \52781 , \8050 );
nor \U$52440 ( \52783 , \52780 , \52782 );
xor \U$52441 ( \52784 , \52776 , \52783 );
and \U$52442 ( \52785 , \7079 , RI9871758_126);
and \U$52443 ( \52786 , RI9871848_128, \7077 );
nor \U$52444 ( \52787 , \52785 , \52786 );
and \U$52445 ( \52788 , \52787 , \6709 );
not \U$52446 ( \52789 , \52787 );
and \U$52447 ( \52790 , \52789 , \6710 );
nor \U$52448 ( \52791 , \52788 , \52790 );
and \U$52449 ( \52792 , \52784 , \52791 );
and \U$52450 ( \52793 , \52776 , \52783 );
nor \U$52451 ( \52794 , \52792 , \52793 );
and \U$52452 ( \52795 , \6453 , RI9871398_118);
and \U$52453 ( \52796 , RI9871488_120, \6451 );
nor \U$52454 ( \52797 , \52795 , \52796 );
and \U$52455 ( \52798 , \52797 , \6190 );
not \U$52456 ( \52799 , \52797 );
and \U$52457 ( \52800 , \52799 , \6705 );
nor \U$52458 ( \52801 , \52798 , \52800 );
and \U$52459 ( \52802 , \5318 , RI98710c8_112);
and \U$52460 ( \52803 , RI9870d08_104, \5316 );
nor \U$52461 ( \52804 , \52802 , \52803 );
and \U$52462 ( \52805 , \52804 , \5052 );
not \U$52463 ( \52806 , \52804 );
and \U$52464 ( \52807 , \52806 , \5322 );
nor \U$52465 ( \52808 , \52805 , \52807 );
xor \U$52466 ( \52809 , \52801 , \52808 );
and \U$52467 ( \52810 , \5881 , RI98712a8_116);
and \U$52468 ( \52811 , RI98711b8_114, \5879 );
nor \U$52469 ( \52812 , \52810 , \52811 );
and \U$52470 ( \52813 , \52812 , \5594 );
not \U$52471 ( \52814 , \52812 );
and \U$52472 ( \52815 , \52814 , \5885 );
nor \U$52473 ( \52816 , \52813 , \52815 );
and \U$52474 ( \52817 , \52809 , \52816 );
and \U$52475 ( \52818 , \52801 , \52808 );
or \U$52476 ( \52819 , \52817 , \52818 );
xor \U$52477 ( \52820 , \52794 , \52819 );
and \U$52478 ( \52821 , \4203 , RI9870df8_106);
and \U$52479 ( \52822 , RI9870a38_98, \4201 );
nor \U$52480 ( \52823 , \52821 , \52822 );
and \U$52481 ( \52824 , \52823 , \3923 );
not \U$52482 ( \52825 , \52823 );
and \U$52483 ( \52826 , \52825 , \4207 );
nor \U$52484 ( \52827 , \52824 , \52826 );
and \U$52485 ( \52828 , \4710 , RI9870ee8_108);
and \U$52486 ( \52829 , RI9870c18_102, \4708 );
nor \U$52487 ( \52830 , \52828 , \52829 );
not \U$52488 ( \52831 , \52830 );
not \U$52489 ( \52832 , \4519 );
and \U$52490 ( \52833 , \52831 , \52832 );
and \U$52491 ( \52834 , \52830 , \4521 );
nor \U$52492 ( \52835 , \52833 , \52834 );
xor \U$52493 ( \52836 , \52827 , \52835 );
and \U$52494 ( \52837 , \3683 , RI9870fd8_110);
and \U$52495 ( \52838 , RI9870b28_100, \3681 );
nor \U$52496 ( \52839 , \52837 , \52838 );
not \U$52497 ( \52840 , \52839 );
not \U$52498 ( \52841 , \3412 );
and \U$52499 ( \52842 , \52840 , \52841 );
and \U$52500 ( \52843 , \52839 , \3412 );
nor \U$52501 ( \52844 , \52842 , \52843 );
and \U$52502 ( \52845 , \52836 , \52844 );
and \U$52503 ( \52846 , \52827 , \52835 );
nor \U$52504 ( \52847 , \52845 , \52846 );
and \U$52505 ( \52848 , \52820 , \52847 );
and \U$52506 ( \52849 , \52794 , \52819 );
or \U$52507 ( \52850 , \52848 , \52849 );
not \U$52508 ( \52851 , \2935 );
and \U$52509 ( \52852 , \3254 , RI98700d8_78);
and \U$52510 ( \52853 , RI98701c8_80, \3252 );
nor \U$52511 ( \52854 , \52852 , \52853 );
not \U$52512 ( \52855 , \52854 );
or \U$52513 ( \52856 , \52851 , \52855 );
or \U$52514 ( \52857 , \52854 , \2935 );
nand \U$52515 ( \52858 , \52856 , \52857 );
and \U$52516 ( \52859 , \2274 , RI986fe08_72);
and \U$52517 ( \52860 , RI986fd18_70, \2272 );
nor \U$52518 ( \52861 , \52859 , \52860 );
and \U$52519 ( \52862 , \52861 , \2030 );
not \U$52520 ( \52863 , \52861 );
and \U$52521 ( \52864 , \52863 , \2031 );
nor \U$52522 ( \52865 , \52862 , \52864 );
xor \U$52523 ( \52866 , \52858 , \52865 );
and \U$52524 ( \52867 , \2464 , RI986ffe8_76);
and \U$52525 ( \52868 , RI986fef8_74, \2462 );
nor \U$52526 ( \52869 , \52867 , \52868 );
and \U$52527 ( \52870 , \52869 , \2468 );
not \U$52528 ( \52871 , \52869 );
and \U$52529 ( \52872 , \52871 , \2263 );
nor \U$52530 ( \52873 , \52870 , \52872 );
and \U$52531 ( \52874 , \52866 , \52873 );
and \U$52532 ( \52875 , \52858 , \52865 );
or \U$52533 ( \52876 , \52874 , \52875 );
not \U$52534 ( \52877 , \1128 );
and \U$52535 ( \52878 , \1293 , RI98703a8_84);
and \U$52536 ( \52879 , RI98702b8_82, \1291 );
nor \U$52537 ( \52880 , \52878 , \52879 );
not \U$52538 ( \52881 , \52880 );
or \U$52539 ( \52882 , \52877 , \52881 );
or \U$52540 ( \52883 , \52880 , \1301 );
nand \U$52541 ( \52884 , \52882 , \52883 );
and \U$52542 ( \52885 , \776 , RI9870498_86);
and \U$52543 ( \52886 , RI9870588_88, \774 );
nor \U$52544 ( \52887 , \52885 , \52886 );
and \U$52545 ( \52888 , \52887 , \474 );
not \U$52546 ( \52889 , \52887 );
and \U$52547 ( \52890 , \52889 , \451 );
nor \U$52548 ( \52891 , \52888 , \52890 );
and \U$52549 ( \52892 , \52884 , \52891 );
xor \U$52550 ( \52893 , \52876 , \52892 );
and \U$52551 ( \52894 , \1329 , RI9870768_92);
and \U$52552 ( \52895 , RI9870678_90, \1327 );
nor \U$52553 ( \52896 , \52894 , \52895 );
and \U$52554 ( \52897 , \52896 , \1336 );
not \U$52555 ( \52898 , \52896 );
and \U$52556 ( \52899 , \52898 , \1337 );
nor \U$52557 ( \52900 , \52897 , \52899 );
and \U$52558 ( \52901 , \1311 , RI9870948_96);
and \U$52559 ( \52902 , RI9870858_94, \1309 );
nor \U$52560 ( \52903 , \52901 , \52902 );
and \U$52561 ( \52904 , \52903 , \1458 );
not \U$52562 ( \52905 , \52903 );
and \U$52563 ( \52906 , \52905 , \1318 );
nor \U$52564 ( \52907 , \52904 , \52906 );
xor \U$52565 ( \52908 , \52900 , \52907 );
not \U$52566 ( \52909 , \2034 );
and \U$52567 ( \52910 , \2042 , RI986fb38_66);
and \U$52568 ( \52911 , RI986fc28_68, \2040 );
nor \U$52569 ( \52912 , \52910 , \52911 );
not \U$52570 ( \52913 , \52912 );
or \U$52571 ( \52914 , \52909 , \52913 );
or \U$52572 ( \52915 , \52912 , \2034 );
nand \U$52573 ( \52916 , \52914 , \52915 );
and \U$52574 ( \52917 , \52908 , \52916 );
and \U$52575 ( \52918 , \52900 , \52907 );
or \U$52576 ( \52919 , \52917 , \52918 );
and \U$52577 ( \52920 , \52893 , \52919 );
and \U$52578 ( \52921 , \52876 , \52892 );
or \U$52579 ( \52922 , \52920 , \52921 );
xor \U$52580 ( \52923 , \52850 , \52922 );
and \U$52581 ( \52924 , \12293 , RI986f2c8_48);
and \U$52582 ( \52925 , RI986f1d8_46, \12291 );
nor \U$52583 ( \52926 , \52924 , \52925 );
and \U$52584 ( \52927 , \52926 , \11686 );
not \U$52585 ( \52928 , \52926 );
and \U$52586 ( \52929 , \52928 , \11687 );
nor \U$52587 ( \52930 , \52927 , \52929 );
and \U$52588 ( \52931 , \13045 , RI986e5a8_20);
and \U$52589 ( \52932 , RI986e4b8_18, \13043 );
nor \U$52590 ( \52933 , \52931 , \52932 );
and \U$52591 ( \52934 , \52933 , \12619 );
not \U$52592 ( \52935 , \52933 );
and \U$52593 ( \52936 , \52935 , \13047 );
nor \U$52594 ( \52937 , \52934 , \52936 );
xor \U$52595 ( \52938 , \52930 , \52937 );
and \U$52596 ( \52939 , \11696 , RI986f0e8_44);
and \U$52597 ( \52940 , RI986eff8_42, \11694 );
nor \U$52598 ( \52941 , \52939 , \52940 );
and \U$52599 ( \52942 , \52941 , \11702 );
not \U$52600 ( \52943 , \52941 );
and \U$52601 ( \52944 , \52943 , \10965 );
nor \U$52602 ( \52945 , \52942 , \52944 );
and \U$52603 ( \52946 , \52938 , \52945 );
and \U$52604 ( \52947 , \52930 , \52937 );
nor \U$52605 ( \52948 , \52946 , \52947 );
and \U$52606 ( \52949 , \15780 , RI986fa48_64);
and \U$52607 ( \52950 , RI986f958_62, RI9873648_192);
nor \U$52608 ( \52951 , \52949 , \52950 );
not \U$52609 ( \52952 , \52951 );
not \U$52610 ( \52953 , RI9873558_190);
and \U$52611 ( \52954 , \52952 , \52953 );
and \U$52612 ( \52955 , \52951 , RI9873558_190);
nor \U$52613 ( \52956 , \52954 , \52955 );
and \U$52614 ( \52957 , \14937 , RI986f868_60);
and \U$52615 ( \52958 , RI986f778_58, \14935 );
nor \U$52616 ( \52959 , \52957 , \52958 );
and \U$52617 ( \52960 , \52959 , \14538 );
not \U$52618 ( \52961 , \52959 );
and \U$52619 ( \52962 , \52961 , \14539 );
nor \U$52620 ( \52963 , \52960 , \52962 );
xor \U$52621 ( \52964 , \52956 , \52963 );
and \U$52622 ( \52965 , \13882 , RI986e788_24);
and \U$52623 ( \52966 , RI986e698_22, \13880 );
nor \U$52624 ( \52967 , \52965 , \52966 );
and \U$52625 ( \52968 , \52967 , \13359 );
not \U$52626 ( \52969 , \52967 );
and \U$52627 ( \52970 , \52969 , \13358 );
nor \U$52628 ( \52971 , \52968 , \52970 );
and \U$52629 ( \52972 , \52964 , \52971 );
and \U$52630 ( \52973 , \52956 , \52963 );
nor \U$52631 ( \52974 , \52972 , \52973 );
xor \U$52632 ( \52975 , \52948 , \52974 );
and \U$52633 ( \52976 , \9505 , RI986ef08_40);
and \U$52634 ( \52977 , RI986ee18_38, \9503 );
nor \U$52635 ( \52978 , \52976 , \52977 );
and \U$52636 ( \52979 , \52978 , \9510 );
not \U$52637 ( \52980 , \52978 );
and \U$52638 ( \52981 , \52980 , \9513 );
nor \U$52639 ( \52982 , \52979 , \52981 );
and \U$52640 ( \52983 , \9237 , RI986e968_28);
and \U$52641 ( \52984 , RI986e878_26, \9235 );
nor \U$52642 ( \52985 , \52983 , \52984 );
and \U$52643 ( \52986 , \52985 , \9241 );
not \U$52644 ( \52987 , \52985 );
and \U$52645 ( \52988 , \52987 , \8836 );
nor \U$52646 ( \52989 , \52986 , \52988 );
xor \U$52647 ( \52990 , \52982 , \52989 );
and \U$52648 ( \52991 , \10424 , RI986ec38_34);
and \U$52649 ( \52992 , RI986ed28_36, \10422 );
nor \U$52650 ( \52993 , \52991 , \52992 );
and \U$52651 ( \52994 , \52993 , \9840 );
not \U$52652 ( \52995 , \52993 );
and \U$52653 ( \52996 , \52995 , \10428 );
nor \U$52654 ( \52997 , \52994 , \52996 );
and \U$52655 ( \52998 , \52990 , \52997 );
and \U$52656 ( \52999 , \52982 , \52989 );
or \U$52657 ( \53000 , \52998 , \52999 );
and \U$52658 ( \53001 , \52975 , \53000 );
and \U$52659 ( \53002 , \52948 , \52974 );
or \U$52660 ( \53003 , \53001 , \53002 );
and \U$52661 ( \53004 , \52923 , \53003 );
and \U$52662 ( \53005 , \52850 , \52922 );
nor \U$52663 ( \53006 , \53004 , \53005 );
not \U$52664 ( \53007 , \52484 );
xor \U$52665 ( \53008 , \52502 , \52492 );
not \U$52666 ( \53009 , \53008 );
or \U$52667 ( \53010 , \53007 , \53009 );
or \U$52668 ( \53011 , \53008 , \52484 );
nand \U$52669 ( \53012 , \53010 , \53011 );
not \U$52670 ( \53013 , \52456 );
xor \U$52671 ( \53014 , \52474 , \52464 );
not \U$52672 ( \53015 , \53014 );
or \U$52673 ( \53016 , \53013 , \53015 );
or \U$52674 ( \53017 , \53014 , \52456 );
nand \U$52675 ( \53018 , \53016 , \53017 );
xor \U$52676 ( \53019 , \53012 , \53018 );
xor \U$52677 ( \53020 , \52569 , \52576 );
xor \U$52678 ( \53021 , \53020 , \52584 );
and \U$52679 ( \53022 , \53019 , \53021 );
and \U$52680 ( \53023 , \53012 , \53018 );
nor \U$52681 ( \53024 , \53022 , \53023 );
not \U$52682 ( \53025 , \52346 );
xor \U$52683 ( \53026 , \52365 , \52354 );
not \U$52684 ( \53027 , \53026 );
or \U$52685 ( \53028 , \53025 , \53027 );
or \U$52686 ( \53029 , \53026 , \52346 );
nand \U$52687 ( \53030 , \53028 , \53029 );
nand \U$52688 ( \53031 , RI9870498_86, \436 );
and \U$52689 ( \53032 , \53031 , \444 );
not \U$52690 ( \53033 , \53031 );
and \U$52691 ( \53034 , \53033 , \443 );
nor \U$52692 ( \53035 , \53032 , \53034 );
xor \U$52693 ( \53036 , \53030 , \53035 );
not \U$52694 ( \53037 , \52374 );
xor \U$52695 ( \53038 , \52393 , \52382 );
not \U$52696 ( \53039 , \53038 );
or \U$52697 ( \53040 , \53037 , \53039 );
or \U$52698 ( \53041 , \53038 , \52374 );
nand \U$52699 ( \53042 , \53040 , \53041 );
and \U$52700 ( \53043 , \53036 , \53042 );
and \U$52701 ( \53044 , \53030 , \53035 );
nor \U$52702 ( \53045 , \53043 , \53044 );
xor \U$52703 ( \53046 , \53024 , \53045 );
xor \U$52704 ( \53047 , \52543 , \52550 );
xor \U$52705 ( \53048 , \53047 , \52558 );
not \U$52706 ( \53049 , \53048 );
not \U$52707 ( \53050 , \52522 );
not \U$52708 ( \53051 , \52533 );
or \U$52709 ( \53052 , \53050 , \53051 );
or \U$52710 ( \53053 , \52522 , \52533 );
nand \U$52711 ( \53054 , \53052 , \53053 );
not \U$52712 ( \53055 , \53054 );
not \U$52713 ( \53056 , \52515 );
and \U$52714 ( \53057 , \53055 , \53056 );
and \U$52715 ( \53058 , \53054 , \52515 );
nor \U$52716 ( \53059 , \53057 , \53058 );
not \U$52717 ( \53060 , \53059 );
and \U$52718 ( \53061 , \53049 , \53060 );
and \U$52719 ( \53062 , \53059 , \53048 );
xor \U$52720 ( \53063 , \52407 , \52415 );
xor \U$52721 ( \53064 , \53063 , \52423 );
nor \U$52722 ( \53065 , \53062 , \53064 );
nor \U$52723 ( \53066 , \53061 , \53065 );
and \U$52724 ( \53067 , \53046 , \53066 );
and \U$52725 ( \53068 , \53024 , \53045 );
or \U$52726 ( \53069 , \53067 , \53068 );
xor \U$52727 ( \53070 , \53006 , \53069 );
xor \U$52728 ( \53071 , \52627 , \52629 );
xor \U$52729 ( \53072 , \53071 , \52632 );
not \U$52730 ( \53073 , \52616 );
not \U$52731 ( \53074 , \52622 );
or \U$52732 ( \53075 , \53073 , \53074 );
or \U$52733 ( \53076 , \52616 , \52622 );
nand \U$52734 ( \53077 , \53075 , \53076 );
not \U$52735 ( \53078 , \53077 );
not \U$52736 ( \53079 , \52614 );
and \U$52737 ( \53080 , \53078 , \53079 );
and \U$52738 ( \53081 , \53077 , \52614 );
nor \U$52739 ( \53082 , \53080 , \53081 );
xor \U$52740 ( \53083 , \53072 , \53082 );
xor \U$52741 ( \53084 , \52596 , \52598 );
xor \U$52742 ( \53085 , \53084 , \52601 );
and \U$52743 ( \53086 , \53083 , \53085 );
and \U$52744 ( \53087 , \53072 , \53082 );
or \U$52745 ( \53088 , \53086 , \53087 );
and \U$52746 ( \53089 , \53070 , \53088 );
and \U$52747 ( \53090 , \53006 , \53069 );
nor \U$52748 ( \53091 , \53089 , \53090 );
xor \U$52749 ( \53092 , \51635 , \51642 );
xor \U$52750 ( \53093 , \53092 , \51650 );
xor \U$52751 ( \53094 , \52325 , \52334 );
xor \U$52752 ( \53095 , \53093 , \53094 );
not \U$52753 ( \53096 , \53095 );
xor \U$52754 ( \53097 , \52428 , \52507 );
xor \U$52755 ( \53098 , \53097 , \52590 );
not \U$52756 ( \53099 , \53098 );
or \U$52757 ( \53100 , \53096 , \53099 );
or \U$52758 ( \53101 , \53098 , \53095 );
xor \U$52759 ( \53102 , \52604 , \52624 );
xor \U$52760 ( \53103 , \53102 , \52635 );
nand \U$52761 ( \53104 , \53101 , \53103 );
nand \U$52762 ( \53105 , \53100 , \53104 );
xnor \U$52763 ( \53106 , \53091 , \53105 );
not \U$52764 ( \53107 , \53106 );
or \U$52765 ( \53108 , \52769 , \53107 );
or \U$52766 ( \53109 , \53106 , \52768 );
nand \U$52767 ( \53110 , \53108 , \53109 );
nand \U$52768 ( \53111 , \52739 , \53110 );
nand \U$52769 ( \53112 , \52718 , \53111 );
not \U$52770 ( \53113 , \52751 );
not \U$52771 ( \53114 , \52757 );
or \U$52772 ( \53115 , \53113 , \53114 );
or \U$52773 ( \53116 , \52757 , \52751 );
nand \U$52774 ( \53117 , \53115 , \53116 );
not \U$52775 ( \53118 , \53117 );
not \U$52776 ( \53119 , \52749 );
and \U$52777 ( \53120 , \53118 , \53119 );
and \U$52778 ( \53121 , \53117 , \52749 );
nor \U$52779 ( \53122 , \53120 , \53121 );
xor \U$52780 ( \53123 , \52794 , \52819 );
xor \U$52781 ( \53124 , \53123 , \52847 );
xor \U$52782 ( \53125 , \52876 , \52892 );
xor \U$52783 ( \53126 , \53125 , \52919 );
and \U$52784 ( \53127 , \53124 , \53126 );
xor \U$52785 ( \53128 , \53030 , \53035 );
xor \U$52786 ( \53129 , \53128 , \53042 );
xor \U$52787 ( \53130 , \52876 , \52892 );
xor \U$52788 ( \53131 , \53130 , \52919 );
and \U$52789 ( \53132 , \53129 , \53131 );
and \U$52790 ( \53133 , \53124 , \53129 );
or \U$52791 ( \53134 , \53127 , \53132 , \53133 );
not \U$52792 ( \53135 , \53134 );
xor \U$52793 ( \53136 , \53122 , \53135 );
xor \U$52794 ( \53137 , \53072 , \53082 );
xor \U$52795 ( \53138 , \53137 , \53085 );
and \U$52796 ( \53139 , \53136 , \53138 );
and \U$52797 ( \53140 , \53122 , \53135 );
or \U$52798 ( \53141 , \53139 , \53140 );
xor \U$52799 ( \53142 , \53024 , \53045 );
xor \U$52800 ( \53143 , \53142 , \53066 );
not \U$52801 ( \53144 , \53143 );
xor \U$52802 ( \53145 , \52850 , \52922 );
xor \U$52803 ( \53146 , \53145 , \53003 );
nand \U$52804 ( \53147 , \53144 , \53146 );
or \U$52805 ( \53148 , \53141 , \53147 );
not \U$52806 ( \53149 , \53147 );
not \U$52807 ( \53150 , \53141 );
or \U$52808 ( \53151 , \53149 , \53150 );
xor \U$52809 ( \53152 , \52956 , \52963 );
xor \U$52810 ( \53153 , \53152 , \52971 );
xor \U$52811 ( \53154 , \52930 , \52937 );
xor \U$52812 ( \53155 , \53154 , \52945 );
or \U$52813 ( \53156 , \53153 , \53155 );
not \U$52814 ( \53157 , \53155 );
not \U$52815 ( \53158 , \53153 );
or \U$52816 ( \53159 , \53157 , \53158 );
xor \U$52817 ( \53160 , \52982 , \52989 );
xor \U$52818 ( \53161 , \53160 , \52997 );
nand \U$52819 ( \53162 , \53159 , \53161 );
nand \U$52820 ( \53163 , \53156 , \53162 );
xor \U$52821 ( \53164 , \52884 , \52891 );
not \U$52822 ( \53165 , \53164 );
xor \U$52823 ( \53166 , \52858 , \52865 );
xor \U$52824 ( \53167 , \53166 , \52873 );
not \U$52825 ( \53168 , \53167 );
or \U$52826 ( \53169 , \53165 , \53168 );
or \U$52827 ( \53170 , \53167 , \53164 );
xor \U$52828 ( \53171 , \52900 , \52907 );
xor \U$52829 ( \53172 , \53171 , \52916 );
nand \U$52830 ( \53173 , \53170 , \53172 );
nand \U$52831 ( \53174 , \53169 , \53173 );
xor \U$52832 ( \53175 , \53163 , \53174 );
xor \U$52833 ( \53176 , \52827 , \52835 );
xor \U$52834 ( \53177 , \53176 , \52844 );
xor \U$52835 ( \53178 , \52776 , \52783 );
xor \U$52836 ( \53179 , \53178 , \52791 );
or \U$52837 ( \53180 , \53177 , \53179 );
not \U$52838 ( \53181 , \53179 );
not \U$52839 ( \53182 , \53177 );
or \U$52840 ( \53183 , \53181 , \53182 );
xor \U$52841 ( \53184 , \52801 , \52808 );
xor \U$52842 ( \53185 , \53184 , \52816 );
nand \U$52843 ( \53186 , \53183 , \53185 );
nand \U$52844 ( \53187 , \53180 , \53186 );
and \U$52845 ( \53188 , \53175 , \53187 );
and \U$52846 ( \53189 , \53163 , \53174 );
or \U$52847 ( \53190 , \53188 , \53189 );
and \U$52848 ( \53191 , \9505 , RI986e878_26);
and \U$52849 ( \53192 , RI986ef08_40, \9503 );
nor \U$52850 ( \53193 , \53191 , \53192 );
and \U$52851 ( \53194 , \53193 , \9510 );
not \U$52852 ( \53195 , \53193 );
and \U$52853 ( \53196 , \53195 , \9513 );
nor \U$52854 ( \53197 , \53194 , \53196 );
and \U$52855 ( \53198 , \10424 , RI986ee18_38);
and \U$52856 ( \53199 , RI986ec38_34, \10422 );
nor \U$52857 ( \53200 , \53198 , \53199 );
and \U$52858 ( \53201 , \53200 , \9840 );
not \U$52859 ( \53202 , \53200 );
and \U$52860 ( \53203 , \53202 , \10428 );
nor \U$52861 ( \53204 , \53201 , \53203 );
xor \U$52862 ( \53205 , \53197 , \53204 );
and \U$52863 ( \53206 , \11696 , RI986ed28_36);
and \U$52864 ( \53207 , RI986f0e8_44, \11694 );
nor \U$52865 ( \53208 , \53206 , \53207 );
and \U$52866 ( \53209 , \53208 , \10965 );
not \U$52867 ( \53210 , \53208 );
and \U$52868 ( \53211 , \53210 , \11702 );
nor \U$52869 ( \53212 , \53209 , \53211 );
and \U$52870 ( \53213 , \53205 , \53212 );
and \U$52871 ( \53214 , \53197 , \53204 );
or \U$52872 ( \53215 , \53213 , \53214 );
not \U$52873 ( \53216 , RI9873558_190);
and \U$52874 ( \53217 , \15780 , RI986f778_58);
and \U$52875 ( \53218 , RI986fa48_64, RI9873648_192);
nor \U$52876 ( \53219 , \53217 , \53218 );
not \U$52877 ( \53220 , \53219 );
or \U$52878 ( \53221 , \53216 , \53220 );
or \U$52879 ( \53222 , \53219 , RI9873558_190);
nand \U$52880 ( \53223 , \53221 , \53222 );
xor \U$52881 ( \53224 , \53223 , \451 );
and \U$52882 ( \53225 , \14937 , RI986e698_22);
and \U$52883 ( \53226 , RI986f868_60, \14935 );
nor \U$52884 ( \53227 , \53225 , \53226 );
and \U$52885 ( \53228 , \53227 , \14539 );
not \U$52886 ( \53229 , \53227 );
and \U$52887 ( \53230 , \53229 , \14538 );
nor \U$52888 ( \53231 , \53228 , \53230 );
and \U$52889 ( \53232 , \53224 , \53231 );
and \U$52890 ( \53233 , \53223 , \451 );
or \U$52891 ( \53234 , \53232 , \53233 );
xor \U$52892 ( \53235 , \53215 , \53234 );
and \U$52893 ( \53236 , \13045 , RI986f1d8_46);
and \U$52894 ( \53237 , RI986e5a8_20, \13043 );
nor \U$52895 ( \53238 , \53236 , \53237 );
and \U$52896 ( \53239 , \53238 , \13047 );
not \U$52897 ( \53240 , \53238 );
and \U$52898 ( \53241 , \53240 , \12619 );
nor \U$52899 ( \53242 , \53239 , \53241 );
and \U$52900 ( \53243 , \12293 , RI986eff8_42);
and \U$52901 ( \53244 , RI986f2c8_48, \12291 );
nor \U$52902 ( \53245 , \53243 , \53244 );
and \U$52903 ( \53246 , \53245 , \11687 );
not \U$52904 ( \53247 , \53245 );
and \U$52905 ( \53248 , \53247 , \11686 );
nor \U$52906 ( \53249 , \53246 , \53248 );
xor \U$52907 ( \53250 , \53242 , \53249 );
and \U$52908 ( \53251 , \13882 , RI986e4b8_18);
and \U$52909 ( \53252 , RI986e788_24, \13880 );
nor \U$52910 ( \53253 , \53251 , \53252 );
and \U$52911 ( \53254 , \53253 , \13358 );
not \U$52912 ( \53255 , \53253 );
and \U$52913 ( \53256 , \53255 , \13359 );
nor \U$52914 ( \53257 , \53254 , \53256 );
and \U$52915 ( \53258 , \53250 , \53257 );
and \U$52916 ( \53259 , \53242 , \53249 );
or \U$52917 ( \53260 , \53258 , \53259 );
and \U$52918 ( \53261 , \53235 , \53260 );
and \U$52919 ( \53262 , \53215 , \53234 );
or \U$52920 ( \53263 , \53261 , \53262 );
and \U$52921 ( \53264 , \2274 , RI986fc28_68);
and \U$52922 ( \53265 , RI986fe08_72, \2272 );
nor \U$52923 ( \53266 , \53264 , \53265 );
and \U$52924 ( \53267 , \53266 , \2030 );
not \U$52925 ( \53268 , \53266 );
and \U$52926 ( \53269 , \53268 , \2031 );
nor \U$52927 ( \53270 , \53267 , \53269 );
and \U$52928 ( \53271 , \1311 , RI9870678_90);
and \U$52929 ( \53272 , RI9870948_96, \1309 );
nor \U$52930 ( \53273 , \53271 , \53272 );
and \U$52931 ( \53274 , \53273 , \1458 );
not \U$52932 ( \53275 , \53273 );
and \U$52933 ( \53276 , \53275 , \1318 );
nor \U$52934 ( \53277 , \53274 , \53276 );
xor \U$52935 ( \53278 , \53270 , \53277 );
not \U$52936 ( \53279 , \2034 );
and \U$52937 ( \53280 , \2042 , RI9870858_94);
and \U$52938 ( \53281 , RI986fb38_66, \2040 );
nor \U$52939 ( \53282 , \53280 , \53281 );
not \U$52940 ( \53283 , \53282 );
or \U$52941 ( \53284 , \53279 , \53283 );
or \U$52942 ( \53285 , \53282 , \2034 );
nand \U$52943 ( \53286 , \53284 , \53285 );
and \U$52944 ( \53287 , \53278 , \53286 );
and \U$52945 ( \53288 , \53270 , \53277 );
or \U$52946 ( \53289 , \53287 , \53288 );
not \U$52947 ( \53290 , \1301 );
and \U$52948 ( \53291 , \1293 , RI9870588_88);
and \U$52949 ( \53292 , RI98703a8_84, \1291 );
nor \U$52950 ( \53293 , \53291 , \53292 );
not \U$52951 ( \53294 , \53293 );
or \U$52952 ( \53295 , \53290 , \53294 );
or \U$52953 ( \53296 , \53293 , \1128 );
nand \U$52954 ( \53297 , \53295 , \53296 );
nand \U$52955 ( \53298 , RI9870498_86, \774 );
and \U$52956 ( \53299 , \53298 , \474 );
not \U$52957 ( \53300 , \53298 );
and \U$52958 ( \53301 , \53300 , \451 );
nor \U$52959 ( \53302 , \53299 , \53301 );
xor \U$52960 ( \53303 , \53297 , \53302 );
and \U$52961 ( \53304 , \1329 , RI98702b8_82);
and \U$52962 ( \53305 , RI9870768_92, \1327 );
nor \U$52963 ( \53306 , \53304 , \53305 );
and \U$52964 ( \53307 , \53306 , \1336 );
not \U$52965 ( \53308 , \53306 );
and \U$52966 ( \53309 , \53308 , \1337 );
nor \U$52967 ( \53310 , \53307 , \53309 );
and \U$52968 ( \53311 , \53303 , \53310 );
and \U$52969 ( \53312 , \53297 , \53302 );
or \U$52970 ( \53313 , \53311 , \53312 );
xor \U$52971 ( \53314 , \53289 , \53313 );
and \U$52972 ( \53315 , \2464 , RI986fd18_70);
and \U$52973 ( \53316 , RI986ffe8_76, \2462 );
nor \U$52974 ( \53317 , \53315 , \53316 );
and \U$52975 ( \53318 , \53317 , \2468 );
not \U$52976 ( \53319 , \53317 );
and \U$52977 ( \53320 , \53319 , \2263 );
nor \U$52978 ( \53321 , \53318 , \53320 );
not \U$52979 ( \53322 , \2935 );
and \U$52980 ( \53323 , \3254 , RI986fef8_74);
and \U$52981 ( \53324 , RI98700d8_78, \3252 );
nor \U$52982 ( \53325 , \53323 , \53324 );
not \U$52983 ( \53326 , \53325 );
or \U$52984 ( \53327 , \53322 , \53326 );
or \U$52985 ( \53328 , \53325 , \3406 );
nand \U$52986 ( \53329 , \53327 , \53328 );
xor \U$52987 ( \53330 , \53321 , \53329 );
not \U$52988 ( \53331 , \3412 );
and \U$52989 ( \53332 , \3683 , RI98701c8_80);
and \U$52990 ( \53333 , RI9870fd8_110, \3681 );
nor \U$52991 ( \53334 , \53332 , \53333 );
not \U$52992 ( \53335 , \53334 );
or \U$52993 ( \53336 , \53331 , \53335 );
or \U$52994 ( \53337 , \53334 , \3918 );
nand \U$52995 ( \53338 , \53336 , \53337 );
and \U$52996 ( \53339 , \53330 , \53338 );
and \U$52997 ( \53340 , \53321 , \53329 );
or \U$52998 ( \53341 , \53339 , \53340 );
and \U$52999 ( \53342 , \53314 , \53341 );
and \U$53000 ( \53343 , \53289 , \53313 );
or \U$53001 ( \53344 , \53342 , \53343 );
xor \U$53002 ( \53345 , \53263 , \53344 );
and \U$53003 ( \53346 , \7079 , RI9871488_120);
and \U$53004 ( \53347 , RI9871758_126, \7077 );
nor \U$53005 ( \53348 , \53346 , \53347 );
and \U$53006 ( \53349 , \53348 , \6710 );
not \U$53007 ( \53350 , \53348 );
and \U$53008 ( \53351 , \53350 , \6709 );
nor \U$53009 ( \53352 , \53349 , \53351 );
and \U$53010 ( \53353 , \5881 , RI9870d08_104);
and \U$53011 ( \53354 , RI98712a8_116, \5879 );
nor \U$53012 ( \53355 , \53353 , \53354 );
and \U$53013 ( \53356 , \53355 , \5594 );
not \U$53014 ( \53357 , \53355 );
and \U$53015 ( \53358 , \53357 , \5885 );
nor \U$53016 ( \53359 , \53356 , \53358 );
xor \U$53017 ( \53360 , \53352 , \53359 );
and \U$53018 ( \53361 , \6453 , RI98711b8_114);
and \U$53019 ( \53362 , RI9871398_118, \6451 );
nor \U$53020 ( \53363 , \53361 , \53362 );
and \U$53021 ( \53364 , \53363 , \6190 );
not \U$53022 ( \53365 , \53363 );
and \U$53023 ( \53366 , \53365 , \6180 );
nor \U$53024 ( \53367 , \53364 , \53366 );
and \U$53025 ( \53368 , \53360 , \53367 );
and \U$53026 ( \53369 , \53352 , \53359 );
or \U$53027 ( \53370 , \53368 , \53369 );
and \U$53028 ( \53371 , \5318 , RI9870c18_102);
and \U$53029 ( \53372 , RI98710c8_112, \5316 );
nor \U$53030 ( \53373 , \53371 , \53372 );
and \U$53031 ( \53374 , \53373 , \5052 );
not \U$53032 ( \53375 , \53373 );
and \U$53033 ( \53376 , \53375 , \5322 );
nor \U$53034 ( \53377 , \53374 , \53376 );
and \U$53035 ( \53378 , \4203 , RI9870b28_100);
and \U$53036 ( \53379 , RI9870df8_106, \4201 );
nor \U$53037 ( \53380 , \53378 , \53379 );
and \U$53038 ( \53381 , \53380 , \4207 );
not \U$53039 ( \53382 , \53380 );
and \U$53040 ( \53383 , \53382 , \3923 );
nor \U$53041 ( \53384 , \53381 , \53383 );
xor \U$53042 ( \53385 , \53377 , \53384 );
not \U$53043 ( \53386 , \4521 );
and \U$53044 ( \53387 , \4710 , RI9870a38_98);
and \U$53045 ( \53388 , RI9870ee8_108, \4708 );
nor \U$53046 ( \53389 , \53387 , \53388 );
not \U$53047 ( \53390 , \53389 );
or \U$53048 ( \53391 , \53386 , \53390 );
or \U$53049 ( \53392 , \53389 , \4521 );
nand \U$53050 ( \53393 , \53391 , \53392 );
and \U$53051 ( \53394 , \53385 , \53393 );
and \U$53052 ( \53395 , \53377 , \53384 );
or \U$53053 ( \53396 , \53394 , \53395 );
xor \U$53054 ( \53397 , \53370 , \53396 );
and \U$53055 ( \53398 , \8486 , RI9871668_124);
and \U$53056 ( \53399 , RI986eb48_32, \8484 );
nor \U$53057 ( \53400 , \53398 , \53399 );
and \U$53058 ( \53401 , \53400 , \8050 );
not \U$53059 ( \53402 , \53400 );
and \U$53060 ( \53403 , \53402 , \8051 );
nor \U$53061 ( \53404 , \53401 , \53403 );
and \U$53062 ( \53405 , \7729 , RI9871848_128);
and \U$53063 ( \53406 , RI9871578_122, \7727 );
nor \U$53064 ( \53407 , \53405 , \53406 );
and \U$53065 ( \53408 , \53407 , \7480 );
not \U$53066 ( \53409 , \53407 );
and \U$53067 ( \53410 , \53409 , \7733 );
nor \U$53068 ( \53411 , \53408 , \53410 );
xor \U$53069 ( \53412 , \53404 , \53411 );
and \U$53070 ( \53413 , \9237 , RI986ea58_30);
and \U$53071 ( \53414 , RI986e968_28, \9235 );
nor \U$53072 ( \53415 , \53413 , \53414 );
and \U$53073 ( \53416 , \53415 , \9241 );
not \U$53074 ( \53417 , \53415 );
and \U$53075 ( \53418 , \53417 , \8836 );
nor \U$53076 ( \53419 , \53416 , \53418 );
and \U$53077 ( \53420 , \53412 , \53419 );
and \U$53078 ( \53421 , \53404 , \53411 );
or \U$53079 ( \53422 , \53420 , \53421 );
and \U$53080 ( \53423 , \53397 , \53422 );
and \U$53081 ( \53424 , \53370 , \53396 );
or \U$53082 ( \53425 , \53423 , \53424 );
and \U$53083 ( \53426 , \53345 , \53425 );
and \U$53084 ( \53427 , \53263 , \53344 );
or \U$53085 ( \53428 , \53426 , \53427 );
xor \U$53086 ( \53429 , \53190 , \53428 );
not \U$53087 ( \53430 , \53059 );
xor \U$53088 ( \53431 , \53064 , \53048 );
not \U$53089 ( \53432 , \53431 );
or \U$53090 ( \53433 , \53430 , \53432 );
or \U$53091 ( \53434 , \53431 , \53059 );
nand \U$53092 ( \53435 , \53433 , \53434 );
not \U$53093 ( \53436 , \443 );
xnor \U$53094 ( \53437 , \52447 , \52436 );
not \U$53095 ( \53438 , \53437 );
or \U$53096 ( \53439 , \53436 , \53438 );
or \U$53097 ( \53440 , \53437 , \443 );
nand \U$53098 ( \53441 , \53439 , \53440 );
xor \U$53099 ( \53442 , \53435 , \53441 );
xor \U$53100 ( \53443 , \53012 , \53018 );
xor \U$53101 ( \53444 , \53443 , \53021 );
and \U$53102 ( \53445 , \53442 , \53444 );
and \U$53103 ( \53446 , \53435 , \53441 );
or \U$53104 ( \53447 , \53445 , \53446 );
and \U$53105 ( \53448 , \53429 , \53447 );
and \U$53106 ( \53449 , \53190 , \53428 );
or \U$53107 ( \53450 , \53448 , \53449 );
nand \U$53108 ( \53451 , \53151 , \53450 );
nand \U$53109 ( \53452 , \53148 , \53451 );
xor \U$53110 ( \53453 , \52339 , \52593 );
xor \U$53111 ( \53454 , \53453 , \52638 );
xor \U$53112 ( \53455 , \53452 , \53454 );
xnor \U$53113 ( \53456 , \53103 , \53098 );
not \U$53114 ( \53457 , \53456 );
not \U$53115 ( \53458 , \53095 );
and \U$53116 ( \53459 , \53457 , \53458 );
and \U$53117 ( \53460 , \53456 , \53095 );
nor \U$53118 ( \53461 , \53459 , \53460 );
xor \U$53119 ( \53462 , \53006 , \53069 );
xor \U$53120 ( \53463 , \53462 , \53088 );
or \U$53121 ( \53464 , \53461 , \53463 );
not \U$53122 ( \53465 , \53463 );
not \U$53123 ( \53466 , \53461 );
or \U$53124 ( \53467 , \53465 , \53466 );
xor \U$53125 ( \53468 , \52759 , \52760 );
xor \U$53126 ( \53469 , \53468 , \52765 );
nand \U$53127 ( \53470 , \53467 , \53469 );
nand \U$53128 ( \53471 , \53464 , \53470 );
and \U$53129 ( \53472 , \53455 , \53471 );
and \U$53130 ( \53473 , \53452 , \53454 );
or \U$53131 ( \53474 , \53472 , \53473 );
and \U$53132 ( \53475 , \53112 , \53474 );
not \U$53133 ( \53476 , \53111 );
and \U$53134 ( \53477 , \52717 , \53476 );
nor \U$53135 ( \53478 , \53475 , \53477 );
not \U$53136 ( \53479 , \53478 );
xor \U$53137 ( \53480 , \52323 , \52696 );
xor \U$53138 ( \53481 , \53480 , \52701 );
xor \U$53139 ( \53482 , \52724 , \52734 );
and \U$53140 ( \53483 , \53482 , \52737 );
and \U$53141 ( \53484 , \52724 , \52734 );
or \U$53142 ( \53485 , \53483 , \53484 );
and \U$53143 ( \53486 , \53105 , \53091 );
or \U$53144 ( \53487 , \53105 , \53091 );
and \U$53145 ( \53488 , \52768 , \53487 );
nor \U$53146 ( \53489 , \53486 , \53488 );
or \U$53147 ( \53490 , \53485 , \53489 );
not \U$53148 ( \53491 , \53489 );
not \U$53149 ( \53492 , \53485 );
or \U$53150 ( \53493 , \53491 , \53492 );
xor \U$53151 ( \53494 , \51917 , \51919 );
xor \U$53152 ( \53495 , \53494 , \51924 );
xor \U$53153 ( \53496 , \52311 , \52318 );
xor \U$53154 ( \53497 , \53495 , \53496 );
nand \U$53155 ( \53498 , \53493 , \53497 );
nand \U$53156 ( \53499 , \53490 , \53498 );
xor \U$53157 ( \53500 , \53481 , \53499 );
xor \U$53158 ( \53501 , \51927 , \52249 );
xor \U$53159 ( \53502 , \53501 , \52264 );
xor \U$53160 ( \53503 , \53500 , \53502 );
not \U$53161 ( \53504 , \53503 );
or \U$53162 ( \53505 , \53479 , \53504 );
or \U$53163 ( \53506 , \53503 , \53478 );
nand \U$53164 ( \53507 , \53505 , \53506 );
not \U$53165 ( \53508 , \52717 );
not \U$53166 ( \53509 , \53474 );
not \U$53167 ( \53510 , \53111 );
and \U$53168 ( \53511 , \53509 , \53510 );
and \U$53169 ( \53512 , \53474 , \53111 );
nor \U$53170 ( \53513 , \53511 , \53512 );
not \U$53171 ( \53514 , \53513 );
or \U$53172 ( \53515 , \53508 , \53514 );
or \U$53173 ( \53516 , \53513 , \52717 );
nand \U$53174 ( \53517 , \53515 , \53516 );
not \U$53175 ( \53518 , \53517 );
xnor \U$53176 ( \53519 , \53489 , \53485 );
not \U$53177 ( \53520 , \53519 );
not \U$53178 ( \53521 , \53497 );
and \U$53179 ( \53522 , \53520 , \53521 );
and \U$53180 ( \53523 , \53519 , \53497 );
nor \U$53181 ( \53524 , \53522 , \53523 );
nor \U$53182 ( \53525 , \53518 , \53524 );
and \U$53183 ( \53526 , \53507 , \53525 );
xor \U$53184 ( \53527 , \53525 , \53507 );
not \U$53185 ( \53528 , \53450 );
not \U$53186 ( \53529 , \53141 );
or \U$53187 ( \53530 , \53528 , \53529 );
or \U$53188 ( \53531 , \53141 , \53450 );
nand \U$53189 ( \53532 , \53530 , \53531 );
not \U$53190 ( \53533 , \53532 );
not \U$53191 ( \53534 , \53147 );
and \U$53192 ( \53535 , \53533 , \53534 );
and \U$53193 ( \53536 , \53532 , \53147 );
nor \U$53194 ( \53537 , \53535 , \53536 );
not \U$53195 ( \53538 , \53537 );
and \U$53196 ( \53539 , \8486 , RI9871578_122);
and \U$53197 ( \53540 , RI9871668_124, \8484 );
nor \U$53198 ( \53541 , \53539 , \53540 );
and \U$53199 ( \53542 , \53541 , \8050 );
not \U$53200 ( \53543 , \53541 );
and \U$53201 ( \53544 , \53543 , \8051 );
nor \U$53202 ( \53545 , \53542 , \53544 );
and \U$53203 ( \53546 , \7079 , RI9871398_118);
and \U$53204 ( \53547 , RI9871488_120, \7077 );
nor \U$53205 ( \53548 , \53546 , \53547 );
and \U$53206 ( \53549 , \53548 , \6710 );
not \U$53207 ( \53550 , \53548 );
and \U$53208 ( \53551 , \53550 , \6709 );
nor \U$53209 ( \53552 , \53549 , \53551 );
xor \U$53210 ( \53553 , \53545 , \53552 );
and \U$53211 ( \53554 , \7729 , RI9871758_126);
and \U$53212 ( \53555 , RI9871848_128, \7727 );
nor \U$53213 ( \53556 , \53554 , \53555 );
and \U$53214 ( \53557 , \53556 , \7480 );
not \U$53215 ( \53558 , \53556 );
and \U$53216 ( \53559 , \53558 , \7733 );
nor \U$53217 ( \53560 , \53557 , \53559 );
and \U$53218 ( \53561 , \53553 , \53560 );
and \U$53219 ( \53562 , \53545 , \53552 );
or \U$53220 ( \53563 , \53561 , \53562 );
not \U$53221 ( \53564 , \3918 );
and \U$53222 ( \53565 , \3683 , RI98700d8_78);
and \U$53223 ( \53566 , RI98701c8_80, \3681 );
nor \U$53224 ( \53567 , \53565 , \53566 );
not \U$53225 ( \53568 , \53567 );
or \U$53226 ( \53569 , \53564 , \53568 );
or \U$53227 ( \53570 , \53567 , \3918 );
nand \U$53228 ( \53571 , \53569 , \53570 );
and \U$53229 ( \53572 , \4203 , RI9870fd8_110);
and \U$53230 ( \53573 , RI9870b28_100, \4201 );
nor \U$53231 ( \53574 , \53572 , \53573 );
and \U$53232 ( \53575 , \53574 , \4207 );
not \U$53233 ( \53576 , \53574 );
and \U$53234 ( \53577 , \53576 , \3922 );
nor \U$53235 ( \53578 , \53575 , \53577 );
xor \U$53236 ( \53579 , \53571 , \53578 );
not \U$53237 ( \53580 , \4519 );
and \U$53238 ( \53581 , \4710 , RI9870df8_106);
and \U$53239 ( \53582 , RI9870a38_98, \4708 );
nor \U$53240 ( \53583 , \53581 , \53582 );
not \U$53241 ( \53584 , \53583 );
or \U$53242 ( \53585 , \53580 , \53584 );
or \U$53243 ( \53586 , \53583 , \4521 );
nand \U$53244 ( \53587 , \53585 , \53586 );
and \U$53245 ( \53588 , \53579 , \53587 );
and \U$53246 ( \53589 , \53571 , \53578 );
or \U$53247 ( \53590 , \53588 , \53589 );
xor \U$53248 ( \53591 , \53563 , \53590 );
and \U$53249 ( \53592 , \5318 , RI9870ee8_108);
and \U$53250 ( \53593 , RI9870c18_102, \5316 );
nor \U$53251 ( \53594 , \53592 , \53593 );
and \U$53252 ( \53595 , \53594 , \5052 );
not \U$53253 ( \53596 , \53594 );
and \U$53254 ( \53597 , \53596 , \5322 );
nor \U$53255 ( \53598 , \53595 , \53597 );
and \U$53256 ( \53599 , \5881 , RI98710c8_112);
and \U$53257 ( \53600 , RI9870d08_104, \5879 );
nor \U$53258 ( \53601 , \53599 , \53600 );
and \U$53259 ( \53602 , \53601 , \5594 );
not \U$53260 ( \53603 , \53601 );
and \U$53261 ( \53604 , \53603 , \5885 );
nor \U$53262 ( \53605 , \53602 , \53604 );
xor \U$53263 ( \53606 , \53598 , \53605 );
and \U$53264 ( \53607 , \6453 , RI98712a8_116);
and \U$53265 ( \53608 , RI98711b8_114, \6451 );
nor \U$53266 ( \53609 , \53607 , \53608 );
and \U$53267 ( \53610 , \53609 , \6190 );
not \U$53268 ( \53611 , \53609 );
and \U$53269 ( \53612 , \53611 , \6180 );
nor \U$53270 ( \53613 , \53610 , \53612 );
and \U$53271 ( \53614 , \53606 , \53613 );
and \U$53272 ( \53615 , \53598 , \53605 );
or \U$53273 ( \53616 , \53614 , \53615 );
xor \U$53274 ( \53617 , \53591 , \53616 );
and \U$53275 ( \53618 , \1329 , RI98703a8_84);
and \U$53276 ( \53619 , RI98702b8_82, \1327 );
nor \U$53277 ( \53620 , \53618 , \53619 );
and \U$53278 ( \53621 , \53620 , \1336 );
not \U$53279 ( \53622 , \53620 );
and \U$53280 ( \53623 , \53622 , \1337 );
nor \U$53281 ( \53624 , \53621 , \53623 );
and \U$53282 ( \53625 , \1311 , RI9870768_92);
and \U$53283 ( \53626 , RI9870678_90, \1309 );
nor \U$53284 ( \53627 , \53625 , \53626 );
and \U$53285 ( \53628 , \53627 , \1458 );
not \U$53286 ( \53629 , \53627 );
and \U$53287 ( \53630 , \53629 , \1318 );
nor \U$53288 ( \53631 , \53628 , \53630 );
xor \U$53289 ( \53632 , \53624 , \53631 );
not \U$53290 ( \53633 , \1462 );
and \U$53291 ( \53634 , \2042 , RI9870948_96);
and \U$53292 ( \53635 , RI9870858_94, \2040 );
nor \U$53293 ( \53636 , \53634 , \53635 );
not \U$53294 ( \53637 , \53636 );
or \U$53295 ( \53638 , \53633 , \53637 );
or \U$53296 ( \53639 , \53636 , \1462 );
nand \U$53297 ( \53640 , \53638 , \53639 );
and \U$53298 ( \53641 , \53632 , \53640 );
and \U$53299 ( \53642 , \53624 , \53631 );
or \U$53300 ( \53643 , \53641 , \53642 );
and \U$53301 ( \53644 , \2274 , RI986fb38_66);
and \U$53302 ( \53645 , RI986fc28_68, \2272 );
nor \U$53303 ( \53646 , \53644 , \53645 );
and \U$53304 ( \53647 , \53646 , \2030 );
not \U$53305 ( \53648 , \53646 );
and \U$53306 ( \53649 , \53648 , \2031 );
nor \U$53307 ( \53650 , \53647 , \53649 );
and \U$53308 ( \53651 , \2464 , RI986fe08_72);
and \U$53309 ( \53652 , RI986fd18_70, \2462 );
nor \U$53310 ( \53653 , \53651 , \53652 );
and \U$53311 ( \53654 , \53653 , \2468 );
not \U$53312 ( \53655 , \53653 );
and \U$53313 ( \53656 , \53655 , \2263 );
nor \U$53314 ( \53657 , \53654 , \53656 );
xor \U$53315 ( \53658 , \53650 , \53657 );
not \U$53316 ( \53659 , \2935 );
and \U$53317 ( \53660 , \3254 , RI986ffe8_76);
and \U$53318 ( \53661 , RI986fef8_74, \3252 );
nor \U$53319 ( \53662 , \53660 , \53661 );
not \U$53320 ( \53663 , \53662 );
or \U$53321 ( \53664 , \53659 , \53663 );
or \U$53322 ( \53665 , \53662 , \3406 );
nand \U$53323 ( \53666 , \53664 , \53665 );
and \U$53324 ( \53667 , \53658 , \53666 );
and \U$53325 ( \53668 , \53650 , \53657 );
or \U$53326 ( \53669 , \53667 , \53668 );
xor \U$53327 ( \53670 , \53643 , \53669 );
xor \U$53328 ( \53671 , \53297 , \53302 );
xor \U$53329 ( \53672 , \53671 , \53310 );
xor \U$53330 ( \53673 , \53670 , \53672 );
xor \U$53331 ( \53674 , \53617 , \53673 );
and \U$53332 ( \53675 , \11696 , RI986ec38_34);
and \U$53333 ( \53676 , RI986ed28_36, \11694 );
nor \U$53334 ( \53677 , \53675 , \53676 );
and \U$53335 ( \53678 , \53677 , \10965 );
not \U$53336 ( \53679 , \53677 );
and \U$53337 ( \53680 , \53679 , \11702 );
nor \U$53338 ( \53681 , \53678 , \53680 );
and \U$53339 ( \53682 , \12293 , RI986f0e8_44);
and \U$53340 ( \53683 , RI986eff8_42, \12291 );
nor \U$53341 ( \53684 , \53682 , \53683 );
and \U$53342 ( \53685 , \53684 , \11687 );
not \U$53343 ( \53686 , \53684 );
and \U$53344 ( \53687 , \53686 , \11686 );
nor \U$53345 ( \53688 , \53685 , \53687 );
xor \U$53346 ( \53689 , \53681 , \53688 );
and \U$53347 ( \53690 , \13045 , RI986f2c8_48);
and \U$53348 ( \53691 , RI986f1d8_46, \13043 );
nor \U$53349 ( \53692 , \53690 , \53691 );
and \U$53350 ( \53693 , \53692 , \13047 );
not \U$53351 ( \53694 , \53692 );
and \U$53352 ( \53695 , \53694 , \12619 );
nor \U$53353 ( \53696 , \53693 , \53695 );
and \U$53354 ( \53697 , \53689 , \53696 );
and \U$53355 ( \53698 , \53681 , \53688 );
or \U$53356 ( \53699 , \53697 , \53698 );
and \U$53357 ( \53700 , \13882 , RI986e5a8_20);
and \U$53358 ( \53701 , RI986e4b8_18, \13880 );
nor \U$53359 ( \53702 , \53700 , \53701 );
and \U$53360 ( \53703 , \53702 , \13358 );
not \U$53361 ( \53704 , \53702 );
and \U$53362 ( \53705 , \53704 , \13359 );
nor \U$53363 ( \53706 , \53703 , \53705 );
not \U$53364 ( \53707 , RI9873558_190);
and \U$53365 ( \53708 , \15780 , RI986f868_60);
and \U$53366 ( \53709 , RI986f778_58, RI9873648_192);
nor \U$53367 ( \53710 , \53708 , \53709 );
not \U$53368 ( \53711 , \53710 );
or \U$53369 ( \53712 , \53707 , \53711 );
or \U$53370 ( \53713 , \53710 , RI9873558_190);
nand \U$53371 ( \53714 , \53712 , \53713 );
xor \U$53372 ( \53715 , \53706 , \53714 );
and \U$53373 ( \53716 , \14937 , RI986e788_24);
and \U$53374 ( \53717 , RI986e698_22, \14935 );
nor \U$53375 ( \53718 , \53716 , \53717 );
and \U$53376 ( \53719 , \53718 , \14539 );
not \U$53377 ( \53720 , \53718 );
and \U$53378 ( \53721 , \53720 , \14538 );
nor \U$53379 ( \53722 , \53719 , \53721 );
and \U$53380 ( \53723 , \53715 , \53722 );
and \U$53381 ( \53724 , \53706 , \53714 );
or \U$53382 ( \53725 , \53723 , \53724 );
xor \U$53383 ( \53726 , \53699 , \53725 );
and \U$53384 ( \53727 , \9505 , RI986e968_28);
and \U$53385 ( \53728 , RI986e878_26, \9503 );
nor \U$53386 ( \53729 , \53727 , \53728 );
and \U$53387 ( \53730 , \53729 , \9510 );
not \U$53388 ( \53731 , \53729 );
and \U$53389 ( \53732 , \53731 , \9513 );
nor \U$53390 ( \53733 , \53730 , \53732 );
and \U$53391 ( \53734 , \9237 , RI986eb48_32);
and \U$53392 ( \53735 , RI986ea58_30, \9235 );
nor \U$53393 ( \53736 , \53734 , \53735 );
and \U$53394 ( \53737 , \53736 , \9241 );
not \U$53395 ( \53738 , \53736 );
and \U$53396 ( \53739 , \53738 , \8836 );
nor \U$53397 ( \53740 , \53737 , \53739 );
xor \U$53398 ( \53741 , \53733 , \53740 );
and \U$53399 ( \53742 , \10424 , RI986ef08_40);
and \U$53400 ( \53743 , RI986ee18_38, \10422 );
nor \U$53401 ( \53744 , \53742 , \53743 );
and \U$53402 ( \53745 , \53744 , \9840 );
not \U$53403 ( \53746 , \53744 );
and \U$53404 ( \53747 , \53746 , \10428 );
nor \U$53405 ( \53748 , \53745 , \53747 );
and \U$53406 ( \53749 , \53741 , \53748 );
and \U$53407 ( \53750 , \53733 , \53740 );
or \U$53408 ( \53751 , \53749 , \53750 );
xor \U$53409 ( \53752 , \53726 , \53751 );
and \U$53410 ( \53753 , \53674 , \53752 );
and \U$53411 ( \53754 , \53617 , \53673 );
or \U$53412 ( \53755 , \53753 , \53754 );
xor \U$53413 ( \53756 , \53370 , \53396 );
xor \U$53414 ( \53757 , \53756 , \53422 );
xor \U$53415 ( \53758 , \53215 , \53234 );
xor \U$53416 ( \53759 , \53758 , \53260 );
xor \U$53417 ( \53760 , \53757 , \53759 );
xor \U$53418 ( \53761 , \53289 , \53313 );
xor \U$53419 ( \53762 , \53761 , \53341 );
xor \U$53420 ( \53763 , \53760 , \53762 );
and \U$53421 ( \53764 , \53755 , \53763 );
xnor \U$53422 ( \53765 , \53172 , \53167 );
not \U$53423 ( \53766 , \53765 );
not \U$53424 ( \53767 , \53164 );
and \U$53425 ( \53768 , \53766 , \53767 );
and \U$53426 ( \53769 , \53765 , \53164 );
nor \U$53427 ( \53770 , \53768 , \53769 );
not \U$53428 ( \53771 , \53770 );
not \U$53429 ( \53772 , \53179 );
not \U$53430 ( \53773 , \53185 );
or \U$53431 ( \53774 , \53772 , \53773 );
or \U$53432 ( \53775 , \53179 , \53185 );
nand \U$53433 ( \53776 , \53774 , \53775 );
not \U$53434 ( \53777 , \53776 );
not \U$53435 ( \53778 , \53177 );
and \U$53436 ( \53779 , \53777 , \53778 );
and \U$53437 ( \53780 , \53776 , \53177 );
nor \U$53438 ( \53781 , \53779 , \53780 );
not \U$53439 ( \53782 , \53161 );
not \U$53440 ( \53783 , \53153 );
or \U$53441 ( \53784 , \53782 , \53783 );
or \U$53442 ( \53785 , \53153 , \53161 );
nand \U$53443 ( \53786 , \53784 , \53785 );
not \U$53444 ( \53787 , \53786 );
not \U$53445 ( \53788 , \53155 );
and \U$53446 ( \53789 , \53787 , \53788 );
and \U$53447 ( \53790 , \53786 , \53155 );
nor \U$53448 ( \53791 , \53789 , \53790 );
xor \U$53449 ( \53792 , \53781 , \53791 );
not \U$53450 ( \53793 , \53792 );
or \U$53451 ( \53794 , \53771 , \53793 );
or \U$53452 ( \53795 , \53792 , \53770 );
nand \U$53453 ( \53796 , \53794 , \53795 );
xor \U$53454 ( \53797 , \53757 , \53759 );
xor \U$53455 ( \53798 , \53797 , \53762 );
and \U$53456 ( \53799 , \53796 , \53798 );
and \U$53457 ( \53800 , \53755 , \53796 );
or \U$53458 ( \53801 , \53764 , \53799 , \53800 );
xor \U$53459 ( \53802 , \53681 , \53688 );
xor \U$53460 ( \53803 , \53802 , \53696 );
xor \U$53461 ( \53804 , \53706 , \53714 );
xor \U$53462 ( \53805 , \53804 , \53722 );
and \U$53463 ( \53806 , \53803 , \53805 );
not \U$53464 ( \53807 , \53806 );
xor \U$53465 ( \53808 , \53624 , \53631 );
xor \U$53466 ( \53809 , \53808 , \53640 );
xor \U$53467 ( \53810 , \53571 , \53578 );
xor \U$53468 ( \53811 , \53810 , \53587 );
and \U$53469 ( \53812 , \53809 , \53811 );
xor \U$53470 ( \53813 , \53650 , \53657 );
xor \U$53471 ( \53814 , \53813 , \53666 );
xor \U$53472 ( \53815 , \53571 , \53578 );
xor \U$53473 ( \53816 , \53815 , \53587 );
and \U$53474 ( \53817 , \53814 , \53816 );
and \U$53475 ( \53818 , \53809 , \53814 );
or \U$53476 ( \53819 , \53812 , \53817 , \53818 );
not \U$53477 ( \53820 , \53819 );
or \U$53478 ( \53821 , \53807 , \53820 );
or \U$53479 ( \53822 , \53819 , \53806 );
xor \U$53480 ( \53823 , \53598 , \53605 );
xor \U$53481 ( \53824 , \53823 , \53613 );
xor \U$53482 ( \53825 , \53545 , \53552 );
xor \U$53483 ( \53826 , \53825 , \53560 );
xor \U$53484 ( \53827 , \53824 , \53826 );
xor \U$53485 ( \53828 , \53733 , \53740 );
xor \U$53486 ( \53829 , \53828 , \53748 );
and \U$53487 ( \53830 , \53827 , \53829 );
and \U$53488 ( \53831 , \53824 , \53826 );
or \U$53489 ( \53832 , \53830 , \53831 );
nand \U$53490 ( \53833 , \53822 , \53832 );
nand \U$53491 ( \53834 , \53821 , \53833 );
and \U$53492 ( \53835 , \10424 , RI986e878_26);
and \U$53493 ( \53836 , RI986ef08_40, \10422 );
nor \U$53494 ( \53837 , \53835 , \53836 );
and \U$53495 ( \53838 , \53837 , \9840 );
not \U$53496 ( \53839 , \53837 );
and \U$53497 ( \53840 , \53839 , \10428 );
nor \U$53498 ( \53841 , \53838 , \53840 );
and \U$53499 ( \53842 , \9505 , RI986ea58_30);
and \U$53500 ( \53843 , RI986e968_28, \9503 );
nor \U$53501 ( \53844 , \53842 , \53843 );
and \U$53502 ( \53845 , \53844 , \9510 );
not \U$53503 ( \53846 , \53844 );
and \U$53504 ( \53847 , \53846 , \9513 );
nor \U$53505 ( \53848 , \53845 , \53847 );
xor \U$53506 ( \53849 , \53841 , \53848 );
and \U$53507 ( \53850 , \11696 , RI986ee18_38);
and \U$53508 ( \53851 , RI986ec38_34, \11694 );
nor \U$53509 ( \53852 , \53850 , \53851 );
and \U$53510 ( \53853 , \53852 , \10965 );
not \U$53511 ( \53854 , \53852 );
and \U$53512 ( \53855 , \53854 , \11702 );
nor \U$53513 ( \53856 , \53853 , \53855 );
and \U$53514 ( \53857 , \53849 , \53856 );
and \U$53515 ( \53858 , \53841 , \53848 );
or \U$53516 ( \53859 , \53857 , \53858 );
not \U$53517 ( \53860 , RI9873558_190);
and \U$53518 ( \53861 , \15780 , RI986e698_22);
and \U$53519 ( \53862 , RI986f868_60, RI9873648_192);
nor \U$53520 ( \53863 , \53861 , \53862 );
not \U$53521 ( \53864 , \53863 );
or \U$53522 ( \53865 , \53860 , \53864 );
or \U$53523 ( \53866 , \53863 , RI9873558_190);
nand \U$53524 ( \53867 , \53865 , \53866 );
xor \U$53525 ( \53868 , \53867 , \1301 );
and \U$53526 ( \53869 , \14937 , RI986e4b8_18);
and \U$53527 ( \53870 , RI986e788_24, \14935 );
nor \U$53528 ( \53871 , \53869 , \53870 );
and \U$53529 ( \53872 , \53871 , \14539 );
not \U$53530 ( \53873 , \53871 );
and \U$53531 ( \53874 , \53873 , \14538 );
nor \U$53532 ( \53875 , \53872 , \53874 );
and \U$53533 ( \53876 , \53868 , \53875 );
and \U$53534 ( \53877 , \53867 , \1301 );
or \U$53535 ( \53878 , \53876 , \53877 );
xor \U$53536 ( \53879 , \53859 , \53878 );
and \U$53537 ( \53880 , \12293 , RI986ed28_36);
and \U$53538 ( \53881 , RI986f0e8_44, \12291 );
nor \U$53539 ( \53882 , \53880 , \53881 );
and \U$53540 ( \53883 , \53882 , \11687 );
not \U$53541 ( \53884 , \53882 );
and \U$53542 ( \53885 , \53884 , \11686 );
nor \U$53543 ( \53886 , \53883 , \53885 );
and \U$53544 ( \53887 , \13045 , RI986eff8_42);
and \U$53545 ( \53888 , RI986f2c8_48, \13043 );
nor \U$53546 ( \53889 , \53887 , \53888 );
and \U$53547 ( \53890 , \53889 , \13047 );
not \U$53548 ( \53891 , \53889 );
and \U$53549 ( \53892 , \53891 , \12619 );
nor \U$53550 ( \53893 , \53890 , \53892 );
xor \U$53551 ( \53894 , \53886 , \53893 );
and \U$53552 ( \53895 , \13882 , RI986f1d8_46);
and \U$53553 ( \53896 , RI986e5a8_20, \13880 );
nor \U$53554 ( \53897 , \53895 , \53896 );
and \U$53555 ( \53898 , \53897 , \13358 );
not \U$53556 ( \53899 , \53897 );
and \U$53557 ( \53900 , \53899 , \13359 );
nor \U$53558 ( \53901 , \53898 , \53900 );
and \U$53559 ( \53902 , \53894 , \53901 );
and \U$53560 ( \53903 , \53886 , \53893 );
or \U$53561 ( \53904 , \53902 , \53903 );
and \U$53562 ( \53905 , \53879 , \53904 );
and \U$53563 ( \53906 , \53859 , \53878 );
or \U$53564 ( \53907 , \53905 , \53906 );
and \U$53565 ( \53908 , \2464 , RI986fc28_68);
and \U$53566 ( \53909 , RI986fe08_72, \2462 );
nor \U$53567 ( \53910 , \53908 , \53909 );
and \U$53568 ( \53911 , \53910 , \2468 );
not \U$53569 ( \53912 , \53910 );
and \U$53570 ( \53913 , \53912 , \2263 );
nor \U$53571 ( \53914 , \53911 , \53913 );
not \U$53572 ( \53915 , \2935 );
and \U$53573 ( \53916 , \3254 , RI986fd18_70);
and \U$53574 ( \53917 , RI986ffe8_76, \3252 );
nor \U$53575 ( \53918 , \53916 , \53917 );
not \U$53576 ( \53919 , \53918 );
or \U$53577 ( \53920 , \53915 , \53919 );
or \U$53578 ( \53921 , \53918 , \2935 );
nand \U$53579 ( \53922 , \53920 , \53921 );
xor \U$53580 ( \53923 , \53914 , \53922 );
not \U$53581 ( \53924 , \3412 );
and \U$53582 ( \53925 , \3683 , RI986fef8_74);
and \U$53583 ( \53926 , RI98700d8_78, \3681 );
nor \U$53584 ( \53927 , \53925 , \53926 );
not \U$53585 ( \53928 , \53927 );
or \U$53586 ( \53929 , \53924 , \53928 );
or \U$53587 ( \53930 , \53927 , \3412 );
nand \U$53588 ( \53931 , \53929 , \53930 );
and \U$53589 ( \53932 , \53923 , \53931 );
and \U$53590 ( \53933 , \53914 , \53922 );
or \U$53591 ( \53934 , \53932 , \53933 );
not \U$53592 ( \53935 , \1301 );
and \U$53593 ( \53936 , \1293 , RI9870498_86);
and \U$53594 ( \53937 , RI9870588_88, \1291 );
nor \U$53595 ( \53938 , \53936 , \53937 );
not \U$53596 ( \53939 , \53938 );
or \U$53597 ( \53940 , \53935 , \53939 );
or \U$53598 ( \53941 , \53938 , \1128 );
nand \U$53599 ( \53942 , \53940 , \53941 );
xor \U$53600 ( \53943 , \53934 , \53942 );
not \U$53601 ( \53944 , \2034 );
and \U$53602 ( \53945 , \2042 , RI9870678_90);
and \U$53603 ( \53946 , RI9870948_96, \2040 );
nor \U$53604 ( \53947 , \53945 , \53946 );
not \U$53605 ( \53948 , \53947 );
or \U$53606 ( \53949 , \53944 , \53948 );
or \U$53607 ( \53950 , \53947 , \1462 );
nand \U$53608 ( \53951 , \53949 , \53950 );
and \U$53609 ( \53952 , \1311 , RI98702b8_82);
and \U$53610 ( \53953 , RI9870768_92, \1309 );
nor \U$53611 ( \53954 , \53952 , \53953 );
and \U$53612 ( \53955 , \53954 , \1458 );
not \U$53613 ( \53956 , \53954 );
and \U$53614 ( \53957 , \53956 , \1318 );
nor \U$53615 ( \53958 , \53955 , \53957 );
xor \U$53616 ( \53959 , \53951 , \53958 );
and \U$53617 ( \53960 , \2274 , RI9870858_94);
and \U$53618 ( \53961 , RI986fb38_66, \2272 );
nor \U$53619 ( \53962 , \53960 , \53961 );
and \U$53620 ( \53963 , \53962 , \2030 );
not \U$53621 ( \53964 , \53962 );
and \U$53622 ( \53965 , \53964 , \2031 );
nor \U$53623 ( \53966 , \53963 , \53965 );
and \U$53624 ( \53967 , \53959 , \53966 );
and \U$53625 ( \53968 , \53951 , \53958 );
or \U$53626 ( \53969 , \53967 , \53968 );
and \U$53627 ( \53970 , \53943 , \53969 );
and \U$53628 ( \53971 , \53934 , \53942 );
or \U$53629 ( \53972 , \53970 , \53971 );
xor \U$53630 ( \53973 , \53907 , \53972 );
and \U$53631 ( \53974 , \5881 , RI9870c18_102);
and \U$53632 ( \53975 , RI98710c8_112, \5879 );
nor \U$53633 ( \53976 , \53974 , \53975 );
and \U$53634 ( \53977 , \53976 , \5594 );
not \U$53635 ( \53978 , \53976 );
and \U$53636 ( \53979 , \53978 , \5885 );
nor \U$53637 ( \53980 , \53977 , \53979 );
and \U$53638 ( \53981 , \6453 , RI9870d08_104);
and \U$53639 ( \53982 , RI98712a8_116, \6451 );
nor \U$53640 ( \53983 , \53981 , \53982 );
and \U$53641 ( \53984 , \53983 , \6190 );
not \U$53642 ( \53985 , \53983 );
and \U$53643 ( \53986 , \53985 , \6705 );
nor \U$53644 ( \53987 , \53984 , \53986 );
xor \U$53645 ( \53988 , \53980 , \53987 );
and \U$53646 ( \53989 , \7079 , RI98711b8_114);
and \U$53647 ( \53990 , RI9871398_118, \7077 );
nor \U$53648 ( \53991 , \53989 , \53990 );
and \U$53649 ( \53992 , \53991 , \6710 );
not \U$53650 ( \53993 , \53991 );
and \U$53651 ( \53994 , \53993 , \6709 );
nor \U$53652 ( \53995 , \53992 , \53994 );
and \U$53653 ( \53996 , \53988 , \53995 );
and \U$53654 ( \53997 , \53980 , \53987 );
or \U$53655 ( \53998 , \53996 , \53997 );
and \U$53656 ( \53999 , \4203 , RI98701c8_80);
and \U$53657 ( \54000 , RI9870fd8_110, \4201 );
nor \U$53658 ( \54001 , \53999 , \54000 );
and \U$53659 ( \54002 , \54001 , \4207 );
not \U$53660 ( \54003 , \54001 );
and \U$53661 ( \54004 , \54003 , \3923 );
nor \U$53662 ( \54005 , \54002 , \54004 );
not \U$53663 ( \54006 , \4519 );
and \U$53664 ( \54007 , \4710 , RI9870b28_100);
and \U$53665 ( \54008 , RI9870df8_106, \4708 );
nor \U$53666 ( \54009 , \54007 , \54008 );
not \U$53667 ( \54010 , \54009 );
or \U$53668 ( \54011 , \54006 , \54010 );
or \U$53669 ( \54012 , \54009 , \4521 );
nand \U$53670 ( \54013 , \54011 , \54012 );
xor \U$53671 ( \54014 , \54005 , \54013 );
and \U$53672 ( \54015 , \5318 , RI9870a38_98);
and \U$53673 ( \54016 , RI9870ee8_108, \5316 );
nor \U$53674 ( \54017 , \54015 , \54016 );
and \U$53675 ( \54018 , \54017 , \5052 );
not \U$53676 ( \54019 , \54017 );
and \U$53677 ( \54020 , \54019 , \5322 );
nor \U$53678 ( \54021 , \54018 , \54020 );
and \U$53679 ( \54022 , \54014 , \54021 );
and \U$53680 ( \54023 , \54005 , \54013 );
or \U$53681 ( \54024 , \54022 , \54023 );
xor \U$53682 ( \54025 , \53998 , \54024 );
and \U$53683 ( \54026 , \9237 , RI9871668_124);
and \U$53684 ( \54027 , RI986eb48_32, \9235 );
nor \U$53685 ( \54028 , \54026 , \54027 );
and \U$53686 ( \54029 , \54028 , \9241 );
not \U$53687 ( \54030 , \54028 );
and \U$53688 ( \54031 , \54030 , \8836 );
nor \U$53689 ( \54032 , \54029 , \54031 );
and \U$53690 ( \54033 , \7729 , RI9871488_120);
and \U$53691 ( \54034 , RI9871758_126, \7727 );
nor \U$53692 ( \54035 , \54033 , \54034 );
and \U$53693 ( \54036 , \54035 , \7480 );
not \U$53694 ( \54037 , \54035 );
and \U$53695 ( \54038 , \54037 , \7733 );
nor \U$53696 ( \54039 , \54036 , \54038 );
xor \U$53697 ( \54040 , \54032 , \54039 );
and \U$53698 ( \54041 , \8486 , RI9871848_128);
and \U$53699 ( \54042 , RI9871578_122, \8484 );
nor \U$53700 ( \54043 , \54041 , \54042 );
and \U$53701 ( \54044 , \54043 , \8050 );
not \U$53702 ( \54045 , \54043 );
and \U$53703 ( \54046 , \54045 , \8051 );
nor \U$53704 ( \54047 , \54044 , \54046 );
and \U$53705 ( \54048 , \54040 , \54047 );
and \U$53706 ( \54049 , \54032 , \54039 );
or \U$53707 ( \54050 , \54048 , \54049 );
and \U$53708 ( \54051 , \54025 , \54050 );
and \U$53709 ( \54052 , \53998 , \54024 );
or \U$53710 ( \54053 , \54051 , \54052 );
and \U$53711 ( \54054 , \53973 , \54053 );
and \U$53712 ( \54055 , \53907 , \53972 );
or \U$53713 ( \54056 , \54054 , \54055 );
xor \U$53714 ( \54057 , \53834 , \54056 );
xor \U$53715 ( \54058 , \53242 , \53249 );
xor \U$53716 ( \54059 , \54058 , \53257 );
xor \U$53717 ( \54060 , \53223 , \451 );
xor \U$53718 ( \54061 , \54060 , \53231 );
xor \U$53719 ( \54062 , \54059 , \54061 );
xor \U$53720 ( \54063 , \53270 , \53277 );
xor \U$53721 ( \54064 , \54063 , \53286 );
xor \U$53722 ( \54065 , \53321 , \53329 );
xor \U$53723 ( \54066 , \54065 , \53338 );
xor \U$53724 ( \54067 , \54064 , \54066 );
xor \U$53725 ( \54068 , \53377 , \53384 );
xor \U$53726 ( \54069 , \54068 , \53393 );
xor \U$53727 ( \54070 , \54067 , \54069 );
and \U$53728 ( \54071 , \54062 , \54070 );
xor \U$53729 ( \54072 , \53352 , \53359 );
xor \U$53730 ( \54073 , \54072 , \53367 );
xor \U$53731 ( \54074 , \53404 , \53411 );
xor \U$53732 ( \54075 , \54074 , \53419 );
xor \U$53733 ( \54076 , \53197 , \53204 );
xor \U$53734 ( \54077 , \54076 , \53212 );
xor \U$53735 ( \54078 , \54075 , \54077 );
xor \U$53736 ( \54079 , \54073 , \54078 );
xor \U$53737 ( \54080 , \54064 , \54066 );
xor \U$53738 ( \54081 , \54080 , \54069 );
and \U$53739 ( \54082 , \54079 , \54081 );
and \U$53740 ( \54083 , \54062 , \54079 );
or \U$53741 ( \54084 , \54071 , \54082 , \54083 );
and \U$53742 ( \54085 , \54057 , \54084 );
and \U$53743 ( \54086 , \53834 , \54056 );
or \U$53744 ( \54087 , \54085 , \54086 );
xor \U$53745 ( \54088 , \53801 , \54087 );
xor \U$53746 ( \54089 , \53163 , \53174 );
xor \U$53747 ( \54090 , \54089 , \53187 );
xor \U$53748 ( \54091 , \53263 , \53344 );
xor \U$53749 ( \54092 , \54091 , \53425 );
xor \U$53750 ( \54093 , \53435 , \53441 );
xor \U$53751 ( \54094 , \54093 , \53444 );
xor \U$53752 ( \54095 , \54092 , \54094 );
xor \U$53753 ( \54096 , \54090 , \54095 );
and \U$53754 ( \54097 , \54088 , \54096 );
and \U$53755 ( \54098 , \53801 , \54087 );
or \U$53756 ( \54099 , \54097 , \54098 );
not \U$53757 ( \54100 , \53791 );
not \U$53758 ( \54101 , \53770 );
and \U$53759 ( \54102 , \54100 , \54101 );
and \U$53760 ( \54103 , \53791 , \53770 );
nor \U$53761 ( \54104 , \54103 , \53781 );
nor \U$53762 ( \54105 , \54102 , \54104 );
xor \U$53763 ( \54106 , \53563 , \53590 );
and \U$53764 ( \54107 , \54106 , \53616 );
and \U$53765 ( \54108 , \53563 , \53590 );
or \U$53766 ( \54109 , \54107 , \54108 );
xor \U$53767 ( \54110 , \53699 , \53725 );
and \U$53768 ( \54111 , \54110 , \53751 );
and \U$53769 ( \54112 , \53699 , \53725 );
or \U$53770 ( \54113 , \54111 , \54112 );
xor \U$53771 ( \54114 , \54109 , \54113 );
xor \U$53772 ( \54115 , \53643 , \53669 );
and \U$53773 ( \54116 , \54115 , \53672 );
and \U$53774 ( \54117 , \53643 , \53669 );
or \U$53775 ( \54118 , \54116 , \54117 );
and \U$53776 ( \54119 , \54114 , \54118 );
and \U$53777 ( \54120 , \54109 , \54113 );
nor \U$53778 ( \54121 , \54119 , \54120 );
or \U$53779 ( \54122 , \54105 , \54121 );
not \U$53780 ( \54123 , \54121 );
not \U$53781 ( \54124 , \54105 );
or \U$53782 ( \54125 , \54123 , \54124 );
xor \U$53783 ( \54126 , \53352 , \53359 );
xor \U$53784 ( \54127 , \54126 , \53367 );
and \U$53785 ( \54128 , \54075 , \54127 );
xor \U$53786 ( \54129 , \53352 , \53359 );
xor \U$53787 ( \54130 , \54129 , \53367 );
and \U$53788 ( \54131 , \54077 , \54130 );
and \U$53789 ( \54132 , \54075 , \54077 );
or \U$53790 ( \54133 , \54128 , \54131 , \54132 );
and \U$53791 ( \54134 , \54059 , \54061 );
xor \U$53792 ( \54135 , \54133 , \54134 );
xor \U$53793 ( \54136 , \54064 , \54066 );
and \U$53794 ( \54137 , \54136 , \54069 );
and \U$53795 ( \54138 , \54064 , \54066 );
or \U$53796 ( \54139 , \54137 , \54138 );
and \U$53797 ( \54140 , \54135 , \54139 );
and \U$53798 ( \54141 , \54133 , \54134 );
or \U$53799 ( \54142 , \54140 , \54141 );
nand \U$53800 ( \54143 , \54125 , \54142 );
nand \U$53801 ( \54144 , \54122 , \54143 );
xor \U$53802 ( \54145 , \53163 , \53174 );
xor \U$53803 ( \54146 , \54145 , \53187 );
and \U$53804 ( \54147 , \54092 , \54146 );
xor \U$53805 ( \54148 , \53163 , \53174 );
xor \U$53806 ( \54149 , \54148 , \53187 );
and \U$53807 ( \54150 , \54094 , \54149 );
and \U$53808 ( \54151 , \54092 , \54094 );
or \U$53809 ( \54152 , \54147 , \54150 , \54151 );
xor \U$53810 ( \54153 , \54144 , \54152 );
xor \U$53811 ( \54154 , \53757 , \53759 );
and \U$53812 ( \54155 , \54154 , \53762 );
and \U$53813 ( \54156 , \53757 , \53759 );
or \U$53814 ( \54157 , \54155 , \54156 );
xor \U$53815 ( \54158 , \52948 , \52974 );
xor \U$53816 ( \54159 , \54158 , \53000 );
xor \U$53817 ( \54160 , \54157 , \54159 );
xor \U$53818 ( \54161 , \52876 , \52892 );
xor \U$53819 ( \54162 , \54161 , \52919 );
xor \U$53820 ( \54163 , \53124 , \53129 );
xor \U$53821 ( \54164 , \54162 , \54163 );
and \U$53822 ( \54165 , \54160 , \54164 );
and \U$53823 ( \54166 , \54157 , \54159 );
or \U$53824 ( \54167 , \54165 , \54166 );
xor \U$53825 ( \54168 , \54153 , \54167 );
and \U$53826 ( \54169 , \54099 , \54168 );
not \U$53827 ( \54170 , \53146 );
not \U$53828 ( \54171 , \53143 );
or \U$53829 ( \54172 , \54170 , \54171 );
or \U$53830 ( \54173 , \53143 , \53146 );
nand \U$53831 ( \54174 , \54172 , \54173 );
not \U$53832 ( \54175 , \54174 );
xor \U$53833 ( \54176 , \53122 , \53135 );
xor \U$53834 ( \54177 , \54176 , \53138 );
not \U$53835 ( \54178 , \54177 );
xor \U$53836 ( \54179 , \53190 , \53428 );
xor \U$53837 ( \54180 , \54179 , \53447 );
not \U$53838 ( \54181 , \54180 );
and \U$53839 ( \54182 , \54178 , \54181 );
and \U$53840 ( \54183 , \54177 , \54180 );
nor \U$53841 ( \54184 , \54182 , \54183 );
not \U$53842 ( \54185 , \54184 );
or \U$53843 ( \54186 , \54175 , \54185 );
or \U$53844 ( \54187 , \54184 , \54174 );
nand \U$53845 ( \54188 , \54186 , \54187 );
xor \U$53846 ( \54189 , \54144 , \54152 );
xor \U$53847 ( \54190 , \54189 , \54167 );
and \U$53848 ( \54191 , \54188 , \54190 );
and \U$53849 ( \54192 , \54099 , \54188 );
or \U$53850 ( \54193 , \54169 , \54191 , \54192 );
not \U$53851 ( \54194 , \54193 );
or \U$53852 ( \54195 , \53538 , \54194 );
or \U$53853 ( \54196 , \54193 , \53537 );
nand \U$53854 ( \54197 , \54195 , \54196 );
not \U$53855 ( \54198 , \54197 );
xor \U$53856 ( \54199 , \54144 , \54152 );
and \U$53857 ( \54200 , \54199 , \54167 );
and \U$53858 ( \54201 , \54144 , \54152 );
or \U$53859 ( \54202 , \54200 , \54201 );
not \U$53860 ( \54203 , \54202 );
and \U$53861 ( \54204 , \54180 , \54174 );
not \U$53862 ( \54205 , \54180 );
not \U$53863 ( \54206 , \54174 );
and \U$53864 ( \54207 , \54205 , \54206 );
nor \U$53865 ( \54208 , \54207 , \54177 );
nor \U$53866 ( \54209 , \54204 , \54208 );
not \U$53867 ( \54210 , \54209 );
or \U$53868 ( \54211 , \54203 , \54210 );
or \U$53869 ( \54212 , \54209 , \54202 );
nand \U$53870 ( \54213 , \54211 , \54212 );
not \U$53871 ( \54214 , \54213 );
xnor \U$53872 ( \54215 , \53463 , \53461 );
not \U$53873 ( \54216 , \54215 );
not \U$53874 ( \54217 , \53469 );
and \U$53875 ( \54218 , \54216 , \54217 );
and \U$53876 ( \54219 , \54215 , \53469 );
nor \U$53877 ( \54220 , \54218 , \54219 );
not \U$53878 ( \54221 , \54220 );
and \U$53879 ( \54222 , \54214 , \54221 );
and \U$53880 ( \54223 , \54213 , \54220 );
nor \U$53881 ( \54224 , \54222 , \54223 );
not \U$53882 ( \54225 , \54224 );
and \U$53883 ( \54226 , \54198 , \54225 );
and \U$53884 ( \54227 , \54197 , \54224 );
nor \U$53885 ( \54228 , \54226 , \54227 );
xor \U$53886 ( \54229 , \54144 , \54152 );
xor \U$53887 ( \54230 , \54229 , \54167 );
xor \U$53888 ( \54231 , \54099 , \54188 );
xor \U$53889 ( \54232 , \54230 , \54231 );
not \U$53890 ( \54233 , \54232 );
not \U$53891 ( \54234 , \54121 );
not \U$53892 ( \54235 , \54142 );
or \U$53893 ( \54236 , \54234 , \54235 );
or \U$53894 ( \54237 , \54142 , \54121 );
nand \U$53895 ( \54238 , \54236 , \54237 );
not \U$53896 ( \54239 , \54238 );
not \U$53897 ( \54240 , \54105 );
and \U$53898 ( \54241 , \54239 , \54240 );
and \U$53899 ( \54242 , \54238 , \54105 );
nor \U$53900 ( \54243 , \54241 , \54242 );
not \U$53901 ( \54244 , \54243 );
xor \U$53902 ( \54245 , \53801 , \54087 );
xor \U$53903 ( \54246 , \54245 , \54096 );
nand \U$53904 ( \54247 , \54244 , \54246 );
nand \U$53905 ( \54248 , \54233 , \54247 );
xor \U$53906 ( \54249 , \53841 , \53848 );
xor \U$53907 ( \54250 , \54249 , \53856 );
xor \U$53908 ( \54251 , \53867 , \1301 );
xor \U$53909 ( \54252 , \54251 , \53875 );
and \U$53910 ( \54253 , \54250 , \54252 );
xor \U$53911 ( \54254 , \53886 , \53893 );
xor \U$53912 ( \54255 , \54254 , \53901 );
xor \U$53913 ( \54256 , \53867 , \1301 );
xor \U$53914 ( \54257 , \54256 , \53875 );
and \U$53915 ( \54258 , \54255 , \54257 );
and \U$53916 ( \54259 , \54250 , \54255 );
or \U$53917 ( \54260 , \54253 , \54258 , \54259 );
nand \U$53918 ( \54261 , RI9870498_86, \1291 );
not \U$53919 ( \54262 , \54261 );
not \U$53920 ( \54263 , \1301 );
or \U$53921 ( \54264 , \54262 , \54263 );
or \U$53922 ( \54265 , \1128 , \54261 );
nand \U$53923 ( \54266 , \54264 , \54265 );
xor \U$53924 ( \54267 , \53914 , \53922 );
xor \U$53925 ( \54268 , \54267 , \53931 );
and \U$53926 ( \54269 , \54266 , \54268 );
xor \U$53927 ( \54270 , \53951 , \53958 );
xor \U$53928 ( \54271 , \54270 , \53966 );
xor \U$53929 ( \54272 , \53914 , \53922 );
xor \U$53930 ( \54273 , \54272 , \53931 );
and \U$53931 ( \54274 , \54271 , \54273 );
and \U$53932 ( \54275 , \54266 , \54271 );
or \U$53933 ( \54276 , \54269 , \54274 , \54275 );
xor \U$53934 ( \54277 , \54260 , \54276 );
xor \U$53935 ( \54278 , \54032 , \54039 );
xor \U$53936 ( \54279 , \54278 , \54047 );
xor \U$53937 ( \54280 , \54005 , \54013 );
xor \U$53938 ( \54281 , \54280 , \54021 );
xor \U$53939 ( \54282 , \54279 , \54281 );
xor \U$53940 ( \54283 , \53980 , \53987 );
xor \U$53941 ( \54284 , \54283 , \53995 );
and \U$53942 ( \54285 , \54282 , \54284 );
and \U$53943 ( \54286 , \54279 , \54281 );
or \U$53944 ( \54287 , \54285 , \54286 );
and \U$53945 ( \54288 , \54277 , \54287 );
and \U$53946 ( \54289 , \54260 , \54276 );
or \U$53947 ( \54290 , \54288 , \54289 );
and \U$53948 ( \54291 , \13045 , RI986f0e8_44);
and \U$53949 ( \54292 , RI986eff8_42, \13043 );
nor \U$53950 ( \54293 , \54291 , \54292 );
and \U$53951 ( \54294 , \54293 , \13047 );
not \U$53952 ( \54295 , \54293 );
and \U$53953 ( \54296 , \54295 , \12619 );
nor \U$53954 ( \54297 , \54294 , \54296 );
and \U$53955 ( \54298 , \11696 , RI986ef08_40);
and \U$53956 ( \54299 , RI986ee18_38, \11694 );
nor \U$53957 ( \54300 , \54298 , \54299 );
and \U$53958 ( \54301 , \54300 , \10965 );
not \U$53959 ( \54302 , \54300 );
and \U$53960 ( \54303 , \54302 , \11702 );
nor \U$53961 ( \54304 , \54301 , \54303 );
xor \U$53962 ( \54305 , \54297 , \54304 );
and \U$53963 ( \54306 , \12293 , RI986ec38_34);
and \U$53964 ( \54307 , RI986ed28_36, \12291 );
nor \U$53965 ( \54308 , \54306 , \54307 );
and \U$53966 ( \54309 , \54308 , \11687 );
not \U$53967 ( \54310 , \54308 );
and \U$53968 ( \54311 , \54310 , \11686 );
nor \U$53969 ( \54312 , \54309 , \54311 );
and \U$53970 ( \54313 , \54305 , \54312 );
and \U$53971 ( \54314 , \54297 , \54304 );
or \U$53972 ( \54315 , \54313 , \54314 );
and \U$53973 ( \54316 , \14937 , RI986e5a8_20);
and \U$53974 ( \54317 , RI986e4b8_18, \14935 );
nor \U$53975 ( \54318 , \54316 , \54317 );
and \U$53976 ( \54319 , \54318 , \14539 );
not \U$53977 ( \54320 , \54318 );
and \U$53978 ( \54321 , \54320 , \14538 );
nor \U$53979 ( \54322 , \54319 , \54321 );
not \U$53980 ( \54323 , RI9873558_190);
and \U$53981 ( \54324 , \15780 , RI986e788_24);
and \U$53982 ( \54325 , RI986e698_22, RI9873648_192);
nor \U$53983 ( \54326 , \54324 , \54325 );
not \U$53984 ( \54327 , \54326 );
or \U$53985 ( \54328 , \54323 , \54327 );
or \U$53986 ( \54329 , \54326 , RI9873558_190);
nand \U$53987 ( \54330 , \54328 , \54329 );
xor \U$53988 ( \54331 , \54322 , \54330 );
and \U$53989 ( \54332 , \13882 , RI986f2c8_48);
and \U$53990 ( \54333 , RI986f1d8_46, \13880 );
nor \U$53991 ( \54334 , \54332 , \54333 );
and \U$53992 ( \54335 , \54334 , \13358 );
not \U$53993 ( \54336 , \54334 );
and \U$53994 ( \54337 , \54336 , \13359 );
nor \U$53995 ( \54338 , \54335 , \54337 );
and \U$53996 ( \54339 , \54331 , \54338 );
and \U$53997 ( \54340 , \54322 , \54330 );
or \U$53998 ( \54341 , \54339 , \54340 );
xor \U$53999 ( \54342 , \54315 , \54341 );
and \U$54000 ( \54343 , \9505 , RI986eb48_32);
and \U$54001 ( \54344 , RI986ea58_30, \9503 );
nor \U$54002 ( \54345 , \54343 , \54344 );
and \U$54003 ( \54346 , \54345 , \9510 );
not \U$54004 ( \54347 , \54345 );
and \U$54005 ( \54348 , \54347 , \9513 );
nor \U$54006 ( \54349 , \54346 , \54348 );
and \U$54007 ( \54350 , \9237 , RI9871578_122);
and \U$54008 ( \54351 , RI9871668_124, \9235 );
nor \U$54009 ( \54352 , \54350 , \54351 );
and \U$54010 ( \54353 , \54352 , \9241 );
not \U$54011 ( \54354 , \54352 );
and \U$54012 ( \54355 , \54354 , \8836 );
nor \U$54013 ( \54356 , \54353 , \54355 );
xor \U$54014 ( \54357 , \54349 , \54356 );
and \U$54015 ( \54358 , \10424 , RI986e968_28);
and \U$54016 ( \54359 , RI986e878_26, \10422 );
nor \U$54017 ( \54360 , \54358 , \54359 );
and \U$54018 ( \54361 , \54360 , \9840 );
not \U$54019 ( \54362 , \54360 );
and \U$54020 ( \54363 , \54362 , \10428 );
nor \U$54021 ( \54364 , \54361 , \54363 );
and \U$54022 ( \54365 , \54357 , \54364 );
and \U$54023 ( \54366 , \54349 , \54356 );
or \U$54024 ( \54367 , \54365 , \54366 );
and \U$54025 ( \54368 , \54342 , \54367 );
and \U$54026 ( \54369 , \54315 , \54341 );
or \U$54027 ( \54370 , \54368 , \54369 );
and \U$54028 ( \54371 , \2464 , RI986fb38_66);
and \U$54029 ( \54372 , RI986fc28_68, \2462 );
nor \U$54030 ( \54373 , \54371 , \54372 );
and \U$54031 ( \54374 , \54373 , \2263 );
not \U$54032 ( \54375 , \54373 );
and \U$54033 ( \54376 , \54375 , \2468 );
nor \U$54034 ( \54377 , \54374 , \54376 );
and \U$54035 ( \54378 , \3254 , RI986fe08_72);
and \U$54036 ( \54379 , RI986fd18_70, \3252 );
nor \U$54037 ( \54380 , \54378 , \54379 );
not \U$54038 ( \54381 , \54380 );
not \U$54039 ( \54382 , \3406 );
and \U$54040 ( \54383 , \54381 , \54382 );
and \U$54041 ( \54384 , \54380 , \3406 );
nor \U$54042 ( \54385 , \54383 , \54384 );
xor \U$54043 ( \54386 , \54377 , \54385 );
and \U$54044 ( \54387 , \2274 , RI9870948_96);
and \U$54045 ( \54388 , RI9870858_94, \2272 );
nor \U$54046 ( \54389 , \54387 , \54388 );
and \U$54047 ( \54390 , \54389 , \2031 );
not \U$54048 ( \54391 , \54389 );
and \U$54049 ( \54392 , \54391 , \2030 );
nor \U$54050 ( \54393 , \54390 , \54392 );
and \U$54051 ( \54394 , \54386 , \54393 );
and \U$54052 ( \54395 , \54377 , \54385 );
nor \U$54053 ( \54396 , \54394 , \54395 );
and \U$54054 ( \54397 , \1329 , RI9870588_88);
and \U$54055 ( \54398 , RI98703a8_84, \1327 );
nor \U$54056 ( \54399 , \54397 , \54398 );
and \U$54057 ( \54400 , \54399 , \1336 );
not \U$54058 ( \54401 , \54399 );
and \U$54059 ( \54402 , \54401 , \1337 );
nor \U$54060 ( \54403 , \54400 , \54402 );
xor \U$54061 ( \54404 , \54396 , \54403 );
and \U$54062 ( \54405 , \1311 , RI98703a8_84);
and \U$54063 ( \54406 , RI98702b8_82, \1309 );
nor \U$54064 ( \54407 , \54405 , \54406 );
and \U$54065 ( \54408 , \54407 , \1315 );
not \U$54066 ( \54409 , \54407 );
and \U$54067 ( \54410 , \54409 , \1458 );
nor \U$54068 ( \54411 , \54408 , \54410 );
and \U$54069 ( \54412 , \2042 , RI9870768_92);
and \U$54070 ( \54413 , RI9870678_90, \2040 );
nor \U$54071 ( \54414 , \54412 , \54413 );
not \U$54072 ( \54415 , \54414 );
not \U$54073 ( \54416 , \2034 );
and \U$54074 ( \54417 , \54415 , \54416 );
and \U$54075 ( \54418 , \54414 , \2034 );
nor \U$54076 ( \54419 , \54417 , \54418 );
xor \U$54077 ( \54420 , \54411 , \54419 );
and \U$54078 ( \54421 , \1329 , RI9870498_86);
and \U$54079 ( \54422 , RI9870588_88, \1327 );
nor \U$54080 ( \54423 , \54421 , \54422 );
and \U$54081 ( \54424 , \54423 , \1337 );
not \U$54082 ( \54425 , \54423 );
and \U$54083 ( \54426 , \54425 , \1336 );
nor \U$54084 ( \54427 , \54424 , \54426 );
and \U$54085 ( \54428 , \54420 , \54427 );
and \U$54086 ( \54429 , \54411 , \54419 );
nor \U$54087 ( \54430 , \54428 , \54429 );
and \U$54088 ( \54431 , \54404 , \54430 );
and \U$54089 ( \54432 , \54396 , \54403 );
or \U$54090 ( \54433 , \54431 , \54432 );
xor \U$54091 ( \54434 , \54370 , \54433 );
and \U$54092 ( \54435 , \7079 , RI98712a8_116);
and \U$54093 ( \54436 , RI98711b8_114, \7077 );
nor \U$54094 ( \54437 , \54435 , \54436 );
and \U$54095 ( \54438 , \54437 , \6710 );
not \U$54096 ( \54439 , \54437 );
and \U$54097 ( \54440 , \54439 , \6709 );
nor \U$54098 ( \54441 , \54438 , \54440 );
and \U$54099 ( \54442 , \7729 , RI9871398_118);
and \U$54100 ( \54443 , RI9871488_120, \7727 );
nor \U$54101 ( \54444 , \54442 , \54443 );
and \U$54102 ( \54445 , \54444 , \7480 );
not \U$54103 ( \54446 , \54444 );
and \U$54104 ( \54447 , \54446 , \7733 );
nor \U$54105 ( \54448 , \54445 , \54447 );
xor \U$54106 ( \54449 , \54441 , \54448 );
and \U$54107 ( \54450 , \8486 , RI9871758_126);
and \U$54108 ( \54451 , RI9871848_128, \8484 );
nor \U$54109 ( \54452 , \54450 , \54451 );
and \U$54110 ( \54453 , \54452 , \8050 );
not \U$54111 ( \54454 , \54452 );
and \U$54112 ( \54455 , \54454 , \8051 );
nor \U$54113 ( \54456 , \54453 , \54455 );
and \U$54114 ( \54457 , \54449 , \54456 );
and \U$54115 ( \54458 , \54441 , \54448 );
or \U$54116 ( \54459 , \54457 , \54458 );
and \U$54117 ( \54460 , \3683 , RI986ffe8_76);
and \U$54118 ( \54461 , RI986fef8_74, \3681 );
nor \U$54119 ( \54462 , \54460 , \54461 );
not \U$54120 ( \54463 , \54462 );
not \U$54121 ( \54464 , \3412 );
and \U$54122 ( \54465 , \54463 , \54464 );
and \U$54123 ( \54466 , \54462 , \3918 );
nor \U$54124 ( \54467 , \54465 , \54466 );
and \U$54125 ( \54468 , \4203 , RI98700d8_78);
and \U$54126 ( \54469 , RI98701c8_80, \4201 );
nor \U$54127 ( \54470 , \54468 , \54469 );
and \U$54128 ( \54471 , \54470 , \3922 );
not \U$54129 ( \54472 , \54470 );
and \U$54130 ( \54473 , \54472 , \4207 );
nor \U$54131 ( \54474 , \54471 , \54473 );
or \U$54132 ( \54475 , \54467 , \54474 );
not \U$54133 ( \54476 , \54474 );
not \U$54134 ( \54477 , \54467 );
or \U$54135 ( \54478 , \54476 , \54477 );
not \U$54136 ( \54479 , \4521 );
and \U$54137 ( \54480 , \4710 , RI9870fd8_110);
and \U$54138 ( \54481 , RI9870b28_100, \4708 );
nor \U$54139 ( \54482 , \54480 , \54481 );
not \U$54140 ( \54483 , \54482 );
or \U$54141 ( \54484 , \54479 , \54483 );
or \U$54142 ( \54485 , \54482 , \4521 );
nand \U$54143 ( \54486 , \54484 , \54485 );
nand \U$54144 ( \54487 , \54478 , \54486 );
nand \U$54145 ( \54488 , \54475 , \54487 );
xor \U$54146 ( \54489 , \54459 , \54488 );
and \U$54147 ( \54490 , \6453 , RI98710c8_112);
and \U$54148 ( \54491 , RI9870d08_104, \6451 );
nor \U$54149 ( \54492 , \54490 , \54491 );
and \U$54150 ( \54493 , \54492 , \6190 );
not \U$54151 ( \54494 , \54492 );
and \U$54152 ( \54495 , \54494 , \6180 );
nor \U$54153 ( \54496 , \54493 , \54495 );
and \U$54154 ( \54497 , \5318 , RI9870df8_106);
and \U$54155 ( \54498 , RI9870a38_98, \5316 );
nor \U$54156 ( \54499 , \54497 , \54498 );
and \U$54157 ( \54500 , \54499 , \5052 );
not \U$54158 ( \54501 , \54499 );
and \U$54159 ( \54502 , \54501 , \5322 );
nor \U$54160 ( \54503 , \54500 , \54502 );
xor \U$54161 ( \54504 , \54496 , \54503 );
and \U$54162 ( \54505 , \5881 , RI9870ee8_108);
and \U$54163 ( \54506 , RI9870c18_102, \5879 );
nor \U$54164 ( \54507 , \54505 , \54506 );
and \U$54165 ( \54508 , \54507 , \5594 );
not \U$54166 ( \54509 , \54507 );
and \U$54167 ( \54510 , \54509 , \5885 );
nor \U$54168 ( \54511 , \54508 , \54510 );
and \U$54169 ( \54512 , \54504 , \54511 );
and \U$54170 ( \54513 , \54496 , \54503 );
or \U$54171 ( \54514 , \54512 , \54513 );
and \U$54172 ( \54515 , \54489 , \54514 );
and \U$54173 ( \54516 , \54459 , \54488 );
or \U$54174 ( \54517 , \54515 , \54516 );
and \U$54175 ( \54518 , \54434 , \54517 );
and \U$54176 ( \54519 , \54370 , \54433 );
or \U$54177 ( \54520 , \54518 , \54519 );
xor \U$54178 ( \54521 , \54290 , \54520 );
xor \U$54179 ( \54522 , \53803 , \53805 );
xor \U$54180 ( \54523 , \53824 , \53826 );
xor \U$54181 ( \54524 , \54523 , \53829 );
and \U$54182 ( \54525 , \54522 , \54524 );
xor \U$54183 ( \54526 , \53571 , \53578 );
xor \U$54184 ( \54527 , \54526 , \53587 );
xor \U$54185 ( \54528 , \53809 , \53814 );
xor \U$54186 ( \54529 , \54527 , \54528 );
xor \U$54187 ( \54530 , \53824 , \53826 );
xor \U$54188 ( \54531 , \54530 , \53829 );
and \U$54189 ( \54532 , \54529 , \54531 );
and \U$54190 ( \54533 , \54522 , \54529 );
or \U$54191 ( \54534 , \54525 , \54532 , \54533 );
and \U$54192 ( \54535 , \54521 , \54534 );
and \U$54193 ( \54536 , \54290 , \54520 );
or \U$54194 ( \54537 , \54535 , \54536 );
xor \U$54195 ( \54538 , \54133 , \54134 );
xor \U$54196 ( \54539 , \54538 , \54139 );
xor \U$54197 ( \54540 , \54537 , \54539 );
xor \U$54198 ( \54541 , \53934 , \53942 );
xor \U$54199 ( \54542 , \54541 , \53969 );
xor \U$54200 ( \54543 , \53998 , \54024 );
xor \U$54201 ( \54544 , \54543 , \54050 );
and \U$54202 ( \54545 , \54542 , \54544 );
xor \U$54203 ( \54546 , \53859 , \53878 );
xor \U$54204 ( \54547 , \54546 , \53904 );
xor \U$54205 ( \54548 , \53998 , \54024 );
xor \U$54206 ( \54549 , \54548 , \54050 );
and \U$54207 ( \54550 , \54547 , \54549 );
and \U$54208 ( \54551 , \54542 , \54547 );
or \U$54209 ( \54552 , \54545 , \54550 , \54551 );
xor \U$54210 ( \54553 , \53617 , \53673 );
xor \U$54211 ( \54554 , \54553 , \53752 );
and \U$54212 ( \54555 , \54552 , \54554 );
xor \U$54213 ( \54556 , \54064 , \54066 );
xor \U$54214 ( \54557 , \54556 , \54069 );
xor \U$54215 ( \54558 , \54062 , \54079 );
xor \U$54216 ( \54559 , \54557 , \54558 );
xor \U$54217 ( \54560 , \53617 , \53673 );
xor \U$54218 ( \54561 , \54560 , \53752 );
and \U$54219 ( \54562 , \54559 , \54561 );
and \U$54220 ( \54563 , \54552 , \54559 );
or \U$54221 ( \54564 , \54555 , \54562 , \54563 );
and \U$54222 ( \54565 , \54540 , \54564 );
and \U$54223 ( \54566 , \54537 , \54539 );
or \U$54224 ( \54567 , \54565 , \54566 );
xor \U$54225 ( \54568 , \54157 , \54159 );
xor \U$54226 ( \54569 , \54568 , \54164 );
xor \U$54227 ( \54570 , \54567 , \54569 );
xor \U$54228 ( \54571 , \54109 , \54113 );
xor \U$54229 ( \54572 , \54571 , \54118 );
xor \U$54230 ( \54573 , \53834 , \54056 );
xor \U$54231 ( \54574 , \54573 , \54084 );
and \U$54232 ( \54575 , \54572 , \54574 );
xor \U$54233 ( \54576 , \53757 , \53759 );
xor \U$54234 ( \54577 , \54576 , \53762 );
xor \U$54235 ( \54578 , \53755 , \53796 );
xor \U$54236 ( \54579 , \54577 , \54578 );
xor \U$54237 ( \54580 , \53834 , \54056 );
xor \U$54238 ( \54581 , \54580 , \54084 );
and \U$54239 ( \54582 , \54579 , \54581 );
and \U$54240 ( \54583 , \54572 , \54579 );
or \U$54241 ( \54584 , \54575 , \54582 , \54583 );
and \U$54242 ( \54585 , \54570 , \54584 );
and \U$54243 ( \54586 , \54567 , \54569 );
or \U$54244 ( \54587 , \54585 , \54586 );
and \U$54245 ( \54588 , \54248 , \54587 );
not \U$54246 ( \54589 , \54247 );
and \U$54247 ( \54590 , \54589 , \54232 );
nor \U$54248 ( \54591 , \54588 , \54590 );
or \U$54249 ( \54592 , \54228 , \54591 );
xnor \U$54250 ( \54593 , \54591 , \54228 );
not \U$54251 ( \54594 , \54232 );
not \U$54252 ( \54595 , \54587 );
not \U$54253 ( \54596 , \54247 );
and \U$54254 ( \54597 , \54595 , \54596 );
and \U$54255 ( \54598 , \54587 , \54247 );
nor \U$54256 ( \54599 , \54597 , \54598 );
not \U$54257 ( \54600 , \54599 );
or \U$54258 ( \54601 , \54594 , \54600 );
or \U$54259 ( \54602 , \54599 , \54232 );
nand \U$54260 ( \54603 , \54601 , \54602 );
not \U$54261 ( \54604 , \54243 );
not \U$54262 ( \54605 , \54246 );
or \U$54263 ( \54606 , \54604 , \54605 );
or \U$54264 ( \54607 , \54246 , \54243 );
nand \U$54265 ( \54608 , \54606 , \54607 );
not \U$54266 ( \54609 , \54608 );
xor \U$54267 ( \54610 , \54567 , \54569 );
xor \U$54268 ( \54611 , \54610 , \54584 );
not \U$54269 ( \54612 , \54611 );
or \U$54270 ( \54613 , \54609 , \54612 );
or \U$54271 ( \54614 , \54611 , \54608 );
xor \U$54272 ( \54615 , \53998 , \54024 );
xor \U$54273 ( \54616 , \54615 , \54050 );
xor \U$54274 ( \54617 , \54542 , \54547 );
xor \U$54275 ( \54618 , \54616 , \54617 );
xor \U$54276 ( \54619 , \54260 , \54276 );
xor \U$54277 ( \54620 , \54619 , \54287 );
and \U$54278 ( \54621 , \54618 , \54620 );
xor \U$54279 ( \54622 , \53824 , \53826 );
xor \U$54280 ( \54623 , \54622 , \53829 );
xor \U$54281 ( \54624 , \54522 , \54529 );
xor \U$54282 ( \54625 , \54623 , \54624 );
xor \U$54283 ( \54626 , \54260 , \54276 );
xor \U$54284 ( \54627 , \54626 , \54287 );
and \U$54285 ( \54628 , \54625 , \54627 );
and \U$54286 ( \54629 , \54618 , \54625 );
or \U$54287 ( \54630 , \54621 , \54628 , \54629 );
not \U$54288 ( \54631 , \54630 );
xnor \U$54289 ( \54632 , \53832 , \53819 );
not \U$54290 ( \54633 , \54632 );
not \U$54291 ( \54634 , \53806 );
and \U$54292 ( \54635 , \54633 , \54634 );
and \U$54293 ( \54636 , \54632 , \53806 );
nor \U$54294 ( \54637 , \54635 , \54636 );
or \U$54295 ( \54638 , \54631 , \54637 );
not \U$54296 ( \54639 , \54637 );
not \U$54297 ( \54640 , \54631 );
or \U$54298 ( \54641 , \54639 , \54640 );
xor \U$54299 ( \54642 , \54441 , \54448 );
xor \U$54300 ( \54643 , \54642 , \54456 );
xor \U$54301 ( \54644 , \54297 , \54304 );
xor \U$54302 ( \54645 , \54644 , \54312 );
and \U$54303 ( \54646 , \54643 , \54645 );
xor \U$54304 ( \54647 , \54349 , \54356 );
xor \U$54305 ( \54648 , \54647 , \54364 );
xor \U$54306 ( \54649 , \54297 , \54304 );
xor \U$54307 ( \54650 , \54649 , \54312 );
and \U$54308 ( \54651 , \54648 , \54650 );
and \U$54309 ( \54652 , \54643 , \54648 );
or \U$54310 ( \54653 , \54646 , \54651 , \54652 );
xor \U$54311 ( \54654 , \54377 , \54385 );
xor \U$54312 ( \54655 , \54654 , \54393 );
not \U$54313 ( \54656 , \54474 );
not \U$54314 ( \54657 , \54486 );
or \U$54315 ( \54658 , \54656 , \54657 );
or \U$54316 ( \54659 , \54474 , \54486 );
nand \U$54317 ( \54660 , \54658 , \54659 );
not \U$54318 ( \54661 , \54660 );
not \U$54319 ( \54662 , \54467 );
and \U$54320 ( \54663 , \54661 , \54662 );
and \U$54321 ( \54664 , \54660 , \54467 );
nor \U$54322 ( \54665 , \54663 , \54664 );
or \U$54323 ( \54666 , \54655 , \54665 );
not \U$54324 ( \54667 , \54665 );
not \U$54325 ( \54668 , \54655 );
or \U$54326 ( \54669 , \54667 , \54668 );
xor \U$54327 ( \54670 , \54496 , \54503 );
xor \U$54328 ( \54671 , \54670 , \54511 );
nand \U$54329 ( \54672 , \54669 , \54671 );
nand \U$54330 ( \54673 , \54666 , \54672 );
xor \U$54331 ( \54674 , \54653 , \54673 );
xor \U$54332 ( \54675 , \53867 , \1301 );
xor \U$54333 ( \54676 , \54675 , \53875 );
xor \U$54334 ( \54677 , \54250 , \54255 );
xor \U$54335 ( \54678 , \54676 , \54677 );
and \U$54336 ( \54679 , \54674 , \54678 );
and \U$54337 ( \54680 , \54653 , \54673 );
or \U$54338 ( \54681 , \54679 , \54680 );
and \U$54339 ( \54682 , \10424 , RI986ea58_30);
and \U$54340 ( \54683 , RI986e968_28, \10422 );
nor \U$54341 ( \54684 , \54682 , \54683 );
and \U$54342 ( \54685 , \54684 , \10428 );
not \U$54343 ( \54686 , \54684 );
and \U$54344 ( \54687 , \54686 , \9840 );
nor \U$54345 ( \54688 , \54685 , \54687 );
and \U$54346 ( \54689 , \9505 , RI9871668_124);
and \U$54347 ( \54690 , RI986eb48_32, \9503 );
nor \U$54348 ( \54691 , \54689 , \54690 );
and \U$54349 ( \54692 , \54691 , \9513 );
not \U$54350 ( \54693 , \54691 );
and \U$54351 ( \54694 , \54693 , \9510 );
nor \U$54352 ( \54695 , \54692 , \54694 );
xor \U$54353 ( \54696 , \54688 , \54695 );
and \U$54354 ( \54697 , \11696 , RI986e878_26);
and \U$54355 ( \54698 , RI986ef08_40, \11694 );
nor \U$54356 ( \54699 , \54697 , \54698 );
and \U$54357 ( \54700 , \54699 , \11702 );
not \U$54358 ( \54701 , \54699 );
and \U$54359 ( \54702 , \54701 , \10965 );
nor \U$54360 ( \54703 , \54700 , \54702 );
and \U$54361 ( \54704 , \54696 , \54703 );
and \U$54362 ( \54705 , \54688 , \54695 );
or \U$54363 ( \54706 , \54704 , \54705 );
not \U$54364 ( \54707 , RI9873558_190);
and \U$54365 ( \54708 , \15780 , RI986e4b8_18);
and \U$54366 ( \54709 , RI986e788_24, RI9873648_192);
nor \U$54367 ( \54710 , \54708 , \54709 );
not \U$54368 ( \54711 , \54710 );
or \U$54369 ( \54712 , \54707 , \54711 );
or \U$54370 ( \54713 , \54710 , RI9873558_190);
nand \U$54371 ( \54714 , \54712 , \54713 );
and \U$54372 ( \54715 , \54714 , \1337 );
not \U$54373 ( \54716 , \54714 );
not \U$54374 ( \54717 , \1337 );
and \U$54375 ( \54718 , \54716 , \54717 );
and \U$54376 ( \54719 , \14937 , RI986f1d8_46);
and \U$54377 ( \54720 , RI986e5a8_20, \14935 );
nor \U$54378 ( \54721 , \54719 , \54720 );
and \U$54379 ( \54722 , \54721 , \14538 );
not \U$54380 ( \54723 , \54721 );
and \U$54381 ( \54724 , \54723 , \14539 );
nor \U$54382 ( \54725 , \54722 , \54724 );
nor \U$54383 ( \54726 , \54718 , \54725 );
nor \U$54384 ( \54727 , \54715 , \54726 );
xor \U$54385 ( \54728 , \54706 , \54727 );
and \U$54386 ( \54729 , \13045 , RI986ed28_36);
and \U$54387 ( \54730 , RI986f0e8_44, \13043 );
nor \U$54388 ( \54731 , \54729 , \54730 );
and \U$54389 ( \54732 , \54731 , \12619 );
not \U$54390 ( \54733 , \54731 );
and \U$54391 ( \54734 , \54733 , \13047 );
nor \U$54392 ( \54735 , \54732 , \54734 );
and \U$54393 ( \54736 , \12293 , RI986ee18_38);
and \U$54394 ( \54737 , RI986ec38_34, \12291 );
nor \U$54395 ( \54738 , \54736 , \54737 );
and \U$54396 ( \54739 , \54738 , \11686 );
not \U$54397 ( \54740 , \54738 );
and \U$54398 ( \54741 , \54740 , \11687 );
nor \U$54399 ( \54742 , \54739 , \54741 );
xor \U$54400 ( \54743 , \54735 , \54742 );
and \U$54401 ( \54744 , \13882 , RI986eff8_42);
and \U$54402 ( \54745 , RI986f2c8_48, \13880 );
nor \U$54403 ( \54746 , \54744 , \54745 );
and \U$54404 ( \54747 , \54746 , \13359 );
not \U$54405 ( \54748 , \54746 );
and \U$54406 ( \54749 , \54748 , \13358 );
nor \U$54407 ( \54750 , \54747 , \54749 );
and \U$54408 ( \54751 , \54743 , \54750 );
and \U$54409 ( \54752 , \54735 , \54742 );
or \U$54410 ( \54753 , \54751 , \54752 );
and \U$54411 ( \54754 , \54728 , \54753 );
and \U$54412 ( \54755 , \54706 , \54727 );
or \U$54413 ( \54756 , \54754 , \54755 );
and \U$54414 ( \54757 , \7729 , RI98711b8_114);
and \U$54415 ( \54758 , RI9871398_118, \7727 );
nor \U$54416 ( \54759 , \54757 , \54758 );
and \U$54417 ( \54760 , \54759 , \7733 );
not \U$54418 ( \54761 , \54759 );
and \U$54419 ( \54762 , \54761 , \7480 );
nor \U$54420 ( \54763 , \54760 , \54762 );
not \U$54421 ( \54764 , \54763 );
and \U$54422 ( \54765 , \9237 , RI9871848_128);
and \U$54423 ( \54766 , RI9871578_122, \9235 );
nor \U$54424 ( \54767 , \54765 , \54766 );
and \U$54425 ( \54768 , \54767 , \8836 );
not \U$54426 ( \54769 , \54767 );
and \U$54427 ( \54770 , \54769 , \9241 );
nor \U$54428 ( \54771 , \54768 , \54770 );
not \U$54429 ( \54772 , \54771 );
and \U$54430 ( \54773 , \54764 , \54772 );
and \U$54431 ( \54774 , \54771 , \54763 );
and \U$54432 ( \54775 , \8486 , RI9871488_120);
and \U$54433 ( \54776 , RI9871758_126, \8484 );
nor \U$54434 ( \54777 , \54775 , \54776 );
and \U$54435 ( \54778 , \54777 , \8051 );
not \U$54436 ( \54779 , \54777 );
and \U$54437 ( \54780 , \54779 , \8050 );
nor \U$54438 ( \54781 , \54778 , \54780 );
nor \U$54439 ( \54782 , \54774 , \54781 );
nor \U$54440 ( \54783 , \54773 , \54782 );
and \U$54441 ( \54784 , \7079 , RI9870d08_104);
and \U$54442 ( \54785 , RI98712a8_116, \7077 );
nor \U$54443 ( \54786 , \54784 , \54785 );
and \U$54444 ( \54787 , \54786 , \6709 );
not \U$54445 ( \54788 , \54786 );
and \U$54446 ( \54789 , \54788 , \6710 );
nor \U$54447 ( \54790 , \54787 , \54789 );
and \U$54448 ( \54791 , \5881 , RI9870a38_98);
and \U$54449 ( \54792 , RI9870ee8_108, \5879 );
nor \U$54450 ( \54793 , \54791 , \54792 );
and \U$54451 ( \54794 , \54793 , \5885 );
not \U$54452 ( \54795 , \54793 );
and \U$54453 ( \54796 , \54795 , \5594 );
nor \U$54454 ( \54797 , \54794 , \54796 );
xor \U$54455 ( \54798 , \54790 , \54797 );
and \U$54456 ( \54799 , \6453 , RI9870c18_102);
and \U$54457 ( \54800 , RI98710c8_112, \6451 );
nor \U$54458 ( \54801 , \54799 , \54800 );
and \U$54459 ( \54802 , \54801 , \6180 );
not \U$54460 ( \54803 , \54801 );
and \U$54461 ( \54804 , \54803 , \6190 );
nor \U$54462 ( \54805 , \54802 , \54804 );
and \U$54463 ( \54806 , \54798 , \54805 );
and \U$54464 ( \54807 , \54790 , \54797 );
or \U$54465 ( \54808 , \54806 , \54807 );
xor \U$54466 ( \54809 , \54783 , \54808 );
and \U$54467 ( \54810 , \4710 , RI98701c8_80);
and \U$54468 ( \54811 , RI9870fd8_110, \4708 );
nor \U$54469 ( \54812 , \54810 , \54811 );
not \U$54470 ( \54813 , \54812 );
not \U$54471 ( \54814 , \4519 );
and \U$54472 ( \54815 , \54813 , \54814 );
and \U$54473 ( \54816 , \54812 , \4519 );
nor \U$54474 ( \54817 , \54815 , \54816 );
and \U$54475 ( \54818 , \4203 , RI986fef8_74);
and \U$54476 ( \54819 , RI98700d8_78, \4201 );
nor \U$54477 ( \54820 , \54818 , \54819 );
and \U$54478 ( \54821 , \54820 , \3923 );
not \U$54479 ( \54822 , \54820 );
and \U$54480 ( \54823 , \54822 , \4207 );
nor \U$54481 ( \54824 , \54821 , \54823 );
xor \U$54482 ( \54825 , \54817 , \54824 );
and \U$54483 ( \54826 , \5318 , RI9870b28_100);
and \U$54484 ( \54827 , RI9870df8_106, \5316 );
nor \U$54485 ( \54828 , \54826 , \54827 );
and \U$54486 ( \54829 , \54828 , \5322 );
not \U$54487 ( \54830 , \54828 );
and \U$54488 ( \54831 , \54830 , \5052 );
nor \U$54489 ( \54832 , \54829 , \54831 );
and \U$54490 ( \54833 , \54825 , \54832 );
and \U$54491 ( \54834 , \54817 , \54824 );
or \U$54492 ( \54835 , \54833 , \54834 );
and \U$54493 ( \54836 , \54809 , \54835 );
and \U$54494 ( \54837 , \54783 , \54808 );
or \U$54495 ( \54838 , \54836 , \54837 );
xor \U$54496 ( \54839 , \54756 , \54838 );
and \U$54497 ( \54840 , \2274 , RI9870678_90);
and \U$54498 ( \54841 , RI9870948_96, \2272 );
nor \U$54499 ( \54842 , \54840 , \54841 );
and \U$54500 ( \54843 , \54842 , \2031 );
not \U$54501 ( \54844 , \54842 );
and \U$54502 ( \54845 , \54844 , \2030 );
nor \U$54503 ( \54846 , \54843 , \54845 );
and \U$54504 ( \54847 , \1311 , RI9870588_88);
and \U$54505 ( \54848 , RI98703a8_84, \1309 );
nor \U$54506 ( \54849 , \54847 , \54848 );
and \U$54507 ( \54850 , \54849 , \1315 );
not \U$54508 ( \54851 , \54849 );
and \U$54509 ( \54852 , \54851 , \1319 );
nor \U$54510 ( \54853 , \54850 , \54852 );
xor \U$54511 ( \54854 , \54846 , \54853 );
and \U$54512 ( \54855 , \2042 , RI98702b8_82);
and \U$54513 ( \54856 , RI9870768_92, \2040 );
nor \U$54514 ( \54857 , \54855 , \54856 );
not \U$54515 ( \54858 , \54857 );
not \U$54516 ( \54859 , \1462 );
and \U$54517 ( \54860 , \54858 , \54859 );
and \U$54518 ( \54861 , \54857 , \1462 );
nor \U$54519 ( \54862 , \54860 , \54861 );
and \U$54520 ( \54863 , \54854 , \54862 );
and \U$54521 ( \54864 , \54846 , \54853 );
or \U$54522 ( \54865 , \54863 , \54864 );
and \U$54523 ( \54866 , \2464 , RI9870858_94);
and \U$54524 ( \54867 , RI986fb38_66, \2462 );
nor \U$54525 ( \54868 , \54866 , \54867 );
and \U$54526 ( \54869 , \54868 , \2263 );
not \U$54527 ( \54870 , \54868 );
and \U$54528 ( \54871 , \54870 , \2468 );
nor \U$54529 ( \54872 , \54869 , \54871 );
and \U$54530 ( \54873 , \3254 , RI986fc28_68);
and \U$54531 ( \54874 , RI986fe08_72, \3252 );
nor \U$54532 ( \54875 , \54873 , \54874 );
not \U$54533 ( \54876 , \54875 );
not \U$54534 ( \54877 , \2935 );
and \U$54535 ( \54878 , \54876 , \54877 );
and \U$54536 ( \54879 , \54875 , \2935 );
nor \U$54537 ( \54880 , \54878 , \54879 );
xor \U$54538 ( \54881 , \54872 , \54880 );
and \U$54539 ( \54882 , \3683 , RI986fd18_70);
and \U$54540 ( \54883 , RI986ffe8_76, \3681 );
nor \U$54541 ( \54884 , \54882 , \54883 );
not \U$54542 ( \54885 , \54884 );
not \U$54543 ( \54886 , \3918 );
and \U$54544 ( \54887 , \54885 , \54886 );
and \U$54545 ( \54888 , \54884 , \3412 );
nor \U$54546 ( \54889 , \54887 , \54888 );
and \U$54547 ( \54890 , \54881 , \54889 );
and \U$54548 ( \54891 , \54872 , \54880 );
or \U$54549 ( \54892 , \54890 , \54891 );
xor \U$54550 ( \54893 , \54865 , \54892 );
xor \U$54551 ( \54894 , \54411 , \54419 );
xor \U$54552 ( \54895 , \54894 , \54427 );
and \U$54553 ( \54896 , \54893 , \54895 );
and \U$54554 ( \54897 , \54865 , \54892 );
or \U$54555 ( \54898 , \54896 , \54897 );
and \U$54556 ( \54899 , \54839 , \54898 );
and \U$54557 ( \54900 , \54756 , \54838 );
nor \U$54558 ( \54901 , \54899 , \54900 );
xor \U$54559 ( \54902 , \54681 , \54901 );
xor \U$54560 ( \54903 , \54396 , \54403 );
xor \U$54561 ( \54904 , \54903 , \54430 );
xor \U$54562 ( \54905 , \54279 , \54281 );
xor \U$54563 ( \54906 , \54905 , \54284 );
and \U$54564 ( \54907 , \54904 , \54906 );
xor \U$54565 ( \54908 , \53914 , \53922 );
xor \U$54566 ( \54909 , \54908 , \53931 );
xor \U$54567 ( \54910 , \54266 , \54271 );
xor \U$54568 ( \54911 , \54909 , \54910 );
xor \U$54569 ( \54912 , \54279 , \54281 );
xor \U$54570 ( \54913 , \54912 , \54284 );
and \U$54571 ( \54914 , \54911 , \54913 );
and \U$54572 ( \54915 , \54904 , \54911 );
or \U$54573 ( \54916 , \54907 , \54914 , \54915 );
and \U$54574 ( \54917 , \54902 , \54916 );
and \U$54575 ( \54918 , \54681 , \54901 );
or \U$54576 ( \54919 , \54917 , \54918 );
nand \U$54577 ( \54920 , \54641 , \54919 );
nand \U$54578 ( \54921 , \54638 , \54920 );
xor \U$54579 ( \54922 , \53907 , \53972 );
xor \U$54580 ( \54923 , \54922 , \54053 );
xor \U$54581 ( \54924 , \54290 , \54520 );
xor \U$54582 ( \54925 , \54924 , \54534 );
and \U$54583 ( \54926 , \54923 , \54925 );
xor \U$54584 ( \54927 , \53617 , \53673 );
xor \U$54585 ( \54928 , \54927 , \53752 );
xor \U$54586 ( \54929 , \54552 , \54559 );
xor \U$54587 ( \54930 , \54928 , \54929 );
xor \U$54588 ( \54931 , \54290 , \54520 );
xor \U$54589 ( \54932 , \54931 , \54534 );
and \U$54590 ( \54933 , \54930 , \54932 );
and \U$54591 ( \54934 , \54923 , \54930 );
or \U$54592 ( \54935 , \54926 , \54933 , \54934 );
xor \U$54593 ( \54936 , \54921 , \54935 );
xor \U$54594 ( \54937 , \53834 , \54056 );
xor \U$54595 ( \54938 , \54937 , \54084 );
xor \U$54596 ( \54939 , \54572 , \54579 );
xor \U$54597 ( \54940 , \54938 , \54939 );
and \U$54598 ( \54941 , \54936 , \54940 );
and \U$54599 ( \54942 , \54921 , \54935 );
or \U$54600 ( \54943 , \54941 , \54942 );
nand \U$54601 ( \54944 , \54614 , \54943 );
nand \U$54602 ( \54945 , \54613 , \54944 );
and \U$54603 ( \54946 , \54603 , \54945 );
xor \U$54604 ( \54947 , \54945 , \54603 );
xor \U$54605 ( \54948 , \54756 , \54838 );
xor \U$54606 ( \54949 , \54948 , \54898 );
not \U$54607 ( \54950 , \54949 );
xor \U$54608 ( \54951 , \54653 , \54673 );
xor \U$54609 ( \54952 , \54951 , \54678 );
not \U$54610 ( \54953 , \54952 );
or \U$54611 ( \54954 , \54950 , \54953 );
or \U$54612 ( \54955 , \54952 , \54949 );
nand \U$54613 ( \54956 , \54954 , \54955 );
not \U$54614 ( \54957 , \54956 );
xor \U$54615 ( \54958 , \54688 , \54695 );
xor \U$54616 ( \54959 , \54958 , \54703 );
xor \U$54617 ( \54960 , \54735 , \54742 );
xor \U$54618 ( \54961 , \54960 , \54750 );
or \U$54619 ( \54962 , \54959 , \54961 );
not \U$54620 ( \54963 , \54961 );
not \U$54621 ( \54964 , \54959 );
or \U$54622 ( \54965 , \54963 , \54964 );
not \U$54623 ( \54966 , \54763 );
xor \U$54624 ( \54967 , \54781 , \54771 );
not \U$54625 ( \54968 , \54967 );
or \U$54626 ( \54969 , \54966 , \54968 );
or \U$54627 ( \54970 , \54967 , \54763 );
nand \U$54628 ( \54971 , \54969 , \54970 );
nand \U$54629 ( \54972 , \54965 , \54971 );
nand \U$54630 ( \54973 , \54962 , \54972 );
xor \U$54631 ( \54974 , \54322 , \54330 );
xor \U$54632 ( \54975 , \54974 , \54338 );
xor \U$54633 ( \54976 , \54973 , \54975 );
xor \U$54634 ( \54977 , \54872 , \54880 );
xor \U$54635 ( \54978 , \54977 , \54889 );
xor \U$54636 ( \54979 , \54817 , \54824 );
xor \U$54637 ( \54980 , \54979 , \54832 );
xor \U$54638 ( \54981 , \54978 , \54980 );
xor \U$54639 ( \54982 , \54790 , \54797 );
xor \U$54640 ( \54983 , \54982 , \54805 );
and \U$54641 ( \54984 , \54981 , \54983 );
and \U$54642 ( \54985 , \54978 , \54980 );
nor \U$54643 ( \54986 , \54984 , \54985 );
and \U$54644 ( \54987 , \54976 , \54986 );
and \U$54645 ( \54988 , \54973 , \54975 );
or \U$54646 ( \54989 , \54987 , \54988 );
and \U$54647 ( \54990 , \2274 , RI9870768_92);
and \U$54648 ( \54991 , RI9870678_90, \2272 );
nor \U$54649 ( \54992 , \54990 , \54991 );
and \U$54650 ( \54993 , \54992 , \2031 );
not \U$54651 ( \54994 , \54992 );
and \U$54652 ( \54995 , \54994 , \2030 );
nor \U$54653 ( \54996 , \54993 , \54995 );
not \U$54654 ( \54997 , \54996 );
and \U$54655 ( \54998 , \3254 , RI986fb38_66);
and \U$54656 ( \54999 , RI986fc28_68, \3252 );
nor \U$54657 ( \55000 , \54998 , \54999 );
not \U$54658 ( \55001 , \55000 );
not \U$54659 ( \55002 , \3406 );
and \U$54660 ( \55003 , \55001 , \55002 );
and \U$54661 ( \55004 , \55000 , \2935 );
nor \U$54662 ( \55005 , \55003 , \55004 );
not \U$54663 ( \55006 , \55005 );
and \U$54664 ( \55007 , \54997 , \55006 );
and \U$54665 ( \55008 , \55005 , \54996 );
and \U$54666 ( \55009 , \2464 , RI9870948_96);
and \U$54667 ( \55010 , RI9870858_94, \2462 );
nor \U$54668 ( \55011 , \55009 , \55010 );
and \U$54669 ( \55012 , \55011 , \2263 );
not \U$54670 ( \55013 , \55011 );
and \U$54671 ( \55014 , \55013 , \2468 );
nor \U$54672 ( \55015 , \55012 , \55014 );
nor \U$54673 ( \55016 , \55008 , \55015 );
nor \U$54674 ( \55017 , \55007 , \55016 );
nand \U$54675 ( \55018 , RI9870498_86, \1327 );
and \U$54676 ( \55019 , \55018 , \1337 );
not \U$54677 ( \55020 , \55018 );
and \U$54678 ( \55021 , \55020 , \1336 );
nor \U$54679 ( \55022 , \55019 , \55021 );
xor \U$54680 ( \55023 , \55017 , \55022 );
xor \U$54681 ( \55024 , \54846 , \54853 );
xor \U$54682 ( \55025 , \55024 , \54862 );
and \U$54683 ( \55026 , \55023 , \55025 );
and \U$54684 ( \55027 , \55017 , \55022 );
or \U$54685 ( \55028 , \55026 , \55027 );
and \U$54686 ( \55029 , \7079 , RI98710c8_112);
and \U$54687 ( \55030 , RI9870d08_104, \7077 );
nor \U$54688 ( \55031 , \55029 , \55030 );
and \U$54689 ( \55032 , \55031 , \6710 );
not \U$54690 ( \55033 , \55031 );
and \U$54691 ( \55034 , \55033 , \6709 );
nor \U$54692 ( \55035 , \55032 , \55034 );
and \U$54693 ( \55036 , \7729 , RI98712a8_116);
and \U$54694 ( \55037 , RI98711b8_114, \7727 );
nor \U$54695 ( \55038 , \55036 , \55037 );
and \U$54696 ( \55039 , \55038 , \7480 );
not \U$54697 ( \55040 , \55038 );
and \U$54698 ( \55041 , \55040 , \7733 );
nor \U$54699 ( \55042 , \55039 , \55041 );
xor \U$54700 ( \55043 , \55035 , \55042 );
and \U$54701 ( \55044 , \8486 , RI9871398_118);
and \U$54702 ( \55045 , RI9871488_120, \8484 );
nor \U$54703 ( \55046 , \55044 , \55045 );
and \U$54704 ( \55047 , \55046 , \8050 );
not \U$54705 ( \55048 , \55046 );
and \U$54706 ( \55049 , \55048 , \8051 );
nor \U$54707 ( \55050 , \55047 , \55049 );
and \U$54708 ( \55051 , \55043 , \55050 );
and \U$54709 ( \55052 , \55035 , \55042 );
or \U$54710 ( \55053 , \55051 , \55052 );
and \U$54711 ( \55054 , \5881 , RI9870df8_106);
and \U$54712 ( \55055 , RI9870a38_98, \5879 );
nor \U$54713 ( \55056 , \55054 , \55055 );
and \U$54714 ( \55057 , \55056 , \5885 );
not \U$54715 ( \55058 , \55056 );
and \U$54716 ( \55059 , \55058 , \5594 );
nor \U$54717 ( \55060 , \55057 , \55059 );
and \U$54718 ( \55061 , \6453 , RI9870ee8_108);
and \U$54719 ( \55062 , RI9870c18_102, \6451 );
nor \U$54720 ( \55063 , \55061 , \55062 );
and \U$54721 ( \55064 , \55063 , \6705 );
not \U$54722 ( \55065 , \55063 );
and \U$54723 ( \55066 , \55065 , \6190 );
nor \U$54724 ( \55067 , \55064 , \55066 );
xor \U$54725 ( \55068 , \55060 , \55067 );
and \U$54726 ( \55069 , \5318 , RI9870fd8_110);
and \U$54727 ( \55070 , RI9870b28_100, \5316 );
nor \U$54728 ( \55071 , \55069 , \55070 );
and \U$54729 ( \55072 , \55071 , \5322 );
not \U$54730 ( \55073 , \55071 );
and \U$54731 ( \55074 , \55073 , \5052 );
nor \U$54732 ( \55075 , \55072 , \55074 );
and \U$54733 ( \55076 , \55068 , \55075 );
and \U$54734 ( \55077 , \55060 , \55067 );
nor \U$54735 ( \55078 , \55076 , \55077 );
xor \U$54736 ( \55079 , \55053 , \55078 );
and \U$54737 ( \55080 , \4203 , RI986ffe8_76);
and \U$54738 ( \55081 , RI986fef8_74, \4201 );
nor \U$54739 ( \55082 , \55080 , \55081 );
and \U$54740 ( \55083 , \55082 , \4207 );
not \U$54741 ( \55084 , \55082 );
and \U$54742 ( \55085 , \55084 , \3922 );
nor \U$54743 ( \55086 , \55083 , \55085 );
not \U$54744 ( \55087 , \3412 );
and \U$54745 ( \55088 , \3683 , RI986fe08_72);
and \U$54746 ( \55089 , RI986fd18_70, \3681 );
nor \U$54747 ( \55090 , \55088 , \55089 );
not \U$54748 ( \55091 , \55090 );
or \U$54749 ( \55092 , \55087 , \55091 );
or \U$54750 ( \55093 , \55090 , \3412 );
nand \U$54751 ( \55094 , \55092 , \55093 );
xor \U$54752 ( \55095 , \55086 , \55094 );
not \U$54753 ( \55096 , \4521 );
and \U$54754 ( \55097 , \4710 , RI98700d8_78);
and \U$54755 ( \55098 , RI98701c8_80, \4708 );
nor \U$54756 ( \55099 , \55097 , \55098 );
not \U$54757 ( \55100 , \55099 );
or \U$54758 ( \55101 , \55096 , \55100 );
or \U$54759 ( \55102 , \55099 , \4519 );
nand \U$54760 ( \55103 , \55101 , \55102 );
and \U$54761 ( \55104 , \55095 , \55103 );
and \U$54762 ( \55105 , \55086 , \55094 );
or \U$54763 ( \55106 , \55104 , \55105 );
and \U$54764 ( \55107 , \55079 , \55106 );
and \U$54765 ( \55108 , \55053 , \55078 );
nor \U$54766 ( \55109 , \55107 , \55108 );
or \U$54767 ( \55110 , \55028 , \55109 );
not \U$54768 ( \55111 , \55109 );
not \U$54769 ( \55112 , \55028 );
or \U$54770 ( \55113 , \55111 , \55112 );
and \U$54771 ( \55114 , \12293 , RI986ef08_40);
and \U$54772 ( \55115 , RI986ee18_38, \12291 );
nor \U$54773 ( \55116 , \55114 , \55115 );
and \U$54774 ( \55117 , \55116 , \11686 );
not \U$54775 ( \55118 , \55116 );
and \U$54776 ( \55119 , \55118 , \11687 );
nor \U$54777 ( \55120 , \55117 , \55119 );
and \U$54778 ( \55121 , \13045 , RI986ec38_34);
and \U$54779 ( \55122 , RI986ed28_36, \13043 );
nor \U$54780 ( \55123 , \55121 , \55122 );
and \U$54781 ( \55124 , \55123 , \12619 );
not \U$54782 ( \55125 , \55123 );
and \U$54783 ( \55126 , \55125 , \13047 );
nor \U$54784 ( \55127 , \55124 , \55126 );
xor \U$54785 ( \55128 , \55120 , \55127 );
and \U$54786 ( \55129 , \11696 , RI986e968_28);
and \U$54787 ( \55130 , RI986e878_26, \11694 );
nor \U$54788 ( \55131 , \55129 , \55130 );
and \U$54789 ( \55132 , \55131 , \11702 );
not \U$54790 ( \55133 , \55131 );
and \U$54791 ( \55134 , \55133 , \10965 );
nor \U$54792 ( \55135 , \55132 , \55134 );
and \U$54793 ( \55136 , \55128 , \55135 );
and \U$54794 ( \55137 , \55120 , \55127 );
nor \U$54795 ( \55138 , \55136 , \55137 );
and \U$54796 ( \55139 , \15780 , RI986e5a8_20);
and \U$54797 ( \55140 , RI986e4b8_18, RI9873648_192);
nor \U$54798 ( \55141 , \55139 , \55140 );
not \U$54799 ( \55142 , \55141 );
not \U$54800 ( \55143 , RI9873558_190);
and \U$54801 ( \55144 , \55142 , \55143 );
and \U$54802 ( \55145 , \55141 , RI9873558_190);
nor \U$54803 ( \55146 , \55144 , \55145 );
and \U$54804 ( \55147 , \14937 , RI986f2c8_48);
and \U$54805 ( \55148 , RI986f1d8_46, \14935 );
nor \U$54806 ( \55149 , \55147 , \55148 );
and \U$54807 ( \55150 , \55149 , \14538 );
not \U$54808 ( \55151 , \55149 );
and \U$54809 ( \55152 , \55151 , \14539 );
nor \U$54810 ( \55153 , \55150 , \55152 );
xor \U$54811 ( \55154 , \55146 , \55153 );
and \U$54812 ( \55155 , \13882 , RI986f0e8_44);
and \U$54813 ( \55156 , RI986eff8_42, \13880 );
nor \U$54814 ( \55157 , \55155 , \55156 );
and \U$54815 ( \55158 , \55157 , \13359 );
not \U$54816 ( \55159 , \55157 );
and \U$54817 ( \55160 , \55159 , \13358 );
nor \U$54818 ( \55161 , \55158 , \55160 );
and \U$54819 ( \55162 , \55154 , \55161 );
and \U$54820 ( \55163 , \55146 , \55153 );
nor \U$54821 ( \55164 , \55162 , \55163 );
xor \U$54822 ( \55165 , \55138 , \55164 );
and \U$54823 ( \55166 , \9237 , RI9871758_126);
and \U$54824 ( \55167 , RI9871848_128, \9235 );
nor \U$54825 ( \55168 , \55166 , \55167 );
and \U$54826 ( \55169 , \55168 , \8836 );
not \U$54827 ( \55170 , \55168 );
and \U$54828 ( \55171 , \55170 , \9241 );
nor \U$54829 ( \55172 , \55169 , \55171 );
and \U$54830 ( \55173 , \10424 , RI986eb48_32);
and \U$54831 ( \55174 , RI986ea58_30, \10422 );
nor \U$54832 ( \55175 , \55173 , \55174 );
and \U$54833 ( \55176 , \55175 , \10428 );
not \U$54834 ( \55177 , \55175 );
and \U$54835 ( \55178 , \55177 , \9840 );
nor \U$54836 ( \55179 , \55176 , \55178 );
or \U$54837 ( \55180 , \55172 , \55179 );
not \U$54838 ( \55181 , \55179 );
not \U$54839 ( \55182 , \55172 );
or \U$54840 ( \55183 , \55181 , \55182 );
and \U$54841 ( \55184 , \9505 , RI9871578_122);
and \U$54842 ( \55185 , RI9871668_124, \9503 );
nor \U$54843 ( \55186 , \55184 , \55185 );
and \U$54844 ( \55187 , \55186 , \9510 );
not \U$54845 ( \55188 , \55186 );
and \U$54846 ( \55189 , \55188 , \9513 );
nor \U$54847 ( \55190 , \55187 , \55189 );
nand \U$54848 ( \55191 , \55183 , \55190 );
nand \U$54849 ( \55192 , \55180 , \55191 );
and \U$54850 ( \55193 , \55165 , \55192 );
and \U$54851 ( \55194 , \55138 , \55164 );
or \U$54852 ( \55195 , \55193 , \55194 );
nand \U$54853 ( \55196 , \55113 , \55195 );
nand \U$54854 ( \55197 , \55110 , \55196 );
xor \U$54855 ( \55198 , \54989 , \55197 );
not \U$54856 ( \55199 , \54655 );
not \U$54857 ( \55200 , \54671 );
or \U$54858 ( \55201 , \55199 , \55200 );
or \U$54859 ( \55202 , \54655 , \54671 );
nand \U$54860 ( \55203 , \55201 , \55202 );
not \U$54861 ( \55204 , \55203 );
not \U$54862 ( \55205 , \54665 );
and \U$54863 ( \55206 , \55204 , \55205 );
and \U$54864 ( \55207 , \55203 , \54665 );
nor \U$54865 ( \55208 , \55206 , \55207 );
xor \U$54866 ( \55209 , \54865 , \54892 );
xor \U$54867 ( \55210 , \55209 , \54895 );
or \U$54868 ( \55211 , \55208 , \55210 );
not \U$54869 ( \55212 , \55210 );
not \U$54870 ( \55213 , \55208 );
or \U$54871 ( \55214 , \55212 , \55213 );
xor \U$54872 ( \55215 , \54297 , \54304 );
xor \U$54873 ( \55216 , \55215 , \54312 );
xor \U$54874 ( \55217 , \54643 , \54648 );
xor \U$54875 ( \55218 , \55216 , \55217 );
nand \U$54876 ( \55219 , \55214 , \55218 );
nand \U$54877 ( \55220 , \55211 , \55219 );
xor \U$54878 ( \55221 , \55198 , \55220 );
not \U$54879 ( \55222 , \55221 );
or \U$54880 ( \55223 , \54957 , \55222 );
or \U$54881 ( \55224 , \55221 , \54956 );
xor \U$54882 ( \55225 , \54459 , \54488 );
xor \U$54883 ( \55226 , \55225 , \54514 );
xor \U$54884 ( \55227 , \54315 , \54341 );
xor \U$54885 ( \55228 , \55227 , \54367 );
xor \U$54886 ( \55229 , \55226 , \55228 );
xor \U$54887 ( \55230 , \54279 , \54281 );
xor \U$54888 ( \55231 , \55230 , \54284 );
xor \U$54889 ( \55232 , \54904 , \54911 );
xor \U$54890 ( \55233 , \55231 , \55232 );
xor \U$54891 ( \55234 , \55229 , \55233 );
nand \U$54892 ( \55235 , \55224 , \55234 );
nand \U$54893 ( \55236 , \55223 , \55235 );
xor \U$54894 ( \55237 , \54783 , \54808 );
xor \U$54895 ( \55238 , \55237 , \54835 );
xor \U$54896 ( \55239 , \54706 , \54727 );
xor \U$54897 ( \55240 , \55239 , \54753 );
and \U$54898 ( \55241 , \55238 , \55240 );
not \U$54899 ( \55242 , \55208 );
not \U$54900 ( \55243 , \55218 );
or \U$54901 ( \55244 , \55242 , \55243 );
or \U$54902 ( \55245 , \55208 , \55218 );
nand \U$54903 ( \55246 , \55244 , \55245 );
not \U$54904 ( \55247 , \55246 );
not \U$54905 ( \55248 , \55210 );
and \U$54906 ( \55249 , \55247 , \55248 );
and \U$54907 ( \55250 , \55246 , \55210 );
nor \U$54908 ( \55251 , \55249 , \55250 );
xor \U$54909 ( \55252 , \54706 , \54727 );
xor \U$54910 ( \55253 , \55252 , \54753 );
and \U$54911 ( \55254 , \55251 , \55253 );
and \U$54912 ( \55255 , \55238 , \55251 );
or \U$54913 ( \55256 , \55241 , \55254 , \55255 );
not \U$54914 ( \55257 , \55195 );
not \U$54915 ( \55258 , \55109 );
or \U$54916 ( \55259 , \55257 , \55258 );
or \U$54917 ( \55260 , \55109 , \55195 );
nand \U$54918 ( \55261 , \55259 , \55260 );
not \U$54919 ( \55262 , \55261 );
not \U$54920 ( \55263 , \55028 );
and \U$54921 ( \55264 , \55262 , \55263 );
and \U$54922 ( \55265 , \55261 , \55028 );
nor \U$54923 ( \55266 , \55264 , \55265 );
not \U$54924 ( \55267 , \55266 );
xor \U$54925 ( \55268 , \54973 , \54975 );
xor \U$54926 ( \55269 , \55268 , \54986 );
nand \U$54927 ( \55270 , \55267 , \55269 );
or \U$54928 ( \55271 , \55256 , \55270 );
not \U$54929 ( \55272 , \55270 );
not \U$54930 ( \55273 , \55256 );
or \U$54931 ( \55274 , \55272 , \55273 );
and \U$54932 ( \55275 , \2274 , RI98702b8_82);
and \U$54933 ( \55276 , RI9870768_92, \2272 );
nor \U$54934 ( \55277 , \55275 , \55276 );
and \U$54935 ( \55278 , \55277 , \2031 );
not \U$54936 ( \55279 , \55277 );
and \U$54937 ( \55280 , \55279 , \2030 );
nor \U$54938 ( \55281 , \55278 , \55280 );
not \U$54939 ( \55282 , \55281 );
nand \U$54940 ( \55283 , RI9870498_86, \1309 );
and \U$54941 ( \55284 , \55283 , \1315 );
not \U$54942 ( \55285 , \55283 );
and \U$54943 ( \55286 , \55285 , \1458 );
nor \U$54944 ( \55287 , \55284 , \55286 );
not \U$54945 ( \55288 , \55287 );
and \U$54946 ( \55289 , \55282 , \55288 );
and \U$54947 ( \55290 , \55281 , \55287 );
and \U$54948 ( \55291 , \2042 , RI9870588_88);
and \U$54949 ( \55292 , RI98703a8_84, \2040 );
nor \U$54950 ( \55293 , \55291 , \55292 );
not \U$54951 ( \55294 , \55293 );
not \U$54952 ( \55295 , \1462 );
and \U$54953 ( \55296 , \55294 , \55295 );
and \U$54954 ( \55297 , \55293 , \1462 );
nor \U$54955 ( \55298 , \55296 , \55297 );
nor \U$54956 ( \55299 , \55290 , \55298 );
nor \U$54957 ( \55300 , \55289 , \55299 );
and \U$54958 ( \55301 , \2042 , RI98703a8_84);
and \U$54959 ( \55302 , RI98702b8_82, \2040 );
nor \U$54960 ( \55303 , \55301 , \55302 );
not \U$54961 ( \55304 , \55303 );
not \U$54962 ( \55305 , \2034 );
and \U$54963 ( \55306 , \55304 , \55305 );
and \U$54964 ( \55307 , \55303 , \2034 );
nor \U$54965 ( \55308 , \55306 , \55307 );
xor \U$54966 ( \55309 , \55300 , \55308 );
and \U$54967 ( \55310 , \2464 , RI9870678_90);
and \U$54968 ( \55311 , RI9870948_96, \2462 );
nor \U$54969 ( \55312 , \55310 , \55311 );
and \U$54970 ( \55313 , \55312 , \2263 );
not \U$54971 ( \55314 , \55312 );
and \U$54972 ( \55315 , \55314 , \2468 );
nor \U$54973 ( \55316 , \55313 , \55315 );
not \U$54974 ( \55317 , \55316 );
and \U$54975 ( \55318 , \3683 , RI986fc28_68);
and \U$54976 ( \55319 , RI986fe08_72, \3681 );
nor \U$54977 ( \55320 , \55318 , \55319 );
not \U$54978 ( \55321 , \55320 );
not \U$54979 ( \55322 , \3918 );
and \U$54980 ( \55323 , \55321 , \55322 );
and \U$54981 ( \55324 , \55320 , \3918 );
nor \U$54982 ( \55325 , \55323 , \55324 );
not \U$54983 ( \55326 , \55325 );
and \U$54984 ( \55327 , \55317 , \55326 );
and \U$54985 ( \55328 , \55325 , \55316 );
and \U$54986 ( \55329 , \3254 , RI9870858_94);
and \U$54987 ( \55330 , RI986fb38_66, \3252 );
nor \U$54988 ( \55331 , \55329 , \55330 );
not \U$54989 ( \55332 , \55331 );
not \U$54990 ( \55333 , \3406 );
and \U$54991 ( \55334 , \55332 , \55333 );
and \U$54992 ( \55335 , \55331 , \3406 );
nor \U$54993 ( \55336 , \55334 , \55335 );
nor \U$54994 ( \55337 , \55328 , \55336 );
nor \U$54995 ( \55338 , \55327 , \55337 );
and \U$54996 ( \55339 , \55309 , \55338 );
and \U$54997 ( \55340 , \55300 , \55308 );
or \U$54998 ( \55341 , \55339 , \55340 );
not \U$54999 ( \55342 , \55341 );
and \U$55000 ( \55343 , \10424 , RI9871668_124);
and \U$55001 ( \55344 , RI986eb48_32, \10422 );
nor \U$55002 ( \55345 , \55343 , \55344 );
and \U$55003 ( \55346 , \55345 , \9840 );
not \U$55004 ( \55347 , \55345 );
and \U$55005 ( \55348 , \55347 , \10428 );
nor \U$55006 ( \55349 , \55346 , \55348 );
and \U$55007 ( \55350 , \11696 , RI986ea58_30);
and \U$55008 ( \55351 , RI986e968_28, \11694 );
nor \U$55009 ( \55352 , \55350 , \55351 );
and \U$55010 ( \55353 , \55352 , \10965 );
not \U$55011 ( \55354 , \55352 );
and \U$55012 ( \55355 , \55354 , \11702 );
nor \U$55013 ( \55356 , \55353 , \55355 );
xor \U$55014 ( \55357 , \55349 , \55356 );
and \U$55015 ( \55358 , \9505 , RI9871848_128);
and \U$55016 ( \55359 , RI9871578_122, \9503 );
nor \U$55017 ( \55360 , \55358 , \55359 );
and \U$55018 ( \55361 , \55360 , \9510 );
not \U$55019 ( \55362 , \55360 );
and \U$55020 ( \55363 , \55362 , \9513 );
nor \U$55021 ( \55364 , \55361 , \55363 );
and \U$55022 ( \55365 , \55357 , \55364 );
and \U$55023 ( \55366 , \55349 , \55356 );
nor \U$55024 ( \55367 , \55365 , \55366 );
and \U$55025 ( \55368 , \15780 , RI986f1d8_46);
and \U$55026 ( \55369 , RI986e5a8_20, RI9873648_192);
nor \U$55027 ( \55370 , \55368 , \55369 );
not \U$55028 ( \55371 , \55370 );
not \U$55029 ( \55372 , RI9873558_190);
and \U$55030 ( \55373 , \55371 , \55372 );
and \U$55031 ( \55374 , \55370 , RI9873558_190);
nor \U$55032 ( \55375 , \55373 , \55374 );
not \U$55033 ( \55376 , \55375 );
not \U$55034 ( \55377 , \1458 );
and \U$55035 ( \55378 , \55376 , \55377 );
and \U$55036 ( \55379 , \55375 , \1458 );
and \U$55037 ( \55380 , \14937 , RI986eff8_42);
and \U$55038 ( \55381 , RI986f2c8_48, \14935 );
nor \U$55039 ( \55382 , \55380 , \55381 );
and \U$55040 ( \55383 , \55382 , \14538 );
not \U$55041 ( \55384 , \55382 );
and \U$55042 ( \55385 , \55384 , \14539 );
nor \U$55043 ( \55386 , \55383 , \55385 );
nor \U$55044 ( \55387 , \55379 , \55386 );
nor \U$55045 ( \55388 , \55378 , \55387 );
xor \U$55046 ( \55389 , \55367 , \55388 );
and \U$55047 ( \55390 , \12293 , RI986e878_26);
and \U$55048 ( \55391 , RI986ef08_40, \12291 );
nor \U$55049 ( \55392 , \55390 , \55391 );
and \U$55050 ( \55393 , \55392 , \11686 );
not \U$55051 ( \55394 , \55392 );
and \U$55052 ( \55395 , \55394 , \11687 );
nor \U$55053 ( \55396 , \55393 , \55395 );
not \U$55054 ( \55397 , \55396 );
and \U$55055 ( \55398 , \13045 , RI986ee18_38);
and \U$55056 ( \55399 , RI986ec38_34, \13043 );
nor \U$55057 ( \55400 , \55398 , \55399 );
and \U$55058 ( \55401 , \55400 , \12619 );
not \U$55059 ( \55402 , \55400 );
and \U$55060 ( \55403 , \55402 , \13047 );
nor \U$55061 ( \55404 , \55401 , \55403 );
not \U$55062 ( \55405 , \55404 );
and \U$55063 ( \55406 , \55397 , \55405 );
and \U$55064 ( \55407 , \55404 , \55396 );
and \U$55065 ( \55408 , \13882 , RI986ed28_36);
and \U$55066 ( \55409 , RI986f0e8_44, \13880 );
nor \U$55067 ( \55410 , \55408 , \55409 );
and \U$55068 ( \55411 , \55410 , \13359 );
not \U$55069 ( \55412 , \55410 );
and \U$55070 ( \55413 , \55412 , \13358 );
nor \U$55071 ( \55414 , \55411 , \55413 );
nor \U$55072 ( \55415 , \55407 , \55414 );
nor \U$55073 ( \55416 , \55406 , \55415 );
and \U$55074 ( \55417 , \55389 , \55416 );
and \U$55075 ( \55418 , \55367 , \55388 );
or \U$55076 ( \55419 , \55417 , \55418 );
not \U$55077 ( \55420 , \55419 );
and \U$55078 ( \55421 , \55342 , \55420 );
and \U$55079 ( \55422 , \55341 , \55419 );
and \U$55080 ( \55423 , \7729 , RI9870d08_104);
and \U$55081 ( \55424 , RI98712a8_116, \7727 );
nor \U$55082 ( \55425 , \55423 , \55424 );
and \U$55083 ( \55426 , \55425 , \7480 );
not \U$55084 ( \55427 , \55425 );
and \U$55085 ( \55428 , \55427 , \7733 );
nor \U$55086 ( \55429 , \55426 , \55428 );
and \U$55087 ( \55430 , \8486 , RI98711b8_114);
and \U$55088 ( \55431 , RI9871398_118, \8484 );
nor \U$55089 ( \55432 , \55430 , \55431 );
and \U$55090 ( \55433 , \55432 , \8050 );
not \U$55091 ( \55434 , \55432 );
and \U$55092 ( \55435 , \55434 , \8051 );
nor \U$55093 ( \55436 , \55433 , \55435 );
xor \U$55094 ( \55437 , \55429 , \55436 );
and \U$55095 ( \55438 , \9237 , RI9871488_120);
and \U$55096 ( \55439 , RI9871758_126, \9235 );
nor \U$55097 ( \55440 , \55438 , \55439 );
and \U$55098 ( \55441 , \55440 , \9241 );
not \U$55099 ( \55442 , \55440 );
and \U$55100 ( \55443 , \55442 , \8836 );
nor \U$55101 ( \55444 , \55441 , \55443 );
and \U$55102 ( \55445 , \55437 , \55444 );
and \U$55103 ( \55446 , \55429 , \55436 );
or \U$55104 ( \55447 , \55445 , \55446 );
and \U$55105 ( \55448 , \7079 , RI9870c18_102);
and \U$55106 ( \55449 , RI98710c8_112, \7077 );
nor \U$55107 ( \55450 , \55448 , \55449 );
and \U$55108 ( \55451 , \55450 , \6710 );
not \U$55109 ( \55452 , \55450 );
and \U$55110 ( \55453 , \55452 , \6709 );
nor \U$55111 ( \55454 , \55451 , \55453 );
and \U$55112 ( \55455 , \5881 , RI9870b28_100);
and \U$55113 ( \55456 , RI9870df8_106, \5879 );
nor \U$55114 ( \55457 , \55455 , \55456 );
and \U$55115 ( \55458 , \55457 , \5594 );
not \U$55116 ( \55459 , \55457 );
and \U$55117 ( \55460 , \55459 , \5885 );
nor \U$55118 ( \55461 , \55458 , \55460 );
xor \U$55119 ( \55462 , \55454 , \55461 );
and \U$55120 ( \55463 , \6453 , RI9870a38_98);
and \U$55121 ( \55464 , RI9870ee8_108, \6451 );
nor \U$55122 ( \55465 , \55463 , \55464 );
and \U$55123 ( \55466 , \55465 , \6190 );
not \U$55124 ( \55467 , \55465 );
and \U$55125 ( \55468 , \55467 , \6180 );
nor \U$55126 ( \55469 , \55466 , \55468 );
and \U$55127 ( \55470 , \55462 , \55469 );
and \U$55128 ( \55471 , \55454 , \55461 );
or \U$55129 ( \55472 , \55470 , \55471 );
xor \U$55130 ( \55473 , \55447 , \55472 );
and \U$55131 ( \55474 , \5318 , RI98701c8_80);
and \U$55132 ( \55475 , RI9870fd8_110, \5316 );
nor \U$55133 ( \55476 , \55474 , \55475 );
and \U$55134 ( \55477 , \55476 , \5052 );
not \U$55135 ( \55478 , \55476 );
and \U$55136 ( \55479 , \55478 , \5322 );
nor \U$55137 ( \55480 , \55477 , \55479 );
and \U$55138 ( \55481 , \4203 , RI986fd18_70);
and \U$55139 ( \55482 , RI986ffe8_76, \4201 );
nor \U$55140 ( \55483 , \55481 , \55482 );
and \U$55141 ( \55484 , \55483 , \4207 );
not \U$55142 ( \55485 , \55483 );
and \U$55143 ( \55486 , \55485 , \3922 );
nor \U$55144 ( \55487 , \55484 , \55486 );
xor \U$55145 ( \55488 , \55480 , \55487 );
not \U$55146 ( \55489 , \4521 );
and \U$55147 ( \55490 , \4710 , RI986fef8_74);
and \U$55148 ( \55491 , RI98700d8_78, \4708 );
nor \U$55149 ( \55492 , \55490 , \55491 );
not \U$55150 ( \55493 , \55492 );
or \U$55151 ( \55494 , \55489 , \55493 );
or \U$55152 ( \55495 , \55492 , \4521 );
nand \U$55153 ( \55496 , \55494 , \55495 );
and \U$55154 ( \55497 , \55488 , \55496 );
and \U$55155 ( \55498 , \55480 , \55487 );
or \U$55156 ( \55499 , \55497 , \55498 );
and \U$55157 ( \55500 , \55473 , \55499 );
and \U$55158 ( \55501 , \55447 , \55472 );
nor \U$55159 ( \55502 , \55500 , \55501 );
nor \U$55160 ( \55503 , \55422 , \55502 );
nor \U$55161 ( \55504 , \55421 , \55503 );
not \U$55162 ( \55505 , \1336 );
not \U$55163 ( \55506 , \54714 );
not \U$55164 ( \55507 , \54725 );
or \U$55165 ( \55508 , \55506 , \55507 );
or \U$55166 ( \55509 , \54725 , \54714 );
nand \U$55167 ( \55510 , \55508 , \55509 );
not \U$55168 ( \55511 , \55510 );
or \U$55169 ( \55512 , \55505 , \55511 );
or \U$55170 ( \55513 , \55510 , \1336 );
nand \U$55171 ( \55514 , \55512 , \55513 );
and \U$55172 ( \55515 , \1311 , RI9870498_86);
and \U$55173 ( \55516 , RI9870588_88, \1309 );
nor \U$55174 ( \55517 , \55515 , \55516 );
and \U$55175 ( \55518 , \55517 , \1458 );
not \U$55176 ( \55519 , \55517 );
and \U$55177 ( \55520 , \55519 , \1318 );
nor \U$55178 ( \55521 , \55518 , \55520 );
xor \U$55179 ( \55522 , \55086 , \55094 );
xor \U$55180 ( \55523 , \55522 , \55103 );
and \U$55181 ( \55524 , \55521 , \55523 );
not \U$55182 ( \55525 , \54996 );
xor \U$55183 ( \55526 , \55015 , \55005 );
not \U$55184 ( \55527 , \55526 );
or \U$55185 ( \55528 , \55525 , \55527 );
or \U$55186 ( \55529 , \55526 , \54996 );
nand \U$55187 ( \55530 , \55528 , \55529 );
xor \U$55188 ( \55531 , \55086 , \55094 );
xor \U$55189 ( \55532 , \55531 , \55103 );
and \U$55190 ( \55533 , \55530 , \55532 );
and \U$55191 ( \55534 , \55521 , \55530 );
or \U$55192 ( \55535 , \55524 , \55533 , \55534 );
xor \U$55193 ( \55536 , \55514 , \55535 );
xor \U$55194 ( \55537 , \55060 , \55067 );
xor \U$55195 ( \55538 , \55537 , \55075 );
not \U$55196 ( \55539 , \55179 );
not \U$55197 ( \55540 , \55190 );
or \U$55198 ( \55541 , \55539 , \55540 );
or \U$55199 ( \55542 , \55179 , \55190 );
nand \U$55200 ( \55543 , \55541 , \55542 );
not \U$55201 ( \55544 , \55543 );
not \U$55202 ( \55545 , \55172 );
and \U$55203 ( \55546 , \55544 , \55545 );
and \U$55204 ( \55547 , \55543 , \55172 );
nor \U$55205 ( \55548 , \55546 , \55547 );
or \U$55206 ( \55549 , \55538 , \55548 );
not \U$55207 ( \55550 , \55548 );
not \U$55208 ( \55551 , \55538 );
or \U$55209 ( \55552 , \55550 , \55551 );
xor \U$55210 ( \55553 , \55035 , \55042 );
xor \U$55211 ( \55554 , \55553 , \55050 );
nand \U$55212 ( \55555 , \55552 , \55554 );
nand \U$55213 ( \55556 , \55549 , \55555 );
and \U$55214 ( \55557 , \55536 , \55556 );
and \U$55215 ( \55558 , \55514 , \55535 );
nor \U$55216 ( \55559 , \55557 , \55558 );
xor \U$55217 ( \55560 , \55504 , \55559 );
not \U$55218 ( \55561 , \54961 );
not \U$55219 ( \55562 , \54971 );
or \U$55220 ( \55563 , \55561 , \55562 );
or \U$55221 ( \55564 , \54961 , \54971 );
nand \U$55222 ( \55565 , \55563 , \55564 );
not \U$55223 ( \55566 , \55565 );
not \U$55224 ( \55567 , \54959 );
and \U$55225 ( \55568 , \55566 , \55567 );
and \U$55226 ( \55569 , \55565 , \54959 );
nor \U$55227 ( \55570 , \55568 , \55569 );
not \U$55228 ( \55571 , \55570 );
xor \U$55229 ( \55572 , \55017 , \55022 );
xor \U$55230 ( \55573 , \55572 , \55025 );
not \U$55231 ( \55574 , \55573 );
and \U$55232 ( \55575 , \55571 , \55574 );
and \U$55233 ( \55576 , \55570 , \55573 );
xor \U$55234 ( \55577 , \54978 , \54980 );
xor \U$55235 ( \55578 , \55577 , \54983 );
nor \U$55236 ( \55579 , \55576 , \55578 );
nor \U$55237 ( \55580 , \55575 , \55579 );
and \U$55238 ( \55581 , \55560 , \55580 );
and \U$55239 ( \55582 , \55504 , \55559 );
nor \U$55240 ( \55583 , \55581 , \55582 );
nand \U$55241 ( \55584 , \55274 , \55583 );
nand \U$55242 ( \55585 , \55271 , \55584 );
xor \U$55243 ( \55586 , \55236 , \55585 );
xor \U$55244 ( \55587 , \54681 , \54901 );
xor \U$55245 ( \55588 , \55587 , \54916 );
xor \U$55246 ( \55589 , \54370 , \54433 );
xor \U$55247 ( \55590 , \55589 , \54517 );
xor \U$55248 ( \55591 , \54260 , \54276 );
xor \U$55249 ( \55592 , \55591 , \54287 );
xor \U$55250 ( \55593 , \54618 , \54625 );
xor \U$55251 ( \55594 , \55592 , \55593 );
xor \U$55252 ( \55595 , \55590 , \55594 );
xor \U$55253 ( \55596 , \55588 , \55595 );
xor \U$55254 ( \55597 , \55586 , \55596 );
not \U$55255 ( \55598 , \55597 );
not \U$55256 ( \55599 , \1315 );
xnor \U$55257 ( \55600 , \55386 , \55375 );
not \U$55258 ( \55601 , \55600 );
or \U$55259 ( \55602 , \55599 , \55601 );
or \U$55260 ( \55603 , \55600 , \1318 );
nand \U$55261 ( \55604 , \55602 , \55603 );
xor \U$55262 ( \55605 , \55349 , \55356 );
xor \U$55263 ( \55606 , \55605 , \55364 );
xor \U$55264 ( \55607 , \55604 , \55606 );
not \U$55265 ( \55608 , \55396 );
xor \U$55266 ( \55609 , \55404 , \55414 );
not \U$55267 ( \55610 , \55609 );
or \U$55268 ( \55611 , \55608 , \55610 );
or \U$55269 ( \55612 , \55609 , \55396 );
nand \U$55270 ( \55613 , \55611 , \55612 );
and \U$55271 ( \55614 , \55607 , \55613 );
and \U$55272 ( \55615 , \55604 , \55606 );
nor \U$55273 ( \55616 , \55614 , \55615 );
xor \U$55274 ( \55617 , \55120 , \55127 );
xor \U$55275 ( \55618 , \55617 , \55135 );
or \U$55276 ( \55619 , \55616 , \55618 );
not \U$55277 ( \55620 , \55618 );
not \U$55278 ( \55621 , \55616 );
or \U$55279 ( \55622 , \55620 , \55621 );
xor \U$55280 ( \55623 , \55429 , \55436 );
xor \U$55281 ( \55624 , \55623 , \55444 );
xor \U$55282 ( \55625 , \55480 , \55487 );
xor \U$55283 ( \55626 , \55625 , \55496 );
xor \U$55284 ( \55627 , \55624 , \55626 );
xor \U$55285 ( \55628 , \55454 , \55461 );
xor \U$55286 ( \55629 , \55628 , \55469 );
and \U$55287 ( \55630 , \55627 , \55629 );
and \U$55288 ( \55631 , \55624 , \55626 );
or \U$55289 ( \55632 , \55630 , \55631 );
nand \U$55290 ( \55633 , \55622 , \55632 );
nand \U$55291 ( \55634 , \55619 , \55633 );
and \U$55292 ( \55635 , \7079 , RI9870ee8_108);
and \U$55293 ( \55636 , RI9870c18_102, \7077 );
nor \U$55294 ( \55637 , \55635 , \55636 );
and \U$55295 ( \55638 , \55637 , \6710 );
not \U$55296 ( \55639 , \55637 );
and \U$55297 ( \55640 , \55639 , \6709 );
nor \U$55298 ( \55641 , \55638 , \55640 );
and \U$55299 ( \55642 , \7729 , RI98710c8_112);
and \U$55300 ( \55643 , RI9870d08_104, \7727 );
nor \U$55301 ( \55644 , \55642 , \55643 );
and \U$55302 ( \55645 , \55644 , \7480 );
not \U$55303 ( \55646 , \55644 );
and \U$55304 ( \55647 , \55646 , \7733 );
nor \U$55305 ( \55648 , \55645 , \55647 );
xor \U$55306 ( \55649 , \55641 , \55648 );
and \U$55307 ( \55650 , \8486 , RI98712a8_116);
and \U$55308 ( \55651 , RI98711b8_114, \8484 );
nor \U$55309 ( \55652 , \55650 , \55651 );
and \U$55310 ( \55653 , \55652 , \8050 );
not \U$55311 ( \55654 , \55652 );
and \U$55312 ( \55655 , \55654 , \8051 );
nor \U$55313 ( \55656 , \55653 , \55655 );
and \U$55314 ( \55657 , \55649 , \55656 );
and \U$55315 ( \55658 , \55641 , \55648 );
or \U$55316 ( \55659 , \55657 , \55658 );
not \U$55317 ( \55660 , \3918 );
and \U$55318 ( \55661 , \3683 , RI986fb38_66);
and \U$55319 ( \55662 , RI986fc28_68, \3681 );
nor \U$55320 ( \55663 , \55661 , \55662 );
not \U$55321 ( \55664 , \55663 );
or \U$55322 ( \55665 , \55660 , \55664 );
or \U$55323 ( \55666 , \55663 , \3412 );
nand \U$55324 ( \55667 , \55665 , \55666 );
and \U$55325 ( \55668 , \4203 , RI986fe08_72);
and \U$55326 ( \55669 , RI986fd18_70, \4201 );
nor \U$55327 ( \55670 , \55668 , \55669 );
and \U$55328 ( \55671 , \55670 , \4207 );
not \U$55329 ( \55672 , \55670 );
and \U$55330 ( \55673 , \55672 , \3923 );
nor \U$55331 ( \55674 , \55671 , \55673 );
xor \U$55332 ( \55675 , \55667 , \55674 );
not \U$55333 ( \55676 , \4519 );
and \U$55334 ( \55677 , \4710 , RI986ffe8_76);
and \U$55335 ( \55678 , RI986fef8_74, \4708 );
nor \U$55336 ( \55679 , \55677 , \55678 );
not \U$55337 ( \55680 , \55679 );
or \U$55338 ( \55681 , \55676 , \55680 );
or \U$55339 ( \55682 , \55679 , \4519 );
nand \U$55340 ( \55683 , \55681 , \55682 );
and \U$55341 ( \55684 , \55675 , \55683 );
and \U$55342 ( \55685 , \55667 , \55674 );
or \U$55343 ( \55686 , \55684 , \55685 );
xor \U$55344 ( \55687 , \55659 , \55686 );
and \U$55345 ( \55688 , \5318 , RI98700d8_78);
and \U$55346 ( \55689 , RI98701c8_80, \5316 );
nor \U$55347 ( \55690 , \55688 , \55689 );
and \U$55348 ( \55691 , \55690 , \5052 );
not \U$55349 ( \55692 , \55690 );
and \U$55350 ( \55693 , \55692 , \5322 );
nor \U$55351 ( \55694 , \55691 , \55693 );
and \U$55352 ( \55695 , \5881 , RI9870fd8_110);
and \U$55353 ( \55696 , RI9870b28_100, \5879 );
nor \U$55354 ( \55697 , \55695 , \55696 );
and \U$55355 ( \55698 , \55697 , \5594 );
not \U$55356 ( \55699 , \55697 );
and \U$55357 ( \55700 , \55699 , \5885 );
nor \U$55358 ( \55701 , \55698 , \55700 );
xor \U$55359 ( \55702 , \55694 , \55701 );
and \U$55360 ( \55703 , \6453 , RI9870df8_106);
and \U$55361 ( \55704 , RI9870a38_98, \6451 );
nor \U$55362 ( \55705 , \55703 , \55704 );
and \U$55363 ( \55706 , \55705 , \6190 );
not \U$55364 ( \55707 , \55705 );
and \U$55365 ( \55708 , \55707 , \6180 );
nor \U$55366 ( \55709 , \55706 , \55708 );
and \U$55367 ( \55710 , \55702 , \55709 );
and \U$55368 ( \55711 , \55694 , \55701 );
or \U$55369 ( \55712 , \55710 , \55711 );
and \U$55370 ( \55713 , \55687 , \55712 );
and \U$55371 ( \55714 , \55659 , \55686 );
or \U$55372 ( \55715 , \55713 , \55714 );
and \U$55373 ( \55716 , \9237 , RI9871398_118);
and \U$55374 ( \55717 , RI9871488_120, \9235 );
nor \U$55375 ( \55718 , \55716 , \55717 );
and \U$55376 ( \55719 , \55718 , \9241 );
not \U$55377 ( \55720 , \55718 );
and \U$55378 ( \55721 , \55720 , \8836 );
nor \U$55379 ( \55722 , \55719 , \55721 );
and \U$55380 ( \55723 , \9505 , RI9871758_126);
and \U$55381 ( \55724 , RI9871848_128, \9503 );
nor \U$55382 ( \55725 , \55723 , \55724 );
and \U$55383 ( \55726 , \55725 , \9510 );
not \U$55384 ( \55727 , \55725 );
and \U$55385 ( \55728 , \55727 , \9513 );
nor \U$55386 ( \55729 , \55726 , \55728 );
xor \U$55387 ( \55730 , \55722 , \55729 );
and \U$55388 ( \55731 , \10424 , RI9871578_122);
and \U$55389 ( \55732 , RI9871668_124, \10422 );
nor \U$55390 ( \55733 , \55731 , \55732 );
and \U$55391 ( \55734 , \55733 , \9840 );
not \U$55392 ( \55735 , \55733 );
and \U$55393 ( \55736 , \55735 , \10428 );
nor \U$55394 ( \55737 , \55734 , \55736 );
and \U$55395 ( \55738 , \55730 , \55737 );
and \U$55396 ( \55739 , \55722 , \55729 );
or \U$55397 ( \55740 , \55738 , \55739 );
and \U$55398 ( \55741 , \13882 , RI986ec38_34);
and \U$55399 ( \55742 , RI986ed28_36, \13880 );
nor \U$55400 ( \55743 , \55741 , \55742 );
and \U$55401 ( \55744 , \55743 , \13358 );
not \U$55402 ( \55745 , \55743 );
and \U$55403 ( \55746 , \55745 , \13359 );
nor \U$55404 ( \55747 , \55744 , \55746 );
not \U$55405 ( \55748 , RI9873558_190);
and \U$55406 ( \55749 , \15780 , RI986f2c8_48);
and \U$55407 ( \55750 , RI986f1d8_46, RI9873648_192);
nor \U$55408 ( \55751 , \55749 , \55750 );
not \U$55409 ( \55752 , \55751 );
or \U$55410 ( \55753 , \55748 , \55752 );
or \U$55411 ( \55754 , \55751 , RI9873558_190);
nand \U$55412 ( \55755 , \55753 , \55754 );
xor \U$55413 ( \55756 , \55747 , \55755 );
and \U$55414 ( \55757 , \14937 , RI986f0e8_44);
and \U$55415 ( \55758 , RI986eff8_42, \14935 );
nor \U$55416 ( \55759 , \55757 , \55758 );
and \U$55417 ( \55760 , \55759 , \14539 );
not \U$55418 ( \55761 , \55759 );
and \U$55419 ( \55762 , \55761 , \14538 );
nor \U$55420 ( \55763 , \55760 , \55762 );
and \U$55421 ( \55764 , \55756 , \55763 );
and \U$55422 ( \55765 , \55747 , \55755 );
or \U$55423 ( \55766 , \55764 , \55765 );
xor \U$55424 ( \55767 , \55740 , \55766 );
and \U$55425 ( \55768 , \11696 , RI986eb48_32);
and \U$55426 ( \55769 , RI986ea58_30, \11694 );
nor \U$55427 ( \55770 , \55768 , \55769 );
and \U$55428 ( \55771 , \55770 , \10965 );
not \U$55429 ( \55772 , \55770 );
and \U$55430 ( \55773 , \55772 , \11702 );
nor \U$55431 ( \55774 , \55771 , \55773 );
and \U$55432 ( \55775 , \12293 , RI986e968_28);
and \U$55433 ( \55776 , RI986e878_26, \12291 );
nor \U$55434 ( \55777 , \55775 , \55776 );
and \U$55435 ( \55778 , \55777 , \11687 );
not \U$55436 ( \55779 , \55777 );
and \U$55437 ( \55780 , \55779 , \11686 );
nor \U$55438 ( \55781 , \55778 , \55780 );
xor \U$55439 ( \55782 , \55774 , \55781 );
and \U$55440 ( \55783 , \13045 , RI986ef08_40);
and \U$55441 ( \55784 , RI986ee18_38, \13043 );
nor \U$55442 ( \55785 , \55783 , \55784 );
and \U$55443 ( \55786 , \55785 , \13047 );
not \U$55444 ( \55787 , \55785 );
and \U$55445 ( \55788 , \55787 , \12619 );
nor \U$55446 ( \55789 , \55786 , \55788 );
and \U$55447 ( \55790 , \55782 , \55789 );
and \U$55448 ( \55791 , \55774 , \55781 );
or \U$55449 ( \55792 , \55790 , \55791 );
and \U$55450 ( \55793 , \55767 , \55792 );
and \U$55451 ( \55794 , \55740 , \55766 );
or \U$55452 ( \55795 , \55793 , \55794 );
xor \U$55453 ( \55796 , \55715 , \55795 );
not \U$55454 ( \55797 , \55287 );
xor \U$55455 ( \55798 , \55298 , \55281 );
not \U$55456 ( \55799 , \55798 );
or \U$55457 ( \55800 , \55797 , \55799 );
or \U$55458 ( \55801 , \55798 , \55287 );
nand \U$55459 ( \55802 , \55800 , \55801 );
and \U$55460 ( \55803 , \2274 , RI98703a8_84);
and \U$55461 ( \55804 , RI98702b8_82, \2272 );
nor \U$55462 ( \55805 , \55803 , \55804 );
and \U$55463 ( \55806 , \55805 , \2030 );
not \U$55464 ( \55807 , \55805 );
and \U$55465 ( \55808 , \55807 , \2031 );
nor \U$55466 ( \55809 , \55806 , \55808 );
and \U$55467 ( \55810 , \2464 , RI9870768_92);
and \U$55468 ( \55811 , RI9870678_90, \2462 );
nor \U$55469 ( \55812 , \55810 , \55811 );
and \U$55470 ( \55813 , \55812 , \2468 );
not \U$55471 ( \55814 , \55812 );
and \U$55472 ( \55815 , \55814 , \2263 );
nor \U$55473 ( \55816 , \55813 , \55815 );
xor \U$55474 ( \55817 , \55809 , \55816 );
not \U$55475 ( \55818 , \3406 );
and \U$55476 ( \55819 , \3254 , RI9870948_96);
and \U$55477 ( \55820 , RI9870858_94, \3252 );
nor \U$55478 ( \55821 , \55819 , \55820 );
not \U$55479 ( \55822 , \55821 );
or \U$55480 ( \55823 , \55818 , \55822 );
or \U$55481 ( \55824 , \55821 , \2935 );
nand \U$55482 ( \55825 , \55823 , \55824 );
and \U$55483 ( \55826 , \55817 , \55825 );
and \U$55484 ( \55827 , \55809 , \55816 );
or \U$55485 ( \55828 , \55826 , \55827 );
xor \U$55486 ( \55829 , \55802 , \55828 );
not \U$55487 ( \55830 , \55316 );
xor \U$55488 ( \55831 , \55336 , \55325 );
not \U$55489 ( \55832 , \55831 );
or \U$55490 ( \55833 , \55830 , \55832 );
or \U$55491 ( \55834 , \55831 , \55316 );
nand \U$55492 ( \55835 , \55833 , \55834 );
and \U$55493 ( \55836 , \55829 , \55835 );
and \U$55494 ( \55837 , \55802 , \55828 );
or \U$55495 ( \55838 , \55836 , \55837 );
and \U$55496 ( \55839 , \55796 , \55838 );
and \U$55497 ( \55840 , \55715 , \55795 );
or \U$55498 ( \55841 , \55839 , \55840 );
xor \U$55499 ( \55842 , \55634 , \55841 );
not \U$55500 ( \55843 , \55538 );
not \U$55501 ( \55844 , \55554 );
or \U$55502 ( \55845 , \55843 , \55844 );
or \U$55503 ( \55846 , \55538 , \55554 );
nand \U$55504 ( \55847 , \55845 , \55846 );
not \U$55505 ( \55848 , \55847 );
not \U$55506 ( \55849 , \55548 );
and \U$55507 ( \55850 , \55848 , \55849 );
and \U$55508 ( \55851 , \55847 , \55548 );
nor \U$55509 ( \55852 , \55850 , \55851 );
xor \U$55510 ( \55853 , \55146 , \55153 );
xor \U$55511 ( \55854 , \55853 , \55161 );
or \U$55512 ( \55855 , \55852 , \55854 );
not \U$55513 ( \55856 , \55854 );
not \U$55514 ( \55857 , \55852 );
or \U$55515 ( \55858 , \55856 , \55857 );
xor \U$55516 ( \55859 , \55086 , \55094 );
xor \U$55517 ( \55860 , \55859 , \55103 );
xor \U$55518 ( \55861 , \55521 , \55530 );
xor \U$55519 ( \55862 , \55860 , \55861 );
nand \U$55520 ( \55863 , \55858 , \55862 );
nand \U$55521 ( \55864 , \55855 , \55863 );
and \U$55522 ( \55865 , \55842 , \55864 );
and \U$55523 ( \55866 , \55634 , \55841 );
or \U$55524 ( \55867 , \55865 , \55866 );
xor \U$55525 ( \55868 , \55053 , \55078 );
xor \U$55526 ( \55869 , \55868 , \55106 );
xor \U$55527 ( \55870 , \55138 , \55164 );
xor \U$55528 ( \55871 , \55870 , \55192 );
xor \U$55529 ( \55872 , \55869 , \55871 );
xor \U$55530 ( \55873 , \55300 , \55308 );
xor \U$55531 ( \55874 , \55873 , \55338 );
xor \U$55532 ( \55875 , \55367 , \55388 );
xor \U$55533 ( \55876 , \55875 , \55416 );
or \U$55534 ( \55877 , \55874 , \55876 );
not \U$55535 ( \55878 , \55876 );
not \U$55536 ( \55879 , \55874 );
or \U$55537 ( \55880 , \55878 , \55879 );
xor \U$55538 ( \55881 , \55447 , \55472 );
xor \U$55539 ( \55882 , \55881 , \55499 );
nand \U$55540 ( \55883 , \55880 , \55882 );
nand \U$55541 ( \55884 , \55877 , \55883 );
and \U$55542 ( \55885 , \55872 , \55884 );
and \U$55543 ( \55886 , \55869 , \55871 );
or \U$55544 ( \55887 , \55885 , \55886 );
and \U$55545 ( \55888 , \55867 , \55887 );
xor \U$55546 ( \55889 , \55514 , \55535 );
xor \U$55547 ( \55890 , \55889 , \55556 );
not \U$55548 ( \55891 , \55341 );
xor \U$55549 ( \55892 , \55419 , \55502 );
not \U$55550 ( \55893 , \55892 );
or \U$55551 ( \55894 , \55891 , \55893 );
or \U$55552 ( \55895 , \55892 , \55341 );
nand \U$55553 ( \55896 , \55894 , \55895 );
xor \U$55554 ( \55897 , \55890 , \55896 );
not \U$55555 ( \55898 , \55570 );
xor \U$55556 ( \55899 , \55573 , \55578 );
not \U$55557 ( \55900 , \55899 );
or \U$55558 ( \55901 , \55898 , \55900 );
or \U$55559 ( \55902 , \55899 , \55570 );
nand \U$55560 ( \55903 , \55901 , \55902 );
and \U$55561 ( \55904 , \55897 , \55903 );
and \U$55562 ( \55905 , \55890 , \55896 );
or \U$55563 ( \55906 , \55904 , \55905 );
or \U$55564 ( \55907 , \55867 , \55887 );
and \U$55565 ( \55908 , \55906 , \55907 );
nor \U$55566 ( \55909 , \55888 , \55908 );
xor \U$55567 ( \55910 , \55504 , \55559 );
xor \U$55568 ( \55911 , \55910 , \55580 );
not \U$55569 ( \55912 , \55911 );
not \U$55570 ( \55913 , \55269 );
not \U$55571 ( \55914 , \55266 );
and \U$55572 ( \55915 , \55913 , \55914 );
and \U$55573 ( \55916 , \55269 , \55266 );
nor \U$55574 ( \55917 , \55915 , \55916 );
not \U$55575 ( \55918 , \55917 );
and \U$55576 ( \55919 , \55912 , \55918 );
and \U$55577 ( \55920 , \55911 , \55917 );
xor \U$55578 ( \55921 , \54706 , \54727 );
xor \U$55579 ( \55922 , \55921 , \54753 );
xor \U$55580 ( \55923 , \55238 , \55251 );
xor \U$55581 ( \55924 , \55922 , \55923 );
nor \U$55582 ( \55925 , \55920 , \55924 );
nor \U$55583 ( \55926 , \55919 , \55925 );
xor \U$55584 ( \55927 , \55909 , \55926 );
xnor \U$55585 ( \55928 , \55234 , \55221 );
not \U$55586 ( \55929 , \55928 );
not \U$55587 ( \55930 , \54956 );
and \U$55588 ( \55931 , \55929 , \55930 );
and \U$55589 ( \55932 , \55928 , \54956 );
nor \U$55590 ( \55933 , \55931 , \55932 );
and \U$55591 ( \55934 , \55927 , \55933 );
and \U$55592 ( \55935 , \55909 , \55926 );
nor \U$55593 ( \55936 , \55934 , \55935 );
not \U$55594 ( \55937 , \55936 );
xor \U$55595 ( \55938 , \54989 , \55197 );
and \U$55596 ( \55939 , \55938 , \55220 );
and \U$55597 ( \55940 , \54989 , \55197 );
or \U$55598 ( \55941 , \55939 , \55940 );
not \U$55599 ( \55942 , \55941 );
xor \U$55600 ( \55943 , \55226 , \55228 );
and \U$55601 ( \55944 , \55943 , \55233 );
and \U$55602 ( \55945 , \55226 , \55228 );
nor \U$55603 ( \55946 , \55944 , \55945 );
not \U$55604 ( \55947 , \55946 );
or \U$55605 ( \55948 , \55942 , \55947 );
or \U$55606 ( \55949 , \55946 , \55941 );
nand \U$55607 ( \55950 , \55948 , \55949 );
not \U$55608 ( \55951 , \55950 );
not \U$55609 ( \55952 , \54949 );
nand \U$55610 ( \55953 , \55952 , \54952 );
not \U$55611 ( \55954 , \55953 );
and \U$55612 ( \55955 , \55951 , \55954 );
and \U$55613 ( \55956 , \55950 , \55953 );
nor \U$55614 ( \55957 , \55955 , \55956 );
not \U$55615 ( \55958 , \55957 );
and \U$55616 ( \55959 , \55937 , \55958 );
and \U$55617 ( \55960 , \55936 , \55957 );
nor \U$55618 ( \55961 , \55959 , \55960 );
not \U$55619 ( \55962 , \55961 );
or \U$55620 ( \55963 , \55598 , \55962 );
or \U$55621 ( \55964 , \55961 , \55597 );
nand \U$55622 ( \55965 , \55963 , \55964 );
xor \U$55623 ( \55966 , \55909 , \55926 );
xor \U$55624 ( \55967 , \55966 , \55933 );
not \U$55625 ( \55968 , \55256 );
not \U$55626 ( \55969 , \55583 );
and \U$55627 ( \55970 , \55968 , \55969 );
and \U$55628 ( \55971 , \55256 , \55583 );
nor \U$55629 ( \55972 , \55970 , \55971 );
xnor \U$55630 ( \55973 , \55972 , \55270 );
or \U$55631 ( \55974 , \55967 , \55973 );
not \U$55632 ( \55975 , \55973 );
not \U$55633 ( \55976 , \55967 );
or \U$55634 ( \55977 , \55975 , \55976 );
not \U$55635 ( \55978 , \55632 );
not \U$55636 ( \55979 , \55616 );
or \U$55637 ( \55980 , \55978 , \55979 );
or \U$55638 ( \55981 , \55616 , \55632 );
nand \U$55639 ( \55982 , \55980 , \55981 );
not \U$55640 ( \55983 , \55982 );
not \U$55641 ( \55984 , \55618 );
and \U$55642 ( \55985 , \55983 , \55984 );
and \U$55643 ( \55986 , \55982 , \55618 );
nor \U$55644 ( \55987 , \55985 , \55986 );
not \U$55645 ( \55988 , \55876 );
not \U$55646 ( \55989 , \55882 );
or \U$55647 ( \55990 , \55988 , \55989 );
or \U$55648 ( \55991 , \55882 , \55876 );
nand \U$55649 ( \55992 , \55990 , \55991 );
not \U$55650 ( \55993 , \55992 );
not \U$55651 ( \55994 , \55874 );
and \U$55652 ( \55995 , \55993 , \55994 );
and \U$55653 ( \55996 , \55992 , \55874 );
nor \U$55654 ( \55997 , \55995 , \55996 );
xor \U$55655 ( \55998 , \55987 , \55997 );
not \U$55656 ( \55999 , \55854 );
not \U$55657 ( \56000 , \55862 );
or \U$55658 ( \56001 , \55999 , \56000 );
or \U$55659 ( \56002 , \55862 , \55854 );
nand \U$55660 ( \56003 , \56001 , \56002 );
not \U$55661 ( \56004 , \56003 );
not \U$55662 ( \56005 , \55852 );
and \U$55663 ( \56006 , \56004 , \56005 );
and \U$55664 ( \56007 , \56003 , \55852 );
nor \U$55665 ( \56008 , \56006 , \56007 );
and \U$55666 ( \56009 , \55998 , \56008 );
and \U$55667 ( \56010 , \55987 , \55997 );
nor \U$55668 ( \56011 , \56009 , \56010 );
xor \U$55669 ( \56012 , \55659 , \55686 );
xor \U$55670 ( \56013 , \56012 , \55712 );
xor \U$55671 ( \56014 , \55624 , \55626 );
xor \U$55672 ( \56015 , \56014 , \55629 );
and \U$55673 ( \56016 , \56013 , \56015 );
xor \U$55674 ( \56017 , \55802 , \55828 );
xor \U$55675 ( \56018 , \56017 , \55835 );
xor \U$55676 ( \56019 , \55624 , \55626 );
xor \U$55677 ( \56020 , \56019 , \55629 );
and \U$55678 ( \56021 , \56018 , \56020 );
and \U$55679 ( \56022 , \56013 , \56018 );
or \U$55680 ( \56023 , \56016 , \56021 , \56022 );
and \U$55681 ( \56024 , \9505 , RI9871488_120);
and \U$55682 ( \56025 , RI9871758_126, \9503 );
nor \U$55683 ( \56026 , \56024 , \56025 );
and \U$55684 ( \56027 , \56026 , \9510 );
not \U$55685 ( \56028 , \56026 );
and \U$55686 ( \56029 , \56028 , \9513 );
nor \U$55687 ( \56030 , \56027 , \56029 );
and \U$55688 ( \56031 , \10424 , RI9871848_128);
and \U$55689 ( \56032 , RI9871578_122, \10422 );
nor \U$55690 ( \56033 , \56031 , \56032 );
and \U$55691 ( \56034 , \56033 , \9840 );
not \U$55692 ( \56035 , \56033 );
and \U$55693 ( \56036 , \56035 , \10428 );
nor \U$55694 ( \56037 , \56034 , \56036 );
xor \U$55695 ( \56038 , \56030 , \56037 );
and \U$55696 ( \56039 , \11696 , RI9871668_124);
and \U$55697 ( \56040 , RI986eb48_32, \11694 );
nor \U$55698 ( \56041 , \56039 , \56040 );
and \U$55699 ( \56042 , \56041 , \10965 );
not \U$55700 ( \56043 , \56041 );
and \U$55701 ( \56044 , \56043 , \11702 );
nor \U$55702 ( \56045 , \56042 , \56044 );
and \U$55703 ( \56046 , \56038 , \56045 );
and \U$55704 ( \56047 , \56030 , \56037 );
or \U$55705 ( \56048 , \56046 , \56047 );
not \U$55706 ( \56049 , RI9873558_190);
and \U$55707 ( \56050 , \15780 , RI986eff8_42);
and \U$55708 ( \56051 , RI986f2c8_48, RI9873648_192);
nor \U$55709 ( \56052 , \56050 , \56051 );
not \U$55710 ( \56053 , \56052 );
or \U$55711 ( \56054 , \56049 , \56053 );
or \U$55712 ( \56055 , \56052 , RI9873558_190);
nand \U$55713 ( \56056 , \56054 , \56055 );
xor \U$55714 ( \56057 , \56056 , \1462 );
and \U$55715 ( \56058 , \14937 , RI986ed28_36);
and \U$55716 ( \56059 , RI986f0e8_44, \14935 );
nor \U$55717 ( \56060 , \56058 , \56059 );
and \U$55718 ( \56061 , \56060 , \14539 );
not \U$55719 ( \56062 , \56060 );
and \U$55720 ( \56063 , \56062 , \14538 );
nor \U$55721 ( \56064 , \56061 , \56063 );
and \U$55722 ( \56065 , \56057 , \56064 );
and \U$55723 ( \56066 , \56056 , \1462 );
or \U$55724 ( \56067 , \56065 , \56066 );
xor \U$55725 ( \56068 , \56048 , \56067 );
and \U$55726 ( \56069 , \12293 , RI986ea58_30);
and \U$55727 ( \56070 , RI986e968_28, \12291 );
nor \U$55728 ( \56071 , \56069 , \56070 );
and \U$55729 ( \56072 , \56071 , \11687 );
not \U$55730 ( \56073 , \56071 );
and \U$55731 ( \56074 , \56073 , \11686 );
nor \U$55732 ( \56075 , \56072 , \56074 );
and \U$55733 ( \56076 , \13045 , RI986e878_26);
and \U$55734 ( \56077 , RI986ef08_40, \13043 );
nor \U$55735 ( \56078 , \56076 , \56077 );
and \U$55736 ( \56079 , \56078 , \13047 );
not \U$55737 ( \56080 , \56078 );
and \U$55738 ( \56081 , \56080 , \12619 );
nor \U$55739 ( \56082 , \56079 , \56081 );
xor \U$55740 ( \56083 , \56075 , \56082 );
and \U$55741 ( \56084 , \13882 , RI986ee18_38);
and \U$55742 ( \56085 , RI986ec38_34, \13880 );
nor \U$55743 ( \56086 , \56084 , \56085 );
and \U$55744 ( \56087 , \56086 , \13358 );
not \U$55745 ( \56088 , \56086 );
and \U$55746 ( \56089 , \56088 , \13359 );
nor \U$55747 ( \56090 , \56087 , \56089 );
and \U$55748 ( \56091 , \56083 , \56090 );
and \U$55749 ( \56092 , \56075 , \56082 );
or \U$55750 ( \56093 , \56091 , \56092 );
and \U$55751 ( \56094 , \56068 , \56093 );
and \U$55752 ( \56095 , \56048 , \56067 );
or \U$55753 ( \56096 , \56094 , \56095 );
nand \U$55754 ( \56097 , RI9870498_86, \2040 );
not \U$55755 ( \56098 , \56097 );
not \U$55756 ( \56099 , \1462 );
or \U$55757 ( \56100 , \56098 , \56099 );
or \U$55758 ( \56101 , \1462 , \56097 );
nand \U$55759 ( \56102 , \56100 , \56101 );
and \U$55760 ( \56103 , \2274 , RI9870588_88);
and \U$55761 ( \56104 , RI98703a8_84, \2272 );
nor \U$55762 ( \56105 , \56103 , \56104 );
and \U$55763 ( \56106 , \56105 , \2030 );
not \U$55764 ( \56107 , \56105 );
and \U$55765 ( \56108 , \56107 , \2031 );
nor \U$55766 ( \56109 , \56106 , \56108 );
and \U$55767 ( \56110 , \56102 , \56109 );
not \U$55768 ( \56111 , \1462 );
and \U$55769 ( \56112 , \2042 , RI9870498_86);
and \U$55770 ( \56113 , RI9870588_88, \2040 );
nor \U$55771 ( \56114 , \56112 , \56113 );
not \U$55772 ( \56115 , \56114 );
or \U$55773 ( \56116 , \56111 , \56115 );
or \U$55774 ( \56117 , \56114 , \1462 );
nand \U$55775 ( \56118 , \56116 , \56117 );
xor \U$55776 ( \56119 , \56110 , \56118 );
not \U$55777 ( \56120 , \2935 );
and \U$55778 ( \56121 , \3254 , RI9870678_90);
and \U$55779 ( \56122 , RI9870948_96, \3252 );
nor \U$55780 ( \56123 , \56121 , \56122 );
not \U$55781 ( \56124 , \56123 );
or \U$55782 ( \56125 , \56120 , \56124 );
or \U$55783 ( \56126 , \56123 , \2935 );
nand \U$55784 ( \56127 , \56125 , \56126 );
and \U$55785 ( \56128 , \2464 , RI98702b8_82);
and \U$55786 ( \56129 , RI9870768_92, \2462 );
nor \U$55787 ( \56130 , \56128 , \56129 );
and \U$55788 ( \56131 , \56130 , \2468 );
not \U$55789 ( \56132 , \56130 );
and \U$55790 ( \56133 , \56132 , \2263 );
nor \U$55791 ( \56134 , \56131 , \56133 );
xor \U$55792 ( \56135 , \56127 , \56134 );
not \U$55793 ( \56136 , \3412 );
and \U$55794 ( \56137 , \3683 , RI9870858_94);
and \U$55795 ( \56138 , RI986fb38_66, \3681 );
nor \U$55796 ( \56139 , \56137 , \56138 );
not \U$55797 ( \56140 , \56139 );
or \U$55798 ( \56141 , \56136 , \56140 );
or \U$55799 ( \56142 , \56139 , \3412 );
nand \U$55800 ( \56143 , \56141 , \56142 );
and \U$55801 ( \56144 , \56135 , \56143 );
and \U$55802 ( \56145 , \56127 , \56134 );
or \U$55803 ( \56146 , \56144 , \56145 );
and \U$55804 ( \56147 , \56119 , \56146 );
and \U$55805 ( \56148 , \56110 , \56118 );
or \U$55806 ( \56149 , \56147 , \56148 );
xor \U$55807 ( \56150 , \56096 , \56149 );
and \U$55808 ( \56151 , \9237 , RI98711b8_114);
and \U$55809 ( \56152 , RI9871398_118, \9235 );
nor \U$55810 ( \56153 , \56151 , \56152 );
and \U$55811 ( \56154 , \56153 , \9241 );
not \U$55812 ( \56155 , \56153 );
and \U$55813 ( \56156 , \56155 , \8836 );
nor \U$55814 ( \56157 , \56154 , \56156 );
and \U$55815 ( \56158 , \7729 , RI9870c18_102);
and \U$55816 ( \56159 , RI98710c8_112, \7727 );
nor \U$55817 ( \56160 , \56158 , \56159 );
and \U$55818 ( \56161 , \56160 , \7480 );
not \U$55819 ( \56162 , \56160 );
and \U$55820 ( \56163 , \56162 , \7733 );
nor \U$55821 ( \56164 , \56161 , \56163 );
xor \U$55822 ( \56165 , \56157 , \56164 );
and \U$55823 ( \56166 , \8486 , RI9870d08_104);
and \U$55824 ( \56167 , RI98712a8_116, \8484 );
nor \U$55825 ( \56168 , \56166 , \56167 );
and \U$55826 ( \56169 , \56168 , \8050 );
not \U$55827 ( \56170 , \56168 );
and \U$55828 ( \56171 , \56170 , \8051 );
nor \U$55829 ( \56172 , \56169 , \56171 );
and \U$55830 ( \56173 , \56165 , \56172 );
and \U$55831 ( \56174 , \56157 , \56164 );
or \U$55832 ( \56175 , \56173 , \56174 );
and \U$55833 ( \56176 , \6453 , RI9870b28_100);
and \U$55834 ( \56177 , RI9870df8_106, \6451 );
nor \U$55835 ( \56178 , \56176 , \56177 );
and \U$55836 ( \56179 , \56178 , \6190 );
not \U$55837 ( \56180 , \56178 );
and \U$55838 ( \56181 , \56180 , \6705 );
nor \U$55839 ( \56182 , \56179 , \56181 );
and \U$55840 ( \56183 , \5881 , RI98701c8_80);
and \U$55841 ( \56184 , RI9870fd8_110, \5879 );
nor \U$55842 ( \56185 , \56183 , \56184 );
and \U$55843 ( \56186 , \56185 , \5594 );
not \U$55844 ( \56187 , \56185 );
and \U$55845 ( \56188 , \56187 , \5885 );
nor \U$55846 ( \56189 , \56186 , \56188 );
xor \U$55847 ( \56190 , \56182 , \56189 );
and \U$55848 ( \56191 , \7079 , RI9870a38_98);
and \U$55849 ( \56192 , RI9870ee8_108, \7077 );
nor \U$55850 ( \56193 , \56191 , \56192 );
and \U$55851 ( \56194 , \56193 , \6710 );
not \U$55852 ( \56195 , \56193 );
and \U$55853 ( \56196 , \56195 , \6709 );
nor \U$55854 ( \56197 , \56194 , \56196 );
and \U$55855 ( \56198 , \56190 , \56197 );
and \U$55856 ( \56199 , \56182 , \56189 );
or \U$55857 ( \56200 , \56198 , \56199 );
xor \U$55858 ( \56201 , \56175 , \56200 );
not \U$55859 ( \56202 , \4519 );
and \U$55860 ( \56203 , \4710 , RI986fd18_70);
and \U$55861 ( \56204 , RI986ffe8_76, \4708 );
nor \U$55862 ( \56205 , \56203 , \56204 );
not \U$55863 ( \56206 , \56205 );
or \U$55864 ( \56207 , \56202 , \56206 );
or \U$55865 ( \56208 , \56205 , \4521 );
nand \U$55866 ( \56209 , \56207 , \56208 );
and \U$55867 ( \56210 , \4203 , RI986fc28_68);
and \U$55868 ( \56211 , RI986fe08_72, \4201 );
nor \U$55869 ( \56212 , \56210 , \56211 );
and \U$55870 ( \56213 , \56212 , \4207 );
not \U$55871 ( \56214 , \56212 );
and \U$55872 ( \56215 , \56214 , \3923 );
nor \U$55873 ( \56216 , \56213 , \56215 );
xor \U$55874 ( \56217 , \56209 , \56216 );
and \U$55875 ( \56218 , \5318 , RI986fef8_74);
and \U$55876 ( \56219 , RI98700d8_78, \5316 );
nor \U$55877 ( \56220 , \56218 , \56219 );
and \U$55878 ( \56221 , \56220 , \5052 );
not \U$55879 ( \56222 , \56220 );
and \U$55880 ( \56223 , \56222 , \5322 );
nor \U$55881 ( \56224 , \56221 , \56223 );
and \U$55882 ( \56225 , \56217 , \56224 );
and \U$55883 ( \56226 , \56209 , \56216 );
or \U$55884 ( \56227 , \56225 , \56226 );
and \U$55885 ( \56228 , \56201 , \56227 );
and \U$55886 ( \56229 , \56175 , \56200 );
or \U$55887 ( \56230 , \56228 , \56229 );
and \U$55888 ( \56231 , \56150 , \56230 );
and \U$55889 ( \56232 , \56096 , \56149 );
or \U$55890 ( \56233 , \56231 , \56232 );
xor \U$55891 ( \56234 , \56023 , \56233 );
xor \U$55892 ( \56235 , \55774 , \55781 );
xor \U$55893 ( \56236 , \56235 , \55789 );
xor \U$55894 ( \56237 , \55641 , \55648 );
xor \U$55895 ( \56238 , \56237 , \55656 );
xor \U$55896 ( \56239 , \56236 , \56238 );
xor \U$55897 ( \56240 , \55722 , \55729 );
xor \U$55898 ( \56241 , \56240 , \55737 );
and \U$55899 ( \56242 , \56239 , \56241 );
and \U$55900 ( \56243 , \56236 , \56238 );
or \U$55901 ( \56244 , \56242 , \56243 );
xor \U$55902 ( \56245 , \55809 , \55816 );
xor \U$55903 ( \56246 , \56245 , \55825 );
xor \U$55904 ( \56247 , \55667 , \55674 );
xor \U$55905 ( \56248 , \56247 , \55683 );
and \U$55906 ( \56249 , \56246 , \56248 );
xor \U$55907 ( \56250 , \55694 , \55701 );
xor \U$55908 ( \56251 , \56250 , \55709 );
xor \U$55909 ( \56252 , \55667 , \55674 );
xor \U$55910 ( \56253 , \56252 , \55683 );
and \U$55911 ( \56254 , \56251 , \56253 );
and \U$55912 ( \56255 , \56246 , \56251 );
or \U$55913 ( \56256 , \56249 , \56254 , \56255 );
xor \U$55914 ( \56257 , \56244 , \56256 );
xor \U$55915 ( \56258 , \55604 , \55606 );
xor \U$55916 ( \56259 , \56258 , \55613 );
and \U$55917 ( \56260 , \56257 , \56259 );
and \U$55918 ( \56261 , \56244 , \56256 );
or \U$55919 ( \56262 , \56260 , \56261 );
and \U$55920 ( \56263 , \56234 , \56262 );
and \U$55921 ( \56264 , \56023 , \56233 );
or \U$55922 ( \56265 , \56263 , \56264 );
xor \U$55923 ( \56266 , \56011 , \56265 );
xor \U$55924 ( \56267 , \55890 , \55896 );
xor \U$55925 ( \56268 , \56267 , \55903 );
and \U$55926 ( \56269 , \56266 , \56268 );
and \U$55927 ( \56270 , \56011 , \56265 );
or \U$55928 ( \56271 , \56269 , \56270 );
not \U$55929 ( \56272 , \55906 );
xnor \U$55930 ( \56273 , \55887 , \55867 );
not \U$55931 ( \56274 , \56273 );
or \U$55932 ( \56275 , \56272 , \56274 );
or \U$55933 ( \56276 , \56273 , \55906 );
nand \U$55934 ( \56277 , \56275 , \56276 );
xor \U$55935 ( \56278 , \56271 , \56277 );
not \U$55936 ( \56279 , \55917 );
xor \U$55937 ( \56280 , \55924 , \55911 );
not \U$55938 ( \56281 , \56280 );
or \U$55939 ( \56282 , \56279 , \56281 );
or \U$55940 ( \56283 , \56280 , \55917 );
nand \U$55941 ( \56284 , \56282 , \56283 );
and \U$55942 ( \56285 , \56278 , \56284 );
and \U$55943 ( \56286 , \56271 , \56277 );
or \U$55944 ( \56287 , \56285 , \56286 );
nand \U$55945 ( \56288 , \55977 , \56287 );
nand \U$55946 ( \56289 , \55974 , \56288 );
and \U$55947 ( \56290 , \55965 , \56289 );
xor \U$55948 ( \56291 , \56289 , \55965 );
xor \U$55949 ( \56292 , \56271 , \56277 );
xor \U$55950 ( \56293 , \56292 , \56284 );
not \U$55951 ( \56294 , \56293 );
xor \U$55952 ( \56295 , \55634 , \55841 );
xor \U$55953 ( \56296 , \56295 , \55864 );
xor \U$55954 ( \56297 , \56011 , \56265 );
xor \U$55955 ( \56298 , \56297 , \56268 );
and \U$55956 ( \56299 , \56296 , \56298 );
not \U$55957 ( \56300 , \56299 );
xor \U$55958 ( \56301 , \55987 , \55997 );
xor \U$55959 ( \56302 , \56301 , \56008 );
not \U$55960 ( \56303 , \56302 );
xor \U$55961 ( \56304 , \56023 , \56233 );
xor \U$55962 ( \56305 , \56304 , \56262 );
nand \U$55963 ( \56306 , \56303 , \56305 );
not \U$55964 ( \56307 , \56306 );
xor \U$55965 ( \56308 , \55869 , \55871 );
xor \U$55966 ( \56309 , \56308 , \55884 );
and \U$55967 ( \56310 , \56307 , \56309 );
xor \U$55968 ( \56311 , \56030 , \56037 );
xor \U$55969 ( \56312 , \56311 , \56045 );
xor \U$55970 ( \56313 , \56056 , \1462 );
xor \U$55971 ( \56314 , \56313 , \56064 );
and \U$55972 ( \56315 , \56312 , \56314 );
xor \U$55973 ( \56316 , \56075 , \56082 );
xor \U$55974 ( \56317 , \56316 , \56090 );
xor \U$55975 ( \56318 , \56056 , \1462 );
xor \U$55976 ( \56319 , \56318 , \56064 );
and \U$55977 ( \56320 , \56317 , \56319 );
and \U$55978 ( \56321 , \56312 , \56317 );
or \U$55979 ( \56322 , \56315 , \56320 , \56321 );
xor \U$55980 ( \56323 , \55747 , \55755 );
xor \U$55981 ( \56324 , \56323 , \55763 );
xor \U$55982 ( \56325 , \56322 , \56324 );
xor \U$55983 ( \56326 , \56182 , \56189 );
xor \U$55984 ( \56327 , \56326 , \56197 );
xor \U$55985 ( \56328 , \56209 , \56216 );
xor \U$55986 ( \56329 , \56328 , \56224 );
xor \U$55987 ( \56330 , \56327 , \56329 );
xor \U$55988 ( \56331 , \56157 , \56164 );
xor \U$55989 ( \56332 , \56331 , \56172 );
and \U$55990 ( \56333 , \56330 , \56332 );
and \U$55991 ( \56334 , \56327 , \56329 );
or \U$55992 ( \56335 , \56333 , \56334 );
and \U$55993 ( \56336 , \56325 , \56335 );
and \U$55994 ( \56337 , \56322 , \56324 );
or \U$55995 ( \56338 , \56336 , \56337 );
and \U$55996 ( \56339 , \6453 , RI9870fd8_110);
and \U$55997 ( \56340 , RI9870b28_100, \6451 );
nor \U$55998 ( \56341 , \56339 , \56340 );
and \U$55999 ( \56342 , \56341 , \6190 );
not \U$56000 ( \56343 , \56341 );
and \U$56001 ( \56344 , \56343 , \6180 );
nor \U$56002 ( \56345 , \56342 , \56344 );
and \U$56003 ( \56346 , \5318 , RI986ffe8_76);
and \U$56004 ( \56347 , RI986fef8_74, \5316 );
nor \U$56005 ( \56348 , \56346 , \56347 );
and \U$56006 ( \56349 , \56348 , \5052 );
not \U$56007 ( \56350 , \56348 );
and \U$56008 ( \56351 , \56350 , \5322 );
nor \U$56009 ( \56352 , \56349 , \56351 );
xor \U$56010 ( \56353 , \56345 , \56352 );
and \U$56011 ( \56354 , \5881 , RI98700d8_78);
and \U$56012 ( \56355 , RI98701c8_80, \5879 );
nor \U$56013 ( \56356 , \56354 , \56355 );
and \U$56014 ( \56357 , \56356 , \5594 );
not \U$56015 ( \56358 , \56356 );
and \U$56016 ( \56359 , \56358 , \5885 );
nor \U$56017 ( \56360 , \56357 , \56359 );
and \U$56018 ( \56361 , \56353 , \56360 );
and \U$56019 ( \56362 , \56345 , \56352 );
or \U$56020 ( \56363 , \56361 , \56362 );
not \U$56021 ( \56364 , \3918 );
and \U$56022 ( \56365 , \3683 , RI9870948_96);
and \U$56023 ( \56366 , RI9870858_94, \3681 );
nor \U$56024 ( \56367 , \56365 , \56366 );
not \U$56025 ( \56368 , \56367 );
or \U$56026 ( \56369 , \56364 , \56368 );
or \U$56027 ( \56370 , \56367 , \3412 );
nand \U$56028 ( \56371 , \56369 , \56370 );
and \U$56029 ( \56372 , \4203 , RI986fb38_66);
and \U$56030 ( \56373 , RI986fc28_68, \4201 );
nor \U$56031 ( \56374 , \56372 , \56373 );
and \U$56032 ( \56375 , \56374 , \4207 );
not \U$56033 ( \56376 , \56374 );
and \U$56034 ( \56377 , \56376 , \3922 );
nor \U$56035 ( \56378 , \56375 , \56377 );
xor \U$56036 ( \56379 , \56371 , \56378 );
not \U$56037 ( \56380 , \4519 );
and \U$56038 ( \56381 , \4710 , RI986fe08_72);
and \U$56039 ( \56382 , RI986fd18_70, \4708 );
nor \U$56040 ( \56383 , \56381 , \56382 );
not \U$56041 ( \56384 , \56383 );
or \U$56042 ( \56385 , \56380 , \56384 );
or \U$56043 ( \56386 , \56383 , \4521 );
nand \U$56044 ( \56387 , \56385 , \56386 );
and \U$56045 ( \56388 , \56379 , \56387 );
and \U$56046 ( \56389 , \56371 , \56378 );
or \U$56047 ( \56390 , \56388 , \56389 );
xor \U$56048 ( \56391 , \56363 , \56390 );
and \U$56049 ( \56392 , \8486 , RI98710c8_112);
and \U$56050 ( \56393 , RI9870d08_104, \8484 );
nor \U$56051 ( \56394 , \56392 , \56393 );
and \U$56052 ( \56395 , \56394 , \8050 );
not \U$56053 ( \56396 , \56394 );
and \U$56054 ( \56397 , \56396 , \8051 );
nor \U$56055 ( \56398 , \56395 , \56397 );
and \U$56056 ( \56399 , \7079 , RI9870df8_106);
and \U$56057 ( \56400 , RI9870a38_98, \7077 );
nor \U$56058 ( \56401 , \56399 , \56400 );
and \U$56059 ( \56402 , \56401 , \6710 );
not \U$56060 ( \56403 , \56401 );
and \U$56061 ( \56404 , \56403 , \6709 );
nor \U$56062 ( \56405 , \56402 , \56404 );
xor \U$56063 ( \56406 , \56398 , \56405 );
and \U$56064 ( \56407 , \7729 , RI9870ee8_108);
and \U$56065 ( \56408 , RI9870c18_102, \7727 );
nor \U$56066 ( \56409 , \56407 , \56408 );
and \U$56067 ( \56410 , \56409 , \7480 );
not \U$56068 ( \56411 , \56409 );
and \U$56069 ( \56412 , \56411 , \7733 );
nor \U$56070 ( \56413 , \56410 , \56412 );
and \U$56071 ( \56414 , \56406 , \56413 );
and \U$56072 ( \56415 , \56398 , \56405 );
or \U$56073 ( \56416 , \56414 , \56415 );
and \U$56074 ( \56417 , \56391 , \56416 );
and \U$56075 ( \56418 , \56363 , \56390 );
or \U$56076 ( \56419 , \56417 , \56418 );
and \U$56077 ( \56420 , \9505 , RI9871398_118);
and \U$56078 ( \56421 , RI9871488_120, \9503 );
nor \U$56079 ( \56422 , \56420 , \56421 );
and \U$56080 ( \56423 , \56422 , \9510 );
not \U$56081 ( \56424 , \56422 );
and \U$56082 ( \56425 , \56424 , \9513 );
nor \U$56083 ( \56426 , \56423 , \56425 );
and \U$56084 ( \56427 , \9237 , RI98712a8_116);
and \U$56085 ( \56428 , RI98711b8_114, \9235 );
nor \U$56086 ( \56429 , \56427 , \56428 );
and \U$56087 ( \56430 , \56429 , \9241 );
not \U$56088 ( \56431 , \56429 );
and \U$56089 ( \56432 , \56431 , \8836 );
nor \U$56090 ( \56433 , \56430 , \56432 );
xor \U$56091 ( \56434 , \56426 , \56433 );
and \U$56092 ( \56435 , \10424 , RI9871758_126);
and \U$56093 ( \56436 , RI9871848_128, \10422 );
nor \U$56094 ( \56437 , \56435 , \56436 );
and \U$56095 ( \56438 , \56437 , \9840 );
not \U$56096 ( \56439 , \56437 );
and \U$56097 ( \56440 , \56439 , \10428 );
nor \U$56098 ( \56441 , \56438 , \56440 );
and \U$56099 ( \56442 , \56434 , \56441 );
and \U$56100 ( \56443 , \56426 , \56433 );
or \U$56101 ( \56444 , \56442 , \56443 );
and \U$56102 ( \56445 , \14937 , RI986ec38_34);
and \U$56103 ( \56446 , RI986ed28_36, \14935 );
nor \U$56104 ( \56447 , \56445 , \56446 );
and \U$56105 ( \56448 , \56447 , \14539 );
not \U$56106 ( \56449 , \56447 );
and \U$56107 ( \56450 , \56449 , \14538 );
nor \U$56108 ( \56451 , \56448 , \56450 );
not \U$56109 ( \56452 , RI9873558_190);
and \U$56110 ( \56453 , \15780 , RI986f0e8_44);
and \U$56111 ( \56454 , RI986eff8_42, RI9873648_192);
nor \U$56112 ( \56455 , \56453 , \56454 );
not \U$56113 ( \56456 , \56455 );
or \U$56114 ( \56457 , \56452 , \56456 );
or \U$56115 ( \56458 , \56455 , RI9873558_190);
nand \U$56116 ( \56459 , \56457 , \56458 );
xor \U$56117 ( \56460 , \56451 , \56459 );
and \U$56118 ( \56461 , \13882 , RI986ef08_40);
and \U$56119 ( \56462 , RI986ee18_38, \13880 );
nor \U$56120 ( \56463 , \56461 , \56462 );
and \U$56121 ( \56464 , \56463 , \13358 );
not \U$56122 ( \56465 , \56463 );
and \U$56123 ( \56466 , \56465 , \13359 );
nor \U$56124 ( \56467 , \56464 , \56466 );
and \U$56125 ( \56468 , \56460 , \56467 );
and \U$56126 ( \56469 , \56451 , \56459 );
or \U$56127 ( \56470 , \56468 , \56469 );
xor \U$56128 ( \56471 , \56444 , \56470 );
and \U$56129 ( \56472 , \11696 , RI9871578_122);
and \U$56130 ( \56473 , RI9871668_124, \11694 );
nor \U$56131 ( \56474 , \56472 , \56473 );
and \U$56132 ( \56475 , \56474 , \10965 );
not \U$56133 ( \56476 , \56474 );
and \U$56134 ( \56477 , \56476 , \11702 );
nor \U$56135 ( \56478 , \56475 , \56477 );
and \U$56136 ( \56479 , \12293 , RI986eb48_32);
and \U$56137 ( \56480 , RI986ea58_30, \12291 );
nor \U$56138 ( \56481 , \56479 , \56480 );
and \U$56139 ( \56482 , \56481 , \11687 );
not \U$56140 ( \56483 , \56481 );
and \U$56141 ( \56484 , \56483 , \11686 );
nor \U$56142 ( \56485 , \56482 , \56484 );
xor \U$56143 ( \56486 , \56478 , \56485 );
and \U$56144 ( \56487 , \13045 , RI986e968_28);
and \U$56145 ( \56488 , RI986e878_26, \13043 );
nor \U$56146 ( \56489 , \56487 , \56488 );
and \U$56147 ( \56490 , \56489 , \13047 );
not \U$56148 ( \56491 , \56489 );
and \U$56149 ( \56492 , \56491 , \12619 );
nor \U$56150 ( \56493 , \56490 , \56492 );
and \U$56151 ( \56494 , \56486 , \56493 );
and \U$56152 ( \56495 , \56478 , \56485 );
or \U$56153 ( \56496 , \56494 , \56495 );
and \U$56154 ( \56497 , \56471 , \56496 );
and \U$56155 ( \56498 , \56444 , \56470 );
or \U$56156 ( \56499 , \56497 , \56498 );
xor \U$56157 ( \56500 , \56419 , \56499 );
not \U$56158 ( \56501 , \2935 );
and \U$56159 ( \56502 , \3254 , RI9870768_92);
and \U$56160 ( \56503 , RI9870678_90, \3252 );
nor \U$56161 ( \56504 , \56502 , \56503 );
not \U$56162 ( \56505 , \56504 );
or \U$56163 ( \56506 , \56501 , \56505 );
or \U$56164 ( \56507 , \56504 , \3406 );
nand \U$56165 ( \56508 , \56506 , \56507 );
and \U$56166 ( \56509 , \2274 , RI9870498_86);
and \U$56167 ( \56510 , RI9870588_88, \2272 );
nor \U$56168 ( \56511 , \56509 , \56510 );
and \U$56169 ( \56512 , \56511 , \2030 );
not \U$56170 ( \56513 , \56511 );
and \U$56171 ( \56514 , \56513 , \2031 );
nor \U$56172 ( \56515 , \56512 , \56514 );
xor \U$56173 ( \56516 , \56508 , \56515 );
and \U$56174 ( \56517 , \2464 , RI98703a8_84);
and \U$56175 ( \56518 , RI98702b8_82, \2462 );
nor \U$56176 ( \56519 , \56517 , \56518 );
and \U$56177 ( \56520 , \56519 , \2468 );
not \U$56178 ( \56521 , \56519 );
and \U$56179 ( \56522 , \56521 , \2263 );
nor \U$56180 ( \56523 , \56520 , \56522 );
and \U$56181 ( \56524 , \56516 , \56523 );
and \U$56182 ( \56525 , \56508 , \56515 );
or \U$56183 ( \56526 , \56524 , \56525 );
xor \U$56184 ( \56527 , \56102 , \56109 );
xor \U$56185 ( \56528 , \56526 , \56527 );
xor \U$56186 ( \56529 , \56127 , \56134 );
xor \U$56187 ( \56530 , \56529 , \56143 );
and \U$56188 ( \56531 , \56528 , \56530 );
and \U$56189 ( \56532 , \56526 , \56527 );
or \U$56190 ( \56533 , \56531 , \56532 );
and \U$56191 ( \56534 , \56500 , \56533 );
and \U$56192 ( \56535 , \56419 , \56499 );
or \U$56193 ( \56536 , \56534 , \56535 );
xor \U$56194 ( \56537 , \56338 , \56536 );
xor \U$56195 ( \56538 , \56110 , \56118 );
xor \U$56196 ( \56539 , \56538 , \56146 );
xor \U$56197 ( \56540 , \56236 , \56238 );
xor \U$56198 ( \56541 , \56540 , \56241 );
and \U$56199 ( \56542 , \56539 , \56541 );
xor \U$56200 ( \56543 , \55667 , \55674 );
xor \U$56201 ( \56544 , \56543 , \55683 );
xor \U$56202 ( \56545 , \56246 , \56251 );
xor \U$56203 ( \56546 , \56544 , \56545 );
xor \U$56204 ( \56547 , \56236 , \56238 );
xor \U$56205 ( \56548 , \56547 , \56241 );
and \U$56206 ( \56549 , \56546 , \56548 );
and \U$56207 ( \56550 , \56539 , \56546 );
or \U$56208 ( \56551 , \56542 , \56549 , \56550 );
and \U$56209 ( \56552 , \56537 , \56551 );
and \U$56210 ( \56553 , \56338 , \56536 );
or \U$56211 ( \56554 , \56552 , \56553 );
xor \U$56212 ( \56555 , \55715 , \55795 );
xor \U$56213 ( \56556 , \56555 , \55838 );
xor \U$56214 ( \56557 , \56554 , \56556 );
xor \U$56215 ( \56558 , \55740 , \55766 );
xor \U$56216 ( \56559 , \56558 , \55792 );
xor \U$56217 ( \56560 , \56244 , \56256 );
xor \U$56218 ( \56561 , \56560 , \56259 );
and \U$56219 ( \56562 , \56559 , \56561 );
xor \U$56220 ( \56563 , \55624 , \55626 );
xor \U$56221 ( \56564 , \56563 , \55629 );
xor \U$56222 ( \56565 , \56013 , \56018 );
xor \U$56223 ( \56566 , \56564 , \56565 );
xor \U$56224 ( \56567 , \56244 , \56256 );
xor \U$56225 ( \56568 , \56567 , \56259 );
and \U$56226 ( \56569 , \56566 , \56568 );
and \U$56227 ( \56570 , \56559 , \56566 );
or \U$56228 ( \56571 , \56562 , \56569 , \56570 );
and \U$56229 ( \56572 , \56557 , \56571 );
and \U$56230 ( \56573 , \56554 , \56556 );
or \U$56231 ( \56574 , \56572 , \56573 );
not \U$56232 ( \56575 , \56309 );
nand \U$56233 ( \56576 , \56575 , \56306 );
and \U$56234 ( \56577 , \56574 , \56576 );
nor \U$56235 ( \56578 , \56310 , \56577 );
not \U$56236 ( \56579 , \56578 );
and \U$56237 ( \56580 , \56300 , \56579 );
and \U$56238 ( \56581 , \56299 , \56578 );
nor \U$56239 ( \56582 , \56580 , \56581 );
not \U$56240 ( \56583 , \56582 );
or \U$56241 ( \56584 , \56294 , \56583 );
or \U$56242 ( \56585 , \56293 , \56582 );
nand \U$56243 ( \56586 , \56584 , \56585 );
xor \U$56244 ( \56587 , \56296 , \56298 );
not \U$56245 ( \56588 , \56587 );
not \U$56246 ( \56589 , \56309 );
not \U$56247 ( \56590 , \56574 );
not \U$56248 ( \56591 , \56306 );
and \U$56249 ( \56592 , \56590 , \56591 );
and \U$56250 ( \56593 , \56574 , \56306 );
nor \U$56251 ( \56594 , \56592 , \56593 );
not \U$56252 ( \56595 , \56594 );
or \U$56253 ( \56596 , \56589 , \56595 );
or \U$56254 ( \56597 , \56594 , \56309 );
nand \U$56255 ( \56598 , \56596 , \56597 );
not \U$56256 ( \56599 , \56598 );
or \U$56257 ( \56600 , \56588 , \56599 );
or \U$56258 ( \56601 , \56598 , \56587 );
not \U$56259 ( \56602 , \56305 );
not \U$56260 ( \56603 , \56302 );
or \U$56261 ( \56604 , \56602 , \56603 );
or \U$56262 ( \56605 , \56302 , \56305 );
nand \U$56263 ( \56606 , \56604 , \56605 );
xor \U$56264 ( \56607 , \56175 , \56200 );
xor \U$56265 ( \56608 , \56607 , \56227 );
xor \U$56266 ( \56609 , \56048 , \56067 );
xor \U$56267 ( \56610 , \56609 , \56093 );
xor \U$56268 ( \56611 , \56608 , \56610 );
xor \U$56269 ( \56612 , \56236 , \56238 );
xor \U$56270 ( \56613 , \56612 , \56241 );
xor \U$56271 ( \56614 , \56539 , \56546 );
xor \U$56272 ( \56615 , \56613 , \56614 );
and \U$56273 ( \56616 , \56611 , \56615 );
and \U$56274 ( \56617 , \56608 , \56610 );
or \U$56275 ( \56618 , \56616 , \56617 );
xor \U$56276 ( \56619 , \56096 , \56149 );
xor \U$56277 ( \56620 , \56619 , \56230 );
xor \U$56278 ( \56621 , \56618 , \56620 );
xor \U$56279 ( \56622 , \56363 , \56390 );
xor \U$56280 ( \56623 , \56622 , \56416 );
xor \U$56281 ( \56624 , \56327 , \56329 );
xor \U$56282 ( \56625 , \56624 , \56332 );
and \U$56283 ( \56626 , \56623 , \56625 );
xor \U$56284 ( \56627 , \56526 , \56527 );
xor \U$56285 ( \56628 , \56627 , \56530 );
xor \U$56286 ( \56629 , \56327 , \56329 );
xor \U$56287 ( \56630 , \56629 , \56332 );
and \U$56288 ( \56631 , \56628 , \56630 );
and \U$56289 ( \56632 , \56623 , \56628 );
or \U$56290 ( \56633 , \56626 , \56631 , \56632 );
and \U$56291 ( \56634 , \9237 , RI9870d08_104);
and \U$56292 ( \56635 , RI98712a8_116, \9235 );
nor \U$56293 ( \56636 , \56634 , \56635 );
and \U$56294 ( \56637 , \56636 , \9241 );
not \U$56295 ( \56638 , \56636 );
and \U$56296 ( \56639 , \56638 , \8836 );
nor \U$56297 ( \56640 , \56637 , \56639 );
and \U$56298 ( \56641 , \7729 , RI9870a38_98);
and \U$56299 ( \56642 , RI9870ee8_108, \7727 );
nor \U$56300 ( \56643 , \56641 , \56642 );
and \U$56301 ( \56644 , \56643 , \7480 );
not \U$56302 ( \56645 , \56643 );
and \U$56303 ( \56646 , \56645 , \7733 );
nor \U$56304 ( \56647 , \56644 , \56646 );
xor \U$56305 ( \56648 , \56640 , \56647 );
and \U$56306 ( \56649 , \8486 , RI9870c18_102);
and \U$56307 ( \56650 , RI98710c8_112, \8484 );
nor \U$56308 ( \56651 , \56649 , \56650 );
and \U$56309 ( \56652 , \56651 , \8050 );
not \U$56310 ( \56653 , \56651 );
and \U$56311 ( \56654 , \56653 , \8051 );
nor \U$56312 ( \56655 , \56652 , \56654 );
and \U$56313 ( \56656 , \56648 , \56655 );
and \U$56314 ( \56657 , \56640 , \56647 );
or \U$56315 ( \56658 , \56656 , \56657 );
and \U$56316 ( \56659 , \5318 , RI986fd18_70);
and \U$56317 ( \56660 , RI986ffe8_76, \5316 );
nor \U$56318 ( \56661 , \56659 , \56660 );
and \U$56319 ( \56662 , \56661 , \5052 );
not \U$56320 ( \56663 , \56661 );
and \U$56321 ( \56664 , \56663 , \5322 );
nor \U$56322 ( \56665 , \56662 , \56664 );
and \U$56323 ( \56666 , \4203 , RI9870858_94);
and \U$56324 ( \56667 , RI986fb38_66, \4201 );
nor \U$56325 ( \56668 , \56666 , \56667 );
and \U$56326 ( \56669 , \56668 , \4207 );
not \U$56327 ( \56670 , \56668 );
and \U$56328 ( \56671 , \56670 , \3923 );
nor \U$56329 ( \56672 , \56669 , \56671 );
xor \U$56330 ( \56673 , \56665 , \56672 );
not \U$56331 ( \56674 , \4521 );
and \U$56332 ( \56675 , \4710 , RI986fc28_68);
and \U$56333 ( \56676 , RI986fe08_72, \4708 );
nor \U$56334 ( \56677 , \56675 , \56676 );
not \U$56335 ( \56678 , \56677 );
or \U$56336 ( \56679 , \56674 , \56678 );
or \U$56337 ( \56680 , \56677 , \4521 );
nand \U$56338 ( \56681 , \56679 , \56680 );
and \U$56339 ( \56682 , \56673 , \56681 );
and \U$56340 ( \56683 , \56665 , \56672 );
or \U$56341 ( \56684 , \56682 , \56683 );
xor \U$56342 ( \56685 , \56658 , \56684 );
and \U$56343 ( \56686 , \7079 , RI9870b28_100);
and \U$56344 ( \56687 , RI9870df8_106, \7077 );
nor \U$56345 ( \56688 , \56686 , \56687 );
and \U$56346 ( \56689 , \56688 , \6710 );
not \U$56347 ( \56690 , \56688 );
and \U$56348 ( \56691 , \56690 , \6709 );
nor \U$56349 ( \56692 , \56689 , \56691 );
and \U$56350 ( \56693 , \5881 , RI986fef8_74);
and \U$56351 ( \56694 , RI98700d8_78, \5879 );
nor \U$56352 ( \56695 , \56693 , \56694 );
and \U$56353 ( \56696 , \56695 , \5594 );
not \U$56354 ( \56697 , \56695 );
and \U$56355 ( \56698 , \56697 , \5885 );
nor \U$56356 ( \56699 , \56696 , \56698 );
xor \U$56357 ( \56700 , \56692 , \56699 );
and \U$56358 ( \56701 , \6453 , RI98701c8_80);
and \U$56359 ( \56702 , RI9870fd8_110, \6451 );
nor \U$56360 ( \56703 , \56701 , \56702 );
and \U$56361 ( \56704 , \56703 , \6190 );
not \U$56362 ( \56705 , \56703 );
and \U$56363 ( \56706 , \56705 , \6705 );
nor \U$56364 ( \56707 , \56704 , \56706 );
and \U$56365 ( \56708 , \56700 , \56707 );
and \U$56366 ( \56709 , \56692 , \56699 );
or \U$56367 ( \56710 , \56708 , \56709 );
and \U$56368 ( \56711 , \56685 , \56710 );
and \U$56369 ( \56712 , \56658 , \56684 );
or \U$56370 ( \56713 , \56711 , \56712 );
and \U$56371 ( \56714 , \9505 , RI98711b8_114);
and \U$56372 ( \56715 , RI9871398_118, \9503 );
nor \U$56373 ( \56716 , \56714 , \56715 );
and \U$56374 ( \56717 , \56716 , \9510 );
not \U$56375 ( \56718 , \56716 );
and \U$56376 ( \56719 , \56718 , \9513 );
nor \U$56377 ( \56720 , \56717 , \56719 );
and \U$56378 ( \56721 , \10424 , RI9871488_120);
and \U$56379 ( \56722 , RI9871758_126, \10422 );
nor \U$56380 ( \56723 , \56721 , \56722 );
and \U$56381 ( \56724 , \56723 , \9840 );
not \U$56382 ( \56725 , \56723 );
and \U$56383 ( \56726 , \56725 , \10428 );
nor \U$56384 ( \56727 , \56724 , \56726 );
xor \U$56385 ( \56728 , \56720 , \56727 );
and \U$56386 ( \56729 , \11696 , RI9871848_128);
and \U$56387 ( \56730 , RI9871578_122, \11694 );
nor \U$56388 ( \56731 , \56729 , \56730 );
and \U$56389 ( \56732 , \56731 , \10965 );
not \U$56390 ( \56733 , \56731 );
and \U$56391 ( \56734 , \56733 , \11702 );
nor \U$56392 ( \56735 , \56732 , \56734 );
and \U$56393 ( \56736 , \56728 , \56735 );
and \U$56394 ( \56737 , \56720 , \56727 );
or \U$56395 ( \56738 , \56736 , \56737 );
not \U$56396 ( \56739 , RI9873558_190);
and \U$56397 ( \56740 , \15780 , RI986ed28_36);
and \U$56398 ( \56741 , RI986f0e8_44, RI9873648_192);
nor \U$56399 ( \56742 , \56740 , \56741 );
not \U$56400 ( \56743 , \56742 );
or \U$56401 ( \56744 , \56739 , \56743 );
or \U$56402 ( \56745 , \56742 , RI9873558_190);
nand \U$56403 ( \56746 , \56744 , \56745 );
xor \U$56404 ( \56747 , \56746 , \2031 );
and \U$56405 ( \56748 , \14937 , RI986ee18_38);
and \U$56406 ( \56749 , RI986ec38_34, \14935 );
nor \U$56407 ( \56750 , \56748 , \56749 );
and \U$56408 ( \56751 , \56750 , \14539 );
not \U$56409 ( \56752 , \56750 );
and \U$56410 ( \56753 , \56752 , \14538 );
nor \U$56411 ( \56754 , \56751 , \56753 );
and \U$56412 ( \56755 , \56747 , \56754 );
and \U$56413 ( \56756 , \56746 , \2031 );
or \U$56414 ( \56757 , \56755 , \56756 );
xor \U$56415 ( \56758 , \56738 , \56757 );
and \U$56416 ( \56759 , \13882 , RI986e878_26);
and \U$56417 ( \56760 , RI986ef08_40, \13880 );
nor \U$56418 ( \56761 , \56759 , \56760 );
and \U$56419 ( \56762 , \56761 , \13358 );
not \U$56420 ( \56763 , \56761 );
and \U$56421 ( \56764 , \56763 , \13359 );
nor \U$56422 ( \56765 , \56762 , \56764 );
and \U$56423 ( \56766 , \12293 , RI9871668_124);
and \U$56424 ( \56767 , RI986eb48_32, \12291 );
nor \U$56425 ( \56768 , \56766 , \56767 );
and \U$56426 ( \56769 , \56768 , \11687 );
not \U$56427 ( \56770 , \56768 );
and \U$56428 ( \56771 , \56770 , \11686 );
nor \U$56429 ( \56772 , \56769 , \56771 );
xor \U$56430 ( \56773 , \56765 , \56772 );
and \U$56431 ( \56774 , \13045 , RI986ea58_30);
and \U$56432 ( \56775 , RI986e968_28, \13043 );
nor \U$56433 ( \56776 , \56774 , \56775 );
and \U$56434 ( \56777 , \56776 , \13047 );
not \U$56435 ( \56778 , \56776 );
and \U$56436 ( \56779 , \56778 , \12619 );
nor \U$56437 ( \56780 , \56777 , \56779 );
and \U$56438 ( \56781 , \56773 , \56780 );
and \U$56439 ( \56782 , \56765 , \56772 );
or \U$56440 ( \56783 , \56781 , \56782 );
and \U$56441 ( \56784 , \56758 , \56783 );
and \U$56442 ( \56785 , \56738 , \56757 );
or \U$56443 ( \56786 , \56784 , \56785 );
xor \U$56444 ( \56787 , \56713 , \56786 );
and \U$56445 ( \56788 , \2464 , RI9870588_88);
and \U$56446 ( \56789 , RI98703a8_84, \2462 );
nor \U$56447 ( \56790 , \56788 , \56789 );
and \U$56448 ( \56791 , \56790 , \2468 );
not \U$56449 ( \56792 , \56790 );
and \U$56450 ( \56793 , \56792 , \2263 );
nor \U$56451 ( \56794 , \56791 , \56793 );
not \U$56452 ( \56795 , \3406 );
and \U$56453 ( \56796 , \3254 , RI98702b8_82);
and \U$56454 ( \56797 , RI9870768_92, \3252 );
nor \U$56455 ( \56798 , \56796 , \56797 );
not \U$56456 ( \56799 , \56798 );
or \U$56457 ( \56800 , \56795 , \56799 );
or \U$56458 ( \56801 , \56798 , \3406 );
nand \U$56459 ( \56802 , \56800 , \56801 );
xor \U$56460 ( \56803 , \56794 , \56802 );
not \U$56461 ( \56804 , \3918 );
and \U$56462 ( \56805 , \3683 , RI9870678_90);
and \U$56463 ( \56806 , RI9870948_96, \3681 );
nor \U$56464 ( \56807 , \56805 , \56806 );
not \U$56465 ( \56808 , \56807 );
or \U$56466 ( \56809 , \56804 , \56808 );
or \U$56467 ( \56810 , \56807 , \3412 );
nand \U$56468 ( \56811 , \56809 , \56810 );
and \U$56469 ( \56812 , \56803 , \56811 );
and \U$56470 ( \56813 , \56794 , \56802 );
or \U$56471 ( \56814 , \56812 , \56813 );
xor \U$56472 ( \56815 , \56508 , \56515 );
xor \U$56473 ( \56816 , \56815 , \56523 );
and \U$56474 ( \56817 , \56814 , \56816 );
xor \U$56475 ( \56818 , \56371 , \56378 );
xor \U$56476 ( \56819 , \56818 , \56387 );
xor \U$56477 ( \56820 , \56508 , \56515 );
xor \U$56478 ( \56821 , \56820 , \56523 );
and \U$56479 ( \56822 , \56819 , \56821 );
and \U$56480 ( \56823 , \56814 , \56819 );
or \U$56481 ( \56824 , \56817 , \56822 , \56823 );
and \U$56482 ( \56825 , \56787 , \56824 );
and \U$56483 ( \56826 , \56713 , \56786 );
or \U$56484 ( \56827 , \56825 , \56826 );
xor \U$56485 ( \56828 , \56633 , \56827 );
xor \U$56486 ( \56829 , \56345 , \56352 );
xor \U$56487 ( \56830 , \56829 , \56360 );
xor \U$56488 ( \56831 , \56426 , \56433 );
xor \U$56489 ( \56832 , \56831 , \56441 );
and \U$56490 ( \56833 , \56830 , \56832 );
xor \U$56491 ( \56834 , \56398 , \56405 );
xor \U$56492 ( \56835 , \56834 , \56413 );
xor \U$56493 ( \56836 , \56426 , \56433 );
xor \U$56494 ( \56837 , \56836 , \56441 );
and \U$56495 ( \56838 , \56835 , \56837 );
and \U$56496 ( \56839 , \56830 , \56835 );
or \U$56497 ( \56840 , \56833 , \56838 , \56839 );
xor \U$56498 ( \56841 , \56478 , \56485 );
xor \U$56499 ( \56842 , \56841 , \56493 );
xor \U$56500 ( \56843 , \56451 , \56459 );
xor \U$56501 ( \56844 , \56843 , \56467 );
and \U$56502 ( \56845 , \56842 , \56844 );
xor \U$56503 ( \56846 , \56840 , \56845 );
xor \U$56504 ( \56847 , \56056 , \1462 );
xor \U$56505 ( \56848 , \56847 , \56064 );
xor \U$56506 ( \56849 , \56312 , \56317 );
xor \U$56507 ( \56850 , \56848 , \56849 );
and \U$56508 ( \56851 , \56846 , \56850 );
and \U$56509 ( \56852 , \56840 , \56845 );
or \U$56510 ( \56853 , \56851 , \56852 );
and \U$56511 ( \56854 , \56828 , \56853 );
and \U$56512 ( \56855 , \56633 , \56827 );
or \U$56513 ( \56856 , \56854 , \56855 );
and \U$56514 ( \56857 , \56621 , \56856 );
and \U$56515 ( \56858 , \56618 , \56620 );
or \U$56516 ( \56859 , \56857 , \56858 );
xor \U$56517 ( \56860 , \56606 , \56859 );
xor \U$56518 ( \56861 , \56554 , \56556 );
xor \U$56519 ( \56862 , \56861 , \56571 );
and \U$56520 ( \56863 , \56860 , \56862 );
and \U$56521 ( \56864 , \56606 , \56859 );
or \U$56522 ( \56865 , \56863 , \56864 );
nand \U$56523 ( \56866 , \56601 , \56865 );
nand \U$56524 ( \56867 , \56600 , \56866 );
and \U$56525 ( \56868 , \56586 , \56867 );
xor \U$56526 ( \56869 , \56867 , \56586 );
xor \U$56527 ( \56870 , \56419 , \56499 );
xor \U$56528 ( \56871 , \56870 , \56533 );
xor \U$56529 ( \56872 , \56608 , \56610 );
xor \U$56530 ( \56873 , \56872 , \56615 );
and \U$56531 ( \56874 , \56871 , \56873 );
xor \U$56532 ( \56875 , \56633 , \56827 );
xor \U$56533 ( \56876 , \56875 , \56853 );
xor \U$56534 ( \56877 , \56608 , \56610 );
xor \U$56535 ( \56878 , \56877 , \56615 );
and \U$56536 ( \56879 , \56876 , \56878 );
and \U$56537 ( \56880 , \56871 , \56876 );
or \U$56538 ( \56881 , \56874 , \56879 , \56880 );
xor \U$56539 ( \56882 , \56244 , \56256 );
xor \U$56540 ( \56883 , \56882 , \56259 );
xor \U$56541 ( \56884 , \56559 , \56566 );
xor \U$56542 ( \56885 , \56883 , \56884 );
xor \U$56543 ( \56886 , \56881 , \56885 );
xor \U$56544 ( \56887 , \56658 , \56684 );
xor \U$56545 ( \56888 , \56887 , \56710 );
xor \U$56546 ( \56889 , \56738 , \56757 );
xor \U$56547 ( \56890 , \56889 , \56783 );
xor \U$56548 ( \56891 , \56888 , \56890 );
xor \U$56549 ( \56892 , \56508 , \56515 );
xor \U$56550 ( \56893 , \56892 , \56523 );
xor \U$56551 ( \56894 , \56814 , \56819 );
xor \U$56552 ( \56895 , \56893 , \56894 );
and \U$56553 ( \56896 , \56891 , \56895 );
and \U$56554 ( \56897 , \56888 , \56890 );
or \U$56555 ( \56898 , \56896 , \56897 );
and \U$56556 ( \56899 , \7079 , RI9870fd8_110);
and \U$56557 ( \56900 , RI9870b28_100, \7077 );
nor \U$56558 ( \56901 , \56899 , \56900 );
and \U$56559 ( \56902 , \56901 , \6710 );
not \U$56560 ( \56903 , \56901 );
and \U$56561 ( \56904 , \56903 , \6709 );
nor \U$56562 ( \56905 , \56902 , \56904 );
and \U$56563 ( \56906 , \7729 , RI9870df8_106);
and \U$56564 ( \56907 , RI9870a38_98, \7727 );
nor \U$56565 ( \56908 , \56906 , \56907 );
and \U$56566 ( \56909 , \56908 , \7480 );
not \U$56567 ( \56910 , \56908 );
and \U$56568 ( \56911 , \56910 , \7733 );
nor \U$56569 ( \56912 , \56909 , \56911 );
xor \U$56570 ( \56913 , \56905 , \56912 );
and \U$56571 ( \56914 , \8486 , RI9870ee8_108);
and \U$56572 ( \56915 , RI9870c18_102, \8484 );
nor \U$56573 ( \56916 , \56914 , \56915 );
and \U$56574 ( \56917 , \56916 , \8050 );
not \U$56575 ( \56918 , \56916 );
and \U$56576 ( \56919 , \56918 , \8051 );
nor \U$56577 ( \56920 , \56917 , \56919 );
and \U$56578 ( \56921 , \56913 , \56920 );
and \U$56579 ( \56922 , \56905 , \56912 );
or \U$56580 ( \56923 , \56921 , \56922 );
and \U$56581 ( \56924 , \5318 , RI986fe08_72);
and \U$56582 ( \56925 , RI986fd18_70, \5316 );
nor \U$56583 ( \56926 , \56924 , \56925 );
and \U$56584 ( \56927 , \56926 , \5052 );
not \U$56585 ( \56928 , \56926 );
and \U$56586 ( \56929 , \56928 , \5322 );
nor \U$56587 ( \56930 , \56927 , \56929 );
and \U$56588 ( \56931 , \5881 , RI986ffe8_76);
and \U$56589 ( \56932 , RI986fef8_74, \5879 );
nor \U$56590 ( \56933 , \56931 , \56932 );
and \U$56591 ( \56934 , \56933 , \5594 );
not \U$56592 ( \56935 , \56933 );
and \U$56593 ( \56936 , \56935 , \5885 );
nor \U$56594 ( \56937 , \56934 , \56936 );
xor \U$56595 ( \56938 , \56930 , \56937 );
and \U$56596 ( \56939 , \6453 , RI98700d8_78);
and \U$56597 ( \56940 , RI98701c8_80, \6451 );
nor \U$56598 ( \56941 , \56939 , \56940 );
and \U$56599 ( \56942 , \56941 , \6190 );
not \U$56600 ( \56943 , \56941 );
and \U$56601 ( \56944 , \56943 , \6705 );
nor \U$56602 ( \56945 , \56942 , \56944 );
and \U$56603 ( \56946 , \56938 , \56945 );
and \U$56604 ( \56947 , \56930 , \56937 );
or \U$56605 ( \56948 , \56946 , \56947 );
xor \U$56606 ( \56949 , \56923 , \56948 );
not \U$56607 ( \56950 , \3412 );
and \U$56608 ( \56951 , \3683 , RI9870768_92);
and \U$56609 ( \56952 , RI9870678_90, \3681 );
nor \U$56610 ( \56953 , \56951 , \56952 );
not \U$56611 ( \56954 , \56953 );
or \U$56612 ( \56955 , \56950 , \56954 );
or \U$56613 ( \56956 , \56953 , \3918 );
nand \U$56614 ( \56957 , \56955 , \56956 );
and \U$56615 ( \56958 , \4203 , RI9870948_96);
and \U$56616 ( \56959 , RI9870858_94, \4201 );
nor \U$56617 ( \56960 , \56958 , \56959 );
and \U$56618 ( \56961 , \56960 , \4207 );
not \U$56619 ( \56962 , \56960 );
and \U$56620 ( \56963 , \56962 , \3923 );
nor \U$56621 ( \56964 , \56961 , \56963 );
xor \U$56622 ( \56965 , \56957 , \56964 );
not \U$56623 ( \56966 , \4519 );
and \U$56624 ( \56967 , \4710 , RI986fb38_66);
and \U$56625 ( \56968 , RI986fc28_68, \4708 );
nor \U$56626 ( \56969 , \56967 , \56968 );
not \U$56627 ( \56970 , \56969 );
or \U$56628 ( \56971 , \56966 , \56970 );
or \U$56629 ( \56972 , \56969 , \4519 );
nand \U$56630 ( \56973 , \56971 , \56972 );
and \U$56631 ( \56974 , \56965 , \56973 );
and \U$56632 ( \56975 , \56957 , \56964 );
or \U$56633 ( \56976 , \56974 , \56975 );
and \U$56634 ( \56977 , \56949 , \56976 );
and \U$56635 ( \56978 , \56923 , \56948 );
or \U$56636 ( \56979 , \56977 , \56978 );
and \U$56637 ( \56980 , \13045 , RI986eb48_32);
and \U$56638 ( \56981 , RI986ea58_30, \13043 );
nor \U$56639 ( \56982 , \56980 , \56981 );
and \U$56640 ( \56983 , \56982 , \13047 );
not \U$56641 ( \56984 , \56982 );
and \U$56642 ( \56985 , \56984 , \12619 );
nor \U$56643 ( \56986 , \56983 , \56985 );
and \U$56644 ( \56987 , \11696 , RI9871758_126);
and \U$56645 ( \56988 , RI9871848_128, \11694 );
nor \U$56646 ( \56989 , \56987 , \56988 );
and \U$56647 ( \56990 , \56989 , \10965 );
not \U$56648 ( \56991 , \56989 );
and \U$56649 ( \56992 , \56991 , \11702 );
nor \U$56650 ( \56993 , \56990 , \56992 );
xor \U$56651 ( \56994 , \56986 , \56993 );
and \U$56652 ( \56995 , \12293 , RI9871578_122);
and \U$56653 ( \56996 , RI9871668_124, \12291 );
nor \U$56654 ( \56997 , \56995 , \56996 );
and \U$56655 ( \56998 , \56997 , \11687 );
not \U$56656 ( \56999 , \56997 );
and \U$56657 ( \57000 , \56999 , \11686 );
nor \U$56658 ( \57001 , \56998 , \57000 );
and \U$56659 ( \57002 , \56994 , \57001 );
and \U$56660 ( \57003 , \56986 , \56993 );
or \U$56661 ( \57004 , \57002 , \57003 );
and \U$56662 ( \57005 , \14937 , RI986ef08_40);
and \U$56663 ( \57006 , RI986ee18_38, \14935 );
nor \U$56664 ( \57007 , \57005 , \57006 );
and \U$56665 ( \57008 , \57007 , \14539 );
not \U$56666 ( \57009 , \57007 );
and \U$56667 ( \57010 , \57009 , \14538 );
nor \U$56668 ( \57011 , \57008 , \57010 );
not \U$56669 ( \57012 , RI9873558_190);
and \U$56670 ( \57013 , \15780 , RI986ec38_34);
and \U$56671 ( \57014 , RI986ed28_36, RI9873648_192);
nor \U$56672 ( \57015 , \57013 , \57014 );
not \U$56673 ( \57016 , \57015 );
or \U$56674 ( \57017 , \57012 , \57016 );
or \U$56675 ( \57018 , \57015 , RI9873558_190);
nand \U$56676 ( \57019 , \57017 , \57018 );
xor \U$56677 ( \57020 , \57011 , \57019 );
and \U$56678 ( \57021 , \13882 , RI986e968_28);
and \U$56679 ( \57022 , RI986e878_26, \13880 );
nor \U$56680 ( \57023 , \57021 , \57022 );
and \U$56681 ( \57024 , \57023 , \13358 );
not \U$56682 ( \57025 , \57023 );
and \U$56683 ( \57026 , \57025 , \13359 );
nor \U$56684 ( \57027 , \57024 , \57026 );
and \U$56685 ( \57028 , \57020 , \57027 );
and \U$56686 ( \57029 , \57011 , \57019 );
or \U$56687 ( \57030 , \57028 , \57029 );
xor \U$56688 ( \57031 , \57004 , \57030 );
and \U$56689 ( \57032 , \9237 , RI98710c8_112);
and \U$56690 ( \57033 , RI9870d08_104, \9235 );
nor \U$56691 ( \57034 , \57032 , \57033 );
and \U$56692 ( \57035 , \57034 , \9241 );
not \U$56693 ( \57036 , \57034 );
and \U$56694 ( \57037 , \57036 , \8836 );
nor \U$56695 ( \57038 , \57035 , \57037 );
and \U$56696 ( \57039 , \9505 , RI98712a8_116);
and \U$56697 ( \57040 , RI98711b8_114, \9503 );
nor \U$56698 ( \57041 , \57039 , \57040 );
and \U$56699 ( \57042 , \57041 , \9510 );
not \U$56700 ( \57043 , \57041 );
and \U$56701 ( \57044 , \57043 , \9513 );
nor \U$56702 ( \57045 , \57042 , \57044 );
xor \U$56703 ( \57046 , \57038 , \57045 );
and \U$56704 ( \57047 , \10424 , RI9871398_118);
and \U$56705 ( \57048 , RI9871488_120, \10422 );
nor \U$56706 ( \57049 , \57047 , \57048 );
and \U$56707 ( \57050 , \57049 , \9840 );
not \U$56708 ( \57051 , \57049 );
and \U$56709 ( \57052 , \57051 , \10428 );
nor \U$56710 ( \57053 , \57050 , \57052 );
and \U$56711 ( \57054 , \57046 , \57053 );
and \U$56712 ( \57055 , \57038 , \57045 );
or \U$56713 ( \57056 , \57054 , \57055 );
and \U$56714 ( \57057 , \57031 , \57056 );
and \U$56715 ( \57058 , \57004 , \57030 );
or \U$56716 ( \57059 , \57057 , \57058 );
xor \U$56717 ( \57060 , \56979 , \57059 );
xor \U$56718 ( \57061 , \56665 , \56672 );
xor \U$56719 ( \57062 , \57061 , \56681 );
nand \U$56720 ( \57063 , RI9870498_86, \2272 );
and \U$56721 ( \57064 , \57063 , \2030 );
not \U$56722 ( \57065 , \57063 );
and \U$56723 ( \57066 , \57065 , \2031 );
nor \U$56724 ( \57067 , \57064 , \57066 );
xor \U$56725 ( \57068 , \57062 , \57067 );
xor \U$56726 ( \57069 , \56794 , \56802 );
xor \U$56727 ( \57070 , \57069 , \56811 );
and \U$56728 ( \57071 , \57068 , \57070 );
and \U$56729 ( \57072 , \57062 , \57067 );
or \U$56730 ( \57073 , \57071 , \57072 );
and \U$56731 ( \57074 , \57060 , \57073 );
and \U$56732 ( \57075 , \56979 , \57059 );
or \U$56733 ( \57076 , \57074 , \57075 );
xor \U$56734 ( \57077 , \56898 , \57076 );
xor \U$56735 ( \57078 , \56692 , \56699 );
xor \U$56736 ( \57079 , \57078 , \56707 );
xor \U$56737 ( \57080 , \56720 , \56727 );
xor \U$56738 ( \57081 , \57080 , \56735 );
and \U$56739 ( \57082 , \57079 , \57081 );
xor \U$56740 ( \57083 , \56640 , \56647 );
xor \U$56741 ( \57084 , \57083 , \56655 );
xor \U$56742 ( \57085 , \56720 , \56727 );
xor \U$56743 ( \57086 , \57085 , \56735 );
and \U$56744 ( \57087 , \57084 , \57086 );
and \U$56745 ( \57088 , \57079 , \57084 );
or \U$56746 ( \57089 , \57082 , \57087 , \57088 );
xor \U$56747 ( \57090 , \56842 , \56844 );
xor \U$56748 ( \57091 , \57089 , \57090 );
xor \U$56749 ( \57092 , \56426 , \56433 );
xor \U$56750 ( \57093 , \57092 , \56441 );
xor \U$56751 ( \57094 , \56830 , \56835 );
xor \U$56752 ( \57095 , \57093 , \57094 );
and \U$56753 ( \57096 , \57091 , \57095 );
and \U$56754 ( \57097 , \57089 , \57090 );
or \U$56755 ( \57098 , \57096 , \57097 );
and \U$56756 ( \57099 , \57077 , \57098 );
and \U$56757 ( \57100 , \56898 , \57076 );
or \U$56758 ( \57101 , \57099 , \57100 );
xor \U$56759 ( \57102 , \56322 , \56324 );
xor \U$56760 ( \57103 , \57102 , \56335 );
xor \U$56761 ( \57104 , \57101 , \57103 );
xor \U$56762 ( \57105 , \56444 , \56470 );
xor \U$56763 ( \57106 , \57105 , \56496 );
xor \U$56764 ( \57107 , \56840 , \56845 );
xor \U$56765 ( \57108 , \57107 , \56850 );
and \U$56766 ( \57109 , \57106 , \57108 );
xor \U$56767 ( \57110 , \56327 , \56329 );
xor \U$56768 ( \57111 , \57110 , \56332 );
xor \U$56769 ( \57112 , \56623 , \56628 );
xor \U$56770 ( \57113 , \57111 , \57112 );
xor \U$56771 ( \57114 , \56840 , \56845 );
xor \U$56772 ( \57115 , \57114 , \56850 );
and \U$56773 ( \57116 , \57113 , \57115 );
and \U$56774 ( \57117 , \57106 , \57113 );
or \U$56775 ( \57118 , \57109 , \57116 , \57117 );
and \U$56776 ( \57119 , \57104 , \57118 );
and \U$56777 ( \57120 , \57101 , \57103 );
or \U$56778 ( \57121 , \57119 , \57120 );
xor \U$56779 ( \57122 , \56886 , \57121 );
xor \U$56780 ( \57123 , \56957 , \56964 );
xor \U$56781 ( \57124 , \57123 , \56973 );
xor \U$56782 ( \57125 , \56930 , \56937 );
xor \U$56783 ( \57126 , \57125 , \56945 );
and \U$56784 ( \57127 , \57124 , \57126 );
xor \U$56785 ( \57128 , \56905 , \56912 );
xor \U$56786 ( \57129 , \57128 , \56920 );
xor \U$56787 ( \57130 , \56930 , \56937 );
xor \U$56788 ( \57131 , \57130 , \56945 );
and \U$56789 ( \57132 , \57129 , \57131 );
and \U$56790 ( \57133 , \57124 , \57129 );
or \U$56791 ( \57134 , \57127 , \57132 , \57133 );
xor \U$56792 ( \57135 , \56765 , \56772 );
xor \U$56793 ( \57136 , \57135 , \56780 );
xor \U$56794 ( \57137 , \57134 , \57136 );
xor \U$56795 ( \57138 , \57011 , \57019 );
xor \U$56796 ( \57139 , \57138 , \57027 );
xor \U$56797 ( \57140 , \57038 , \57045 );
xor \U$56798 ( \57141 , \57140 , \57053 );
xor \U$56799 ( \57142 , \57139 , \57141 );
xor \U$56800 ( \57143 , \56986 , \56993 );
xor \U$56801 ( \57144 , \57143 , \57001 );
and \U$56802 ( \57145 , \57142 , \57144 );
and \U$56803 ( \57146 , \57139 , \57141 );
or \U$56804 ( \57147 , \57145 , \57146 );
and \U$56805 ( \57148 , \57137 , \57147 );
and \U$56806 ( \57149 , \57134 , \57136 );
or \U$56807 ( \57150 , \57148 , \57149 );
and \U$56808 ( \57151 , \9505 , RI9870d08_104);
and \U$56809 ( \57152 , RI98712a8_116, \9503 );
nor \U$56810 ( \57153 , \57151 , \57152 );
and \U$56811 ( \57154 , \57153 , \9510 );
not \U$56812 ( \57155 , \57153 );
and \U$56813 ( \57156 , \57155 , \9513 );
nor \U$56814 ( \57157 , \57154 , \57156 );
and \U$56815 ( \57158 , \10424 , RI98711b8_114);
and \U$56816 ( \57159 , RI9871398_118, \10422 );
nor \U$56817 ( \57160 , \57158 , \57159 );
and \U$56818 ( \57161 , \57160 , \9840 );
not \U$56819 ( \57162 , \57160 );
and \U$56820 ( \57163 , \57162 , \10428 );
nor \U$56821 ( \57164 , \57161 , \57163 );
xor \U$56822 ( \57165 , \57157 , \57164 );
and \U$56823 ( \57166 , \11696 , RI9871488_120);
and \U$56824 ( \57167 , RI9871758_126, \11694 );
nor \U$56825 ( \57168 , \57166 , \57167 );
and \U$56826 ( \57169 , \57168 , \10965 );
not \U$56827 ( \57170 , \57168 );
and \U$56828 ( \57171 , \57170 , \11702 );
nor \U$56829 ( \57172 , \57169 , \57171 );
and \U$56830 ( \57173 , \57165 , \57172 );
and \U$56831 ( \57174 , \57157 , \57164 );
or \U$56832 ( \57175 , \57173 , \57174 );
not \U$56833 ( \57176 , RI9873558_190);
and \U$56834 ( \57177 , \15780 , RI986ee18_38);
and \U$56835 ( \57178 , RI986ec38_34, RI9873648_192);
nor \U$56836 ( \57179 , \57177 , \57178 );
not \U$56837 ( \57180 , \57179 );
or \U$56838 ( \57181 , \57176 , \57180 );
or \U$56839 ( \57182 , \57179 , RI9873558_190);
nand \U$56840 ( \57183 , \57181 , \57182 );
xor \U$56841 ( \57184 , \57183 , \2263 );
and \U$56842 ( \57185 , \14937 , RI986e878_26);
and \U$56843 ( \57186 , RI986ef08_40, \14935 );
nor \U$56844 ( \57187 , \57185 , \57186 );
and \U$56845 ( \57188 , \57187 , \14539 );
not \U$56846 ( \57189 , \57187 );
and \U$56847 ( \57190 , \57189 , \14538 );
nor \U$56848 ( \57191 , \57188 , \57190 );
and \U$56849 ( \57192 , \57184 , \57191 );
and \U$56850 ( \57193 , \57183 , \2263 );
or \U$56851 ( \57194 , \57192 , \57193 );
xor \U$56852 ( \57195 , \57175 , \57194 );
and \U$56853 ( \57196 , \12293 , RI9871848_128);
and \U$56854 ( \57197 , RI9871578_122, \12291 );
nor \U$56855 ( \57198 , \57196 , \57197 );
and \U$56856 ( \57199 , \57198 , \11687 );
not \U$56857 ( \57200 , \57198 );
and \U$56858 ( \57201 , \57200 , \11686 );
nor \U$56859 ( \57202 , \57199 , \57201 );
and \U$56860 ( \57203 , \13045 , RI9871668_124);
and \U$56861 ( \57204 , RI986eb48_32, \13043 );
nor \U$56862 ( \57205 , \57203 , \57204 );
and \U$56863 ( \57206 , \57205 , \13047 );
not \U$56864 ( \57207 , \57205 );
and \U$56865 ( \57208 , \57207 , \12619 );
nor \U$56866 ( \57209 , \57206 , \57208 );
xor \U$56867 ( \57210 , \57202 , \57209 );
and \U$56868 ( \57211 , \13882 , RI986ea58_30);
and \U$56869 ( \57212 , RI986e968_28, \13880 );
nor \U$56870 ( \57213 , \57211 , \57212 );
and \U$56871 ( \57214 , \57213 , \13358 );
not \U$56872 ( \57215 , \57213 );
and \U$56873 ( \57216 , \57215 , \13359 );
nor \U$56874 ( \57217 , \57214 , \57216 );
and \U$56875 ( \57218 , \57210 , \57217 );
and \U$56876 ( \57219 , \57202 , \57209 );
or \U$56877 ( \57220 , \57218 , \57219 );
and \U$56878 ( \57221 , \57195 , \57220 );
and \U$56879 ( \57222 , \57175 , \57194 );
or \U$56880 ( \57223 , \57221 , \57222 );
not \U$56881 ( \57224 , \2935 );
and \U$56882 ( \57225 , \3254 , RI98703a8_84);
and \U$56883 ( \57226 , RI98702b8_82, \3252 );
nor \U$56884 ( \57227 , \57225 , \57226 );
not \U$56885 ( \57228 , \57227 );
or \U$56886 ( \57229 , \57224 , \57228 );
or \U$56887 ( \57230 , \57227 , \3406 );
nand \U$56888 ( \57231 , \57229 , \57230 );
and \U$56889 ( \57232 , \2464 , RI9870498_86);
and \U$56890 ( \57233 , RI9870588_88, \2462 );
nor \U$56891 ( \57234 , \57232 , \57233 );
and \U$56892 ( \57235 , \57234 , \2468 );
not \U$56893 ( \57236 , \57234 );
and \U$56894 ( \57237 , \57236 , \2263 );
nor \U$56895 ( \57238 , \57235 , \57237 );
xor \U$56896 ( \57239 , \57231 , \57238 );
not \U$56897 ( \57240 , \3412 );
and \U$56898 ( \57241 , \3683 , RI98702b8_82);
and \U$56899 ( \57242 , RI9870768_92, \3681 );
nor \U$56900 ( \57243 , \57241 , \57242 );
not \U$56901 ( \57244 , \57243 );
or \U$56902 ( \57245 , \57240 , \57244 );
or \U$56903 ( \57246 , \57243 , \3412 );
nand \U$56904 ( \57247 , \57245 , \57246 );
nand \U$56905 ( \57248 , RI9870498_86, \2462 );
and \U$56906 ( \57249 , \57248 , \2468 );
not \U$56907 ( \57250 , \57248 );
and \U$56908 ( \57251 , \57250 , \2263 );
nor \U$56909 ( \57252 , \57249 , \57251 );
xor \U$56910 ( \57253 , \57247 , \57252 );
not \U$56911 ( \57254 , \2935 );
and \U$56912 ( \57255 , \3254 , RI9870588_88);
and \U$56913 ( \57256 , RI98703a8_84, \3252 );
nor \U$56914 ( \57257 , \57255 , \57256 );
not \U$56915 ( \57258 , \57257 );
or \U$56916 ( \57259 , \57254 , \57258 );
or \U$56917 ( \57260 , \57257 , \2935 );
nand \U$56918 ( \57261 , \57259 , \57260 );
and \U$56919 ( \57262 , \57253 , \57261 );
and \U$56920 ( \57263 , \57247 , \57252 );
or \U$56921 ( \57264 , \57262 , \57263 );
and \U$56922 ( \57265 , \57239 , \57264 );
and \U$56923 ( \57266 , \57231 , \57238 );
or \U$56924 ( \57267 , \57265 , \57266 );
xor \U$56925 ( \57268 , \57223 , \57267 );
and \U$56926 ( \57269 , \8486 , RI9870a38_98);
and \U$56927 ( \57270 , RI9870ee8_108, \8484 );
nor \U$56928 ( \57271 , \57269 , \57270 );
and \U$56929 ( \57272 , \57271 , \8050 );
not \U$56930 ( \57273 , \57271 );
and \U$56931 ( \57274 , \57273 , \8051 );
nor \U$56932 ( \57275 , \57272 , \57274 );
and \U$56933 ( \57276 , \7729 , RI9870b28_100);
and \U$56934 ( \57277 , RI9870df8_106, \7727 );
nor \U$56935 ( \57278 , \57276 , \57277 );
and \U$56936 ( \57279 , \57278 , \7480 );
not \U$56937 ( \57280 , \57278 );
and \U$56938 ( \57281 , \57280 , \7733 );
nor \U$56939 ( \57282 , \57279 , \57281 );
xor \U$56940 ( \57283 , \57275 , \57282 );
and \U$56941 ( \57284 , \9237 , RI9870c18_102);
and \U$56942 ( \57285 , RI98710c8_112, \9235 );
nor \U$56943 ( \57286 , \57284 , \57285 );
and \U$56944 ( \57287 , \57286 , \9241 );
not \U$56945 ( \57288 , \57286 );
and \U$56946 ( \57289 , \57288 , \8836 );
nor \U$56947 ( \57290 , \57287 , \57289 );
and \U$56948 ( \57291 , \57283 , \57290 );
and \U$56949 ( \57292 , \57275 , \57282 );
or \U$56950 ( \57293 , \57291 , \57292 );
and \U$56951 ( \57294 , \5318 , RI986fc28_68);
and \U$56952 ( \57295 , RI986fe08_72, \5316 );
nor \U$56953 ( \57296 , \57294 , \57295 );
and \U$56954 ( \57297 , \57296 , \5052 );
not \U$56955 ( \57298 , \57296 );
and \U$56956 ( \57299 , \57298 , \5322 );
nor \U$56957 ( \57300 , \57297 , \57299 );
and \U$56958 ( \57301 , \4203 , RI9870678_90);
and \U$56959 ( \57302 , RI9870948_96, \4201 );
nor \U$56960 ( \57303 , \57301 , \57302 );
and \U$56961 ( \57304 , \57303 , \4207 );
not \U$56962 ( \57305 , \57303 );
and \U$56963 ( \57306 , \57305 , \3922 );
nor \U$56964 ( \57307 , \57304 , \57306 );
xor \U$56965 ( \57308 , \57300 , \57307 );
not \U$56966 ( \57309 , \4519 );
and \U$56967 ( \57310 , \4710 , RI9870858_94);
and \U$56968 ( \57311 , RI986fb38_66, \4708 );
nor \U$56969 ( \57312 , \57310 , \57311 );
not \U$56970 ( \57313 , \57312 );
or \U$56971 ( \57314 , \57309 , \57313 );
or \U$56972 ( \57315 , \57312 , \4519 );
nand \U$56973 ( \57316 , \57314 , \57315 );
and \U$56974 ( \57317 , \57308 , \57316 );
and \U$56975 ( \57318 , \57300 , \57307 );
or \U$56976 ( \57319 , \57317 , \57318 );
xor \U$56977 ( \57320 , \57293 , \57319 );
and \U$56978 ( \57321 , \5881 , RI986fd18_70);
and \U$56979 ( \57322 , RI986ffe8_76, \5879 );
nor \U$56980 ( \57323 , \57321 , \57322 );
and \U$56981 ( \57324 , \57323 , \5594 );
not \U$56982 ( \57325 , \57323 );
and \U$56983 ( \57326 , \57325 , \5885 );
nor \U$56984 ( \57327 , \57324 , \57326 );
and \U$56985 ( \57328 , \6453 , RI986fef8_74);
and \U$56986 ( \57329 , RI98700d8_78, \6451 );
nor \U$56987 ( \57330 , \57328 , \57329 );
and \U$56988 ( \57331 , \57330 , \6190 );
not \U$56989 ( \57332 , \57330 );
and \U$56990 ( \57333 , \57332 , \6705 );
nor \U$56991 ( \57334 , \57331 , \57333 );
xor \U$56992 ( \57335 , \57327 , \57334 );
and \U$56993 ( \57336 , \7079 , RI98701c8_80);
and \U$56994 ( \57337 , RI9870fd8_110, \7077 );
nor \U$56995 ( \57338 , \57336 , \57337 );
and \U$56996 ( \57339 , \57338 , \6710 );
not \U$56997 ( \57340 , \57338 );
and \U$56998 ( \57341 , \57340 , \6709 );
nor \U$56999 ( \57342 , \57339 , \57341 );
and \U$57000 ( \57343 , \57335 , \57342 );
and \U$57001 ( \57344 , \57327 , \57334 );
or \U$57002 ( \57345 , \57343 , \57344 );
and \U$57003 ( \57346 , \57320 , \57345 );
and \U$57004 ( \57347 , \57293 , \57319 );
or \U$57005 ( \57348 , \57346 , \57347 );
and \U$57006 ( \57349 , \57268 , \57348 );
and \U$57007 ( \57350 , \57223 , \57267 );
or \U$57008 ( \57351 , \57349 , \57350 );
xor \U$57009 ( \57352 , \57150 , \57351 );
xor \U$57010 ( \57353 , \56746 , \2031 );
xor \U$57011 ( \57354 , \57353 , \56754 );
xor \U$57012 ( \57355 , \57062 , \57067 );
xor \U$57013 ( \57356 , \57355 , \57070 );
and \U$57014 ( \57357 , \57354 , \57356 );
xor \U$57015 ( \57358 , \56720 , \56727 );
xor \U$57016 ( \57359 , \57358 , \56735 );
xor \U$57017 ( \57360 , \57079 , \57084 );
xor \U$57018 ( \57361 , \57359 , \57360 );
xor \U$57019 ( \57362 , \57062 , \57067 );
xor \U$57020 ( \57363 , \57362 , \57070 );
and \U$57021 ( \57364 , \57361 , \57363 );
and \U$57022 ( \57365 , \57354 , \57361 );
or \U$57023 ( \57366 , \57357 , \57364 , \57365 );
and \U$57024 ( \57367 , \57352 , \57366 );
and \U$57025 ( \57368 , \57150 , \57351 );
or \U$57026 ( \57369 , \57367 , \57368 );
xor \U$57027 ( \57370 , \56713 , \56786 );
xor \U$57028 ( \57371 , \57370 , \56824 );
xor \U$57029 ( \57372 , \57369 , \57371 );
xor \U$57030 ( \57373 , \56979 , \57059 );
xor \U$57031 ( \57374 , \57373 , \57073 );
xor \U$57032 ( \57375 , \56888 , \56890 );
xor \U$57033 ( \57376 , \57375 , \56895 );
and \U$57034 ( \57377 , \57374 , \57376 );
xor \U$57035 ( \57378 , \57089 , \57090 );
xor \U$57036 ( \57379 , \57378 , \57095 );
xor \U$57037 ( \57380 , \56888 , \56890 );
xor \U$57038 ( \57381 , \57380 , \56895 );
and \U$57039 ( \57382 , \57379 , \57381 );
and \U$57040 ( \57383 , \57374 , \57379 );
or \U$57041 ( \57384 , \57377 , \57382 , \57383 );
and \U$57042 ( \57385 , \57372 , \57384 );
and \U$57043 ( \57386 , \57369 , \57371 );
or \U$57044 ( \57387 , \57385 , \57386 );
xor \U$57045 ( \57388 , \56898 , \57076 );
xor \U$57046 ( \57389 , \57388 , \57098 );
xor \U$57047 ( \57390 , \56840 , \56845 );
xor \U$57048 ( \57391 , \57390 , \56850 );
xor \U$57049 ( \57392 , \57106 , \57113 );
xor \U$57050 ( \57393 , \57391 , \57392 );
and \U$57051 ( \57394 , \57389 , \57393 );
xor \U$57052 ( \57395 , \57387 , \57394 );
xor \U$57053 ( \57396 , \56608 , \56610 );
xor \U$57054 ( \57397 , \57396 , \56615 );
xor \U$57055 ( \57398 , \56871 , \56876 );
xor \U$57056 ( \57399 , \57397 , \57398 );
and \U$57057 ( \57400 , \57395 , \57399 );
and \U$57058 ( \57401 , \57387 , \57394 );
or \U$57059 ( \57402 , \57400 , \57401 );
xnor \U$57060 ( \57403 , \57122 , \57402 );
not \U$57061 ( \57404 , \57403 );
xor \U$57062 ( \57405 , \56338 , \56536 );
xor \U$57063 ( \57406 , \57405 , \56551 );
xor \U$57064 ( \57407 , \56618 , \56620 );
xor \U$57065 ( \57408 , \57407 , \56856 );
xor \U$57066 ( \57409 , \57406 , \57408 );
not \U$57067 ( \57410 , \57409 );
and \U$57068 ( \57411 , \57404 , \57410 );
and \U$57069 ( \57412 , \57403 , \57409 );
nor \U$57070 ( \57413 , \57411 , \57412 );
xor \U$57071 ( \57414 , \57387 , \57394 );
xor \U$57072 ( \57415 , \57414 , \57399 );
xor \U$57073 ( \57416 , \57101 , \57103 );
xor \U$57074 ( \57417 , \57416 , \57118 );
xor \U$57075 ( \57418 , \57415 , \57417 );
xor \U$57076 ( \57419 , \57389 , \57393 );
not \U$57077 ( \57420 , \57419 );
xor \U$57078 ( \57421 , \57369 , \57371 );
xor \U$57079 ( \57422 , \57421 , \57384 );
not \U$57080 ( \57423 , \57422 );
or \U$57081 ( \57424 , \57420 , \57423 );
or \U$57082 ( \57425 , \57422 , \57419 );
xor \U$57083 ( \57426 , \57231 , \57238 );
xor \U$57084 ( \57427 , \57426 , \57264 );
xor \U$57085 ( \57428 , \57175 , \57194 );
xor \U$57086 ( \57429 , \57428 , \57220 );
and \U$57087 ( \57430 , \57427 , \57429 );
xor \U$57088 ( \57431 , \57293 , \57319 );
xor \U$57089 ( \57432 , \57431 , \57345 );
xor \U$57090 ( \57433 , \57175 , \57194 );
xor \U$57091 ( \57434 , \57433 , \57220 );
and \U$57092 ( \57435 , \57432 , \57434 );
and \U$57093 ( \57436 , \57427 , \57432 );
or \U$57094 ( \57437 , \57430 , \57435 , \57436 );
and \U$57095 ( \57438 , \7079 , RI98700d8_78);
and \U$57096 ( \57439 , RI98701c8_80, \7077 );
nor \U$57097 ( \57440 , \57438 , \57439 );
and \U$57098 ( \57441 , \57440 , \6710 );
not \U$57099 ( \57442 , \57440 );
and \U$57100 ( \57443 , \57442 , \6709 );
nor \U$57101 ( \57444 , \57441 , \57443 );
and \U$57102 ( \57445 , \7729 , RI9870fd8_110);
and \U$57103 ( \57446 , RI9870b28_100, \7727 );
nor \U$57104 ( \57447 , \57445 , \57446 );
and \U$57105 ( \57448 , \57447 , \7480 );
not \U$57106 ( \57449 , \57447 );
and \U$57107 ( \57450 , \57449 , \7733 );
nor \U$57108 ( \57451 , \57448 , \57450 );
xor \U$57109 ( \57452 , \57444 , \57451 );
and \U$57110 ( \57453 , \8486 , RI9870df8_106);
and \U$57111 ( \57454 , RI9870a38_98, \8484 );
nor \U$57112 ( \57455 , \57453 , \57454 );
and \U$57113 ( \57456 , \57455 , \8050 );
not \U$57114 ( \57457 , \57455 );
and \U$57115 ( \57458 , \57457 , \8051 );
nor \U$57116 ( \57459 , \57456 , \57458 );
and \U$57117 ( \57460 , \57452 , \57459 );
and \U$57118 ( \57461 , \57444 , \57451 );
or \U$57119 ( \57462 , \57460 , \57461 );
not \U$57120 ( \57463 , \3412 );
and \U$57121 ( \57464 , \3683 , RI98703a8_84);
and \U$57122 ( \57465 , RI98702b8_82, \3681 );
nor \U$57123 ( \57466 , \57464 , \57465 );
not \U$57124 ( \57467 , \57466 );
or \U$57125 ( \57468 , \57463 , \57467 );
or \U$57126 ( \57469 , \57466 , \3412 );
nand \U$57127 ( \57470 , \57468 , \57469 );
and \U$57128 ( \57471 , \4203 , RI9870768_92);
and \U$57129 ( \57472 , RI9870678_90, \4201 );
nor \U$57130 ( \57473 , \57471 , \57472 );
and \U$57131 ( \57474 , \57473 , \4207 );
not \U$57132 ( \57475 , \57473 );
and \U$57133 ( \57476 , \57475 , \3923 );
nor \U$57134 ( \57477 , \57474 , \57476 );
xor \U$57135 ( \57478 , \57470 , \57477 );
not \U$57136 ( \57479 , \4519 );
and \U$57137 ( \57480 , \4710 , RI9870948_96);
and \U$57138 ( \57481 , RI9870858_94, \4708 );
nor \U$57139 ( \57482 , \57480 , \57481 );
not \U$57140 ( \57483 , \57482 );
or \U$57141 ( \57484 , \57479 , \57483 );
or \U$57142 ( \57485 , \57482 , \4521 );
nand \U$57143 ( \57486 , \57484 , \57485 );
and \U$57144 ( \57487 , \57478 , \57486 );
and \U$57145 ( \57488 , \57470 , \57477 );
or \U$57146 ( \57489 , \57487 , \57488 );
xor \U$57147 ( \57490 , \57462 , \57489 );
and \U$57148 ( \57491 , \5318 , RI986fb38_66);
and \U$57149 ( \57492 , RI986fc28_68, \5316 );
nor \U$57150 ( \57493 , \57491 , \57492 );
and \U$57151 ( \57494 , \57493 , \5052 );
not \U$57152 ( \57495 , \57493 );
and \U$57153 ( \57496 , \57495 , \5322 );
nor \U$57154 ( \57497 , \57494 , \57496 );
and \U$57155 ( \57498 , \5881 , RI986fe08_72);
and \U$57156 ( \57499 , RI986fd18_70, \5879 );
nor \U$57157 ( \57500 , \57498 , \57499 );
and \U$57158 ( \57501 , \57500 , \5594 );
not \U$57159 ( \57502 , \57500 );
and \U$57160 ( \57503 , \57502 , \5885 );
nor \U$57161 ( \57504 , \57501 , \57503 );
xor \U$57162 ( \57505 , \57497 , \57504 );
and \U$57163 ( \57506 , \6453 , RI986ffe8_76);
and \U$57164 ( \57507 , RI986fef8_74, \6451 );
nor \U$57165 ( \57508 , \57506 , \57507 );
and \U$57166 ( \57509 , \57508 , \6190 );
not \U$57167 ( \57510 , \57508 );
and \U$57168 ( \57511 , \57510 , \6180 );
nor \U$57169 ( \57512 , \57509 , \57511 );
and \U$57170 ( \57513 , \57505 , \57512 );
and \U$57171 ( \57514 , \57497 , \57504 );
or \U$57172 ( \57515 , \57513 , \57514 );
and \U$57173 ( \57516 , \57490 , \57515 );
and \U$57174 ( \57517 , \57462 , \57489 );
or \U$57175 ( \57518 , \57516 , \57517 );
and \U$57176 ( \57519 , \9237 , RI9870ee8_108);
and \U$57177 ( \57520 , RI9870c18_102, \9235 );
nor \U$57178 ( \57521 , \57519 , \57520 );
and \U$57179 ( \57522 , \57521 , \9241 );
not \U$57180 ( \57523 , \57521 );
and \U$57181 ( \57524 , \57523 , \8836 );
nor \U$57182 ( \57525 , \57522 , \57524 );
and \U$57183 ( \57526 , \9505 , RI98710c8_112);
and \U$57184 ( \57527 , RI9870d08_104, \9503 );
nor \U$57185 ( \57528 , \57526 , \57527 );
and \U$57186 ( \57529 , \57528 , \9510 );
not \U$57187 ( \57530 , \57528 );
and \U$57188 ( \57531 , \57530 , \9513 );
nor \U$57189 ( \57532 , \57529 , \57531 );
xor \U$57190 ( \57533 , \57525 , \57532 );
and \U$57191 ( \57534 , \10424 , RI98712a8_116);
and \U$57192 ( \57535 , RI98711b8_114, \10422 );
nor \U$57193 ( \57536 , \57534 , \57535 );
and \U$57194 ( \57537 , \57536 , \9840 );
not \U$57195 ( \57538 , \57536 );
and \U$57196 ( \57539 , \57538 , \10428 );
nor \U$57197 ( \57540 , \57537 , \57539 );
and \U$57198 ( \57541 , \57533 , \57540 );
and \U$57199 ( \57542 , \57525 , \57532 );
or \U$57200 ( \57543 , \57541 , \57542 );
and \U$57201 ( \57544 , \15780 , RI986ef08_40);
and \U$57202 ( \57545 , RI986ee18_38, RI9873648_192);
nor \U$57203 ( \57546 , \57544 , \57545 );
not \U$57204 ( \57547 , \57546 );
not \U$57205 ( \57548 , RI9873558_190);
and \U$57206 ( \57549 , \57547 , \57548 );
and \U$57207 ( \57550 , \57546 , RI9873558_190);
nor \U$57208 ( \57551 , \57549 , \57550 );
and \U$57209 ( \57552 , \14937 , RI986e968_28);
and \U$57210 ( \57553 , RI986e878_26, \14935 );
nor \U$57211 ( \57554 , \57552 , \57553 );
and \U$57212 ( \57555 , \57554 , \14538 );
not \U$57213 ( \57556 , \57554 );
and \U$57214 ( \57557 , \57556 , \14539 );
nor \U$57215 ( \57558 , \57555 , \57557 );
xor \U$57216 ( \57559 , \57551 , \57558 );
and \U$57217 ( \57560 , \13882 , RI986eb48_32);
and \U$57218 ( \57561 , RI986ea58_30, \13880 );
nor \U$57219 ( \57562 , \57560 , \57561 );
and \U$57220 ( \57563 , \57562 , \13359 );
not \U$57221 ( \57564 , \57562 );
and \U$57222 ( \57565 , \57564 , \13358 );
nor \U$57223 ( \57566 , \57563 , \57565 );
and \U$57224 ( \57567 , \57559 , \57566 );
and \U$57225 ( \57568 , \57551 , \57558 );
nor \U$57226 ( \57569 , \57567 , \57568 );
xor \U$57227 ( \57570 , \57543 , \57569 );
and \U$57228 ( \57571 , \12293 , RI9871758_126);
and \U$57229 ( \57572 , RI9871848_128, \12291 );
nor \U$57230 ( \57573 , \57571 , \57572 );
and \U$57231 ( \57574 , \57573 , \11687 );
not \U$57232 ( \57575 , \57573 );
and \U$57233 ( \57576 , \57575 , \11686 );
nor \U$57234 ( \57577 , \57574 , \57576 );
and \U$57235 ( \57578 , \11696 , RI9871398_118);
and \U$57236 ( \57579 , RI9871488_120, \11694 );
nor \U$57237 ( \57580 , \57578 , \57579 );
and \U$57238 ( \57581 , \57580 , \10965 );
not \U$57239 ( \57582 , \57580 );
and \U$57240 ( \57583 , \57582 , \11702 );
nor \U$57241 ( \57584 , \57581 , \57583 );
xor \U$57242 ( \57585 , \57577 , \57584 );
and \U$57243 ( \57586 , \13045 , RI9871578_122);
and \U$57244 ( \57587 , RI9871668_124, \13043 );
nor \U$57245 ( \57588 , \57586 , \57587 );
and \U$57246 ( \57589 , \57588 , \13047 );
not \U$57247 ( \57590 , \57588 );
and \U$57248 ( \57591 , \57590 , \12619 );
nor \U$57249 ( \57592 , \57589 , \57591 );
and \U$57250 ( \57593 , \57585 , \57592 );
and \U$57251 ( \57594 , \57577 , \57584 );
or \U$57252 ( \57595 , \57593 , \57594 );
and \U$57253 ( \57596 , \57570 , \57595 );
and \U$57254 ( \57597 , \57543 , \57569 );
or \U$57255 ( \57598 , \57596 , \57597 );
xor \U$57256 ( \57599 , \57518 , \57598 );
xor \U$57257 ( \57600 , \57247 , \57252 );
xor \U$57258 ( \57601 , \57600 , \57261 );
xor \U$57259 ( \57602 , \57327 , \57334 );
xor \U$57260 ( \57603 , \57602 , \57342 );
and \U$57261 ( \57604 , \57601 , \57603 );
xor \U$57262 ( \57605 , \57300 , \57307 );
xor \U$57263 ( \57606 , \57605 , \57316 );
xor \U$57264 ( \57607 , \57327 , \57334 );
xor \U$57265 ( \57608 , \57607 , \57342 );
and \U$57266 ( \57609 , \57606 , \57608 );
and \U$57267 ( \57610 , \57601 , \57606 );
or \U$57268 ( \57611 , \57604 , \57609 , \57610 );
and \U$57269 ( \57612 , \57599 , \57611 );
and \U$57270 ( \57613 , \57518 , \57598 );
or \U$57271 ( \57614 , \57612 , \57613 );
xor \U$57272 ( \57615 , \57437 , \57614 );
xor \U$57273 ( \57616 , \57157 , \57164 );
xor \U$57274 ( \57617 , \57616 , \57172 );
xor \U$57275 ( \57618 , \57275 , \57282 );
xor \U$57276 ( \57619 , \57618 , \57290 );
and \U$57277 ( \57620 , \57617 , \57619 );
xor \U$57278 ( \57621 , \57202 , \57209 );
xor \U$57279 ( \57622 , \57621 , \57217 );
xor \U$57280 ( \57623 , \57275 , \57282 );
xor \U$57281 ( \57624 , \57623 , \57290 );
and \U$57282 ( \57625 , \57622 , \57624 );
and \U$57283 ( \57626 , \57617 , \57622 );
or \U$57284 ( \57627 , \57620 , \57625 , \57626 );
xor \U$57285 ( \57628 , \57139 , \57141 );
xor \U$57286 ( \57629 , \57628 , \57144 );
and \U$57287 ( \57630 , \57627 , \57629 );
xor \U$57288 ( \57631 , \56930 , \56937 );
xor \U$57289 ( \57632 , \57631 , \56945 );
xor \U$57290 ( \57633 , \57124 , \57129 );
xor \U$57291 ( \57634 , \57632 , \57633 );
xor \U$57292 ( \57635 , \57139 , \57141 );
xor \U$57293 ( \57636 , \57635 , \57144 );
and \U$57294 ( \57637 , \57634 , \57636 );
and \U$57295 ( \57638 , \57627 , \57634 );
or \U$57296 ( \57639 , \57630 , \57637 , \57638 );
and \U$57297 ( \57640 , \57615 , \57639 );
and \U$57298 ( \57641 , \57437 , \57614 );
or \U$57299 ( \57642 , \57640 , \57641 );
xor \U$57300 ( \57643 , \56923 , \56948 );
xor \U$57301 ( \57644 , \57643 , \56976 );
xor \U$57302 ( \57645 , \57004 , \57030 );
xor \U$57303 ( \57646 , \57645 , \57056 );
and \U$57304 ( \57647 , \57644 , \57646 );
xor \U$57305 ( \57648 , \57062 , \57067 );
xor \U$57306 ( \57649 , \57648 , \57070 );
xor \U$57307 ( \57650 , \57354 , \57361 );
xor \U$57308 ( \57651 , \57649 , \57650 );
xor \U$57309 ( \57652 , \57004 , \57030 );
xor \U$57310 ( \57653 , \57652 , \57056 );
and \U$57311 ( \57654 , \57651 , \57653 );
and \U$57312 ( \57655 , \57644 , \57651 );
or \U$57313 ( \57656 , \57647 , \57654 , \57655 );
xor \U$57314 ( \57657 , \57642 , \57656 );
xor \U$57315 ( \57658 , \56888 , \56890 );
xor \U$57316 ( \57659 , \57658 , \56895 );
xor \U$57317 ( \57660 , \57374 , \57379 );
xor \U$57318 ( \57661 , \57659 , \57660 );
and \U$57319 ( \57662 , \57657 , \57661 );
and \U$57320 ( \57663 , \57642 , \57656 );
or \U$57321 ( \57664 , \57662 , \57663 );
nand \U$57322 ( \57665 , \57425 , \57664 );
nand \U$57323 ( \57666 , \57424 , \57665 );
and \U$57324 ( \57667 , \57418 , \57666 );
and \U$57325 ( \57668 , \57415 , \57417 );
nor \U$57326 ( \57669 , \57667 , \57668 );
or \U$57327 ( \57670 , \57413 , \57669 );
xnor \U$57328 ( \57671 , \57669 , \57413 );
xor \U$57329 ( \57672 , \57642 , \57656 );
xor \U$57330 ( \57673 , \57672 , \57661 );
and \U$57331 ( \57674 , \7729 , RI98701c8_80);
and \U$57332 ( \57675 , RI9870fd8_110, \7727 );
nor \U$57333 ( \57676 , \57674 , \57675 );
and \U$57334 ( \57677 , \57676 , \7733 );
not \U$57335 ( \57678 , \57676 );
and \U$57336 ( \57679 , \57678 , \7480 );
nor \U$57337 ( \57680 , \57677 , \57679 );
and \U$57338 ( \57681 , \8486 , RI9870b28_100);
and \U$57339 ( \57682 , RI9870df8_106, \8484 );
nor \U$57340 ( \57683 , \57681 , \57682 );
and \U$57341 ( \57684 , \57683 , \8051 );
not \U$57342 ( \57685 , \57683 );
and \U$57343 ( \57686 , \57685 , \8050 );
nor \U$57344 ( \57687 , \57684 , \57686 );
or \U$57345 ( \57688 , \57680 , \57687 );
not \U$57346 ( \57689 , \57687 );
not \U$57347 ( \57690 , \57680 );
or \U$57348 ( \57691 , \57689 , \57690 );
and \U$57349 ( \57692 , \9237 , RI9870a38_98);
and \U$57350 ( \57693 , RI9870ee8_108, \9235 );
nor \U$57351 ( \57694 , \57692 , \57693 );
and \U$57352 ( \57695 , \57694 , \9241 );
not \U$57353 ( \57696 , \57694 );
and \U$57354 ( \57697 , \57696 , \8836 );
nor \U$57355 ( \57698 , \57695 , \57697 );
nand \U$57356 ( \57699 , \57691 , \57698 );
nand \U$57357 ( \57700 , \57688 , \57699 );
and \U$57358 ( \57701 , \5318 , RI9870858_94);
and \U$57359 ( \57702 , RI986fb38_66, \5316 );
nor \U$57360 ( \57703 , \57701 , \57702 );
and \U$57361 ( \57704 , \57703 , \5052 );
not \U$57362 ( \57705 , \57703 );
and \U$57363 ( \57706 , \57705 , \5322 );
nor \U$57364 ( \57707 , \57704 , \57706 );
and \U$57365 ( \57708 , \4203 , RI98702b8_82);
and \U$57366 ( \57709 , RI9870768_92, \4201 );
nor \U$57367 ( \57710 , \57708 , \57709 );
and \U$57368 ( \57711 , \57710 , \4207 );
not \U$57369 ( \57712 , \57710 );
and \U$57370 ( \57713 , \57712 , \3923 );
nor \U$57371 ( \57714 , \57711 , \57713 );
xor \U$57372 ( \57715 , \57707 , \57714 );
not \U$57373 ( \57716 , \4521 );
and \U$57374 ( \57717 , \4710 , RI9870678_90);
and \U$57375 ( \57718 , RI9870948_96, \4708 );
nor \U$57376 ( \57719 , \57717 , \57718 );
not \U$57377 ( \57720 , \57719 );
or \U$57378 ( \57721 , \57716 , \57720 );
or \U$57379 ( \57722 , \57719 , \4519 );
nand \U$57380 ( \57723 , \57721 , \57722 );
and \U$57381 ( \57724 , \57715 , \57723 );
and \U$57382 ( \57725 , \57707 , \57714 );
or \U$57383 ( \57726 , \57724 , \57725 );
xor \U$57384 ( \57727 , \57700 , \57726 );
and \U$57385 ( \57728 , \6453 , RI986fd18_70);
and \U$57386 ( \57729 , RI986ffe8_76, \6451 );
nor \U$57387 ( \57730 , \57728 , \57729 );
and \U$57388 ( \57731 , \57730 , \6705 );
not \U$57389 ( \57732 , \57730 );
and \U$57390 ( \57733 , \57732 , \6190 );
nor \U$57391 ( \57734 , \57731 , \57733 );
and \U$57392 ( \57735 , \7079 , RI986fef8_74);
and \U$57393 ( \57736 , RI98700d8_78, \7077 );
nor \U$57394 ( \57737 , \57735 , \57736 );
and \U$57395 ( \57738 , \57737 , \6709 );
not \U$57396 ( \57739 , \57737 );
and \U$57397 ( \57740 , \57739 , \6710 );
nor \U$57398 ( \57741 , \57738 , \57740 );
xor \U$57399 ( \57742 , \57734 , \57741 );
and \U$57400 ( \57743 , \5881 , RI986fc28_68);
and \U$57401 ( \57744 , RI986fe08_72, \5879 );
nor \U$57402 ( \57745 , \57743 , \57744 );
and \U$57403 ( \57746 , \57745 , \5885 );
not \U$57404 ( \57747 , \57745 );
and \U$57405 ( \57748 , \57747 , \5594 );
nor \U$57406 ( \57749 , \57746 , \57748 );
and \U$57407 ( \57750 , \57742 , \57749 );
and \U$57408 ( \57751 , \57734 , \57741 );
nor \U$57409 ( \57752 , \57750 , \57751 );
and \U$57410 ( \57753 , \57727 , \57752 );
and \U$57411 ( \57754 , \57700 , \57726 );
or \U$57412 ( \57755 , \57753 , \57754 );
not \U$57413 ( \57756 , RI9873558_190);
and \U$57414 ( \57757 , \15780 , RI986e878_26);
and \U$57415 ( \57758 , RI986ef08_40, RI9873648_192);
nor \U$57416 ( \57759 , \57757 , \57758 );
not \U$57417 ( \57760 , \57759 );
or \U$57418 ( \57761 , \57756 , \57760 );
or \U$57419 ( \57762 , \57759 , RI9873558_190);
nand \U$57420 ( \57763 , \57761 , \57762 );
xor \U$57421 ( \57764 , \57763 , \3406 );
and \U$57422 ( \57765 , \14937 , RI986ea58_30);
and \U$57423 ( \57766 , RI986e968_28, \14935 );
nor \U$57424 ( \57767 , \57765 , \57766 );
and \U$57425 ( \57768 , \57767 , \14539 );
not \U$57426 ( \57769 , \57767 );
and \U$57427 ( \57770 , \57769 , \14538 );
nor \U$57428 ( \57771 , \57768 , \57770 );
and \U$57429 ( \57772 , \57764 , \57771 );
and \U$57430 ( \57773 , \57763 , \3406 );
or \U$57431 ( \57774 , \57772 , \57773 );
not \U$57432 ( \57775 , \57774 );
and \U$57433 ( \57776 , \10424 , RI9870d08_104);
and \U$57434 ( \57777 , RI98712a8_116, \10422 );
nor \U$57435 ( \57778 , \57776 , \57777 );
and \U$57436 ( \57779 , \57778 , \10428 );
not \U$57437 ( \57780 , \57778 );
and \U$57438 ( \57781 , \57780 , \9840 );
nor \U$57439 ( \57782 , \57779 , \57781 );
and \U$57440 ( \57783 , \11696 , RI98711b8_114);
and \U$57441 ( \57784 , RI9871398_118, \11694 );
nor \U$57442 ( \57785 , \57783 , \57784 );
and \U$57443 ( \57786 , \57785 , \11702 );
not \U$57444 ( \57787 , \57785 );
and \U$57445 ( \57788 , \57787 , \10965 );
nor \U$57446 ( \57789 , \57786 , \57788 );
xor \U$57447 ( \57790 , \57782 , \57789 );
and \U$57448 ( \57791 , \9505 , RI9870c18_102);
and \U$57449 ( \57792 , RI98710c8_112, \9503 );
nor \U$57450 ( \57793 , \57791 , \57792 );
and \U$57451 ( \57794 , \57793 , \9513 );
not \U$57452 ( \57795 , \57793 );
and \U$57453 ( \57796 , \57795 , \9510 );
nor \U$57454 ( \57797 , \57794 , \57796 );
and \U$57455 ( \57798 , \57790 , \57797 );
and \U$57456 ( \57799 , \57782 , \57789 );
nor \U$57457 ( \57800 , \57798 , \57799 );
not \U$57458 ( \57801 , \57800 );
or \U$57459 ( \57802 , \57775 , \57801 );
or \U$57460 ( \57803 , \57800 , \57774 );
and \U$57461 ( \57804 , \13045 , RI9871848_128);
and \U$57462 ( \57805 , RI9871578_122, \13043 );
nor \U$57463 ( \57806 , \57804 , \57805 );
and \U$57464 ( \57807 , \57806 , \12619 );
not \U$57465 ( \57808 , \57806 );
and \U$57466 ( \57809 , \57808 , \13047 );
nor \U$57467 ( \57810 , \57807 , \57809 );
and \U$57468 ( \57811 , \13882 , RI9871668_124);
and \U$57469 ( \57812 , RI986eb48_32, \13880 );
nor \U$57470 ( \57813 , \57811 , \57812 );
and \U$57471 ( \57814 , \57813 , \13359 );
not \U$57472 ( \57815 , \57813 );
and \U$57473 ( \57816 , \57815 , \13358 );
nor \U$57474 ( \57817 , \57814 , \57816 );
xor \U$57475 ( \57818 , \57810 , \57817 );
and \U$57476 ( \57819 , \12293 , RI9871488_120);
and \U$57477 ( \57820 , RI9871758_126, \12291 );
nor \U$57478 ( \57821 , \57819 , \57820 );
and \U$57479 ( \57822 , \57821 , \11686 );
not \U$57480 ( \57823 , \57821 );
and \U$57481 ( \57824 , \57823 , \11687 );
nor \U$57482 ( \57825 , \57822 , \57824 );
and \U$57483 ( \57826 , \57818 , \57825 );
and \U$57484 ( \57827 , \57810 , \57817 );
nor \U$57485 ( \57828 , \57826 , \57827 );
nand \U$57486 ( \57829 , \57803 , \57828 );
nand \U$57487 ( \57830 , \57802 , \57829 );
xor \U$57488 ( \57831 , \57755 , \57830 );
not \U$57489 ( \57832 , \3406 );
and \U$57490 ( \57833 , \3254 , RI9870498_86);
and \U$57491 ( \57834 , RI9870588_88, \3252 );
nor \U$57492 ( \57835 , \57833 , \57834 );
not \U$57493 ( \57836 , \57835 );
or \U$57494 ( \57837 , \57832 , \57836 );
or \U$57495 ( \57838 , \57835 , \3406 );
nand \U$57496 ( \57839 , \57837 , \57838 );
xor \U$57497 ( \57840 , \57497 , \57504 );
xor \U$57498 ( \57841 , \57840 , \57512 );
and \U$57499 ( \57842 , \57839 , \57841 );
xor \U$57500 ( \57843 , \57470 , \57477 );
xor \U$57501 ( \57844 , \57843 , \57486 );
xor \U$57502 ( \57845 , \57497 , \57504 );
xor \U$57503 ( \57846 , \57845 , \57512 );
and \U$57504 ( \57847 , \57844 , \57846 );
and \U$57505 ( \57848 , \57839 , \57844 );
or \U$57506 ( \57849 , \57842 , \57847 , \57848 );
xor \U$57507 ( \57850 , \57831 , \57849 );
xor \U$57508 ( \57851 , \57444 , \57451 );
xor \U$57509 ( \57852 , \57851 , \57459 );
xor \U$57510 ( \57853 , \57525 , \57532 );
xor \U$57511 ( \57854 , \57853 , \57540 );
xor \U$57512 ( \57855 , \57852 , \57854 );
xor \U$57513 ( \57856 , \57577 , \57584 );
xor \U$57514 ( \57857 , \57856 , \57592 );
and \U$57515 ( \57858 , \57855 , \57857 );
and \U$57516 ( \57859 , \57852 , \57854 );
or \U$57517 ( \57860 , \57858 , \57859 );
xor \U$57518 ( \57861 , \57183 , \2263 );
xor \U$57519 ( \57862 , \57861 , \57191 );
xor \U$57520 ( \57863 , \57860 , \57862 );
xor \U$57521 ( \57864 , \57275 , \57282 );
xor \U$57522 ( \57865 , \57864 , \57290 );
xor \U$57523 ( \57866 , \57617 , \57622 );
xor \U$57524 ( \57867 , \57865 , \57866 );
xor \U$57525 ( \57868 , \57863 , \57867 );
and \U$57526 ( \57869 , \57850 , \57868 );
xor \U$57527 ( \57870 , \57462 , \57489 );
xor \U$57528 ( \57871 , \57870 , \57515 );
xor \U$57529 ( \57872 , \57543 , \57569 );
xor \U$57530 ( \57873 , \57872 , \57595 );
xor \U$57531 ( \57874 , \57327 , \57334 );
xor \U$57532 ( \57875 , \57874 , \57342 );
xor \U$57533 ( \57876 , \57601 , \57606 );
xor \U$57534 ( \57877 , \57875 , \57876 );
xor \U$57535 ( \57878 , \57873 , \57877 );
xor \U$57536 ( \57879 , \57871 , \57878 );
xor \U$57537 ( \57880 , \57860 , \57862 );
xor \U$57538 ( \57881 , \57880 , \57867 );
and \U$57539 ( \57882 , \57879 , \57881 );
and \U$57540 ( \57883 , \57850 , \57879 );
or \U$57541 ( \57884 , \57869 , \57882 , \57883 );
xor \U$57542 ( \57885 , \57700 , \57726 );
xor \U$57543 ( \57886 , \57885 , \57752 );
xor \U$57544 ( \57887 , \57852 , \57854 );
xor \U$57545 ( \57888 , \57887 , \57857 );
and \U$57546 ( \57889 , \57886 , \57888 );
xor \U$57547 ( \57890 , \57497 , \57504 );
xor \U$57548 ( \57891 , \57890 , \57512 );
xor \U$57549 ( \57892 , \57839 , \57844 );
xor \U$57550 ( \57893 , \57891 , \57892 );
xor \U$57551 ( \57894 , \57852 , \57854 );
xor \U$57552 ( \57895 , \57894 , \57857 );
and \U$57553 ( \57896 , \57893 , \57895 );
and \U$57554 ( \57897 , \57886 , \57893 );
or \U$57555 ( \57898 , \57889 , \57896 , \57897 );
not \U$57556 ( \57899 , \57898 );
xor \U$57557 ( \57900 , \57810 , \57817 );
xor \U$57558 ( \57901 , \57900 , \57825 );
not \U$57559 ( \57902 , \57901 );
xor \U$57560 ( \57903 , \57763 , \3406 );
xor \U$57561 ( \57904 , \57903 , \57771 );
nand \U$57562 ( \57905 , \57902 , \57904 );
xor \U$57563 ( \57906 , \57551 , \57558 );
xor \U$57564 ( \57907 , \57906 , \57566 );
xor \U$57565 ( \57908 , \57905 , \57907 );
xor \U$57566 ( \57909 , \57734 , \57741 );
xor \U$57567 ( \57910 , \57909 , \57749 );
not \U$57568 ( \57911 , \57910 );
not \U$57569 ( \57912 , \57687 );
not \U$57570 ( \57913 , \57698 );
or \U$57571 ( \57914 , \57912 , \57913 );
or \U$57572 ( \57915 , \57687 , \57698 );
nand \U$57573 ( \57916 , \57914 , \57915 );
not \U$57574 ( \57917 , \57916 );
not \U$57575 ( \57918 , \57680 );
and \U$57576 ( \57919 , \57917 , \57918 );
and \U$57577 ( \57920 , \57916 , \57680 );
nor \U$57578 ( \57921 , \57919 , \57920 );
not \U$57579 ( \57922 , \57921 );
and \U$57580 ( \57923 , \57911 , \57922 );
and \U$57581 ( \57924 , \57921 , \57910 );
xor \U$57582 ( \57925 , \57782 , \57789 );
xor \U$57583 ( \57926 , \57925 , \57797 );
nor \U$57584 ( \57927 , \57924 , \57926 );
nor \U$57585 ( \57928 , \57923 , \57927 );
and \U$57586 ( \57929 , \57908 , \57928 );
and \U$57587 ( \57930 , \57905 , \57907 );
or \U$57588 ( \57931 , \57929 , \57930 );
or \U$57589 ( \57932 , \57899 , \57931 );
not \U$57590 ( \57933 , \57931 );
not \U$57591 ( \57934 , \57899 );
or \U$57592 ( \57935 , \57933 , \57934 );
and \U$57593 ( \57936 , \13045 , RI9871758_126);
and \U$57594 ( \57937 , RI9871848_128, \13043 );
nor \U$57595 ( \57938 , \57936 , \57937 );
and \U$57596 ( \57939 , \57938 , \13047 );
not \U$57597 ( \57940 , \57938 );
and \U$57598 ( \57941 , \57940 , \12619 );
nor \U$57599 ( \57942 , \57939 , \57941 );
and \U$57600 ( \57943 , \11696 , RI98712a8_116);
and \U$57601 ( \57944 , RI98711b8_114, \11694 );
nor \U$57602 ( \57945 , \57943 , \57944 );
and \U$57603 ( \57946 , \57945 , \10965 );
not \U$57604 ( \57947 , \57945 );
and \U$57605 ( \57948 , \57947 , \11702 );
nor \U$57606 ( \57949 , \57946 , \57948 );
xor \U$57607 ( \57950 , \57942 , \57949 );
and \U$57608 ( \57951 , \12293 , RI9871398_118);
and \U$57609 ( \57952 , RI9871488_120, \12291 );
nor \U$57610 ( \57953 , \57951 , \57952 );
and \U$57611 ( \57954 , \57953 , \11687 );
not \U$57612 ( \57955 , \57953 );
and \U$57613 ( \57956 , \57955 , \11686 );
nor \U$57614 ( \57957 , \57954 , \57956 );
and \U$57615 ( \57958 , \57950 , \57957 );
and \U$57616 ( \57959 , \57942 , \57949 );
or \U$57617 ( \57960 , \57958 , \57959 );
and \U$57618 ( \57961 , \13882 , RI9871578_122);
and \U$57619 ( \57962 , RI9871668_124, \13880 );
nor \U$57620 ( \57963 , \57961 , \57962 );
and \U$57621 ( \57964 , \57963 , \13359 );
not \U$57622 ( \57965 , \57963 );
and \U$57623 ( \57966 , \57965 , \13358 );
nor \U$57624 ( \57967 , \57964 , \57966 );
and \U$57625 ( \57968 , \15780 , RI986e968_28);
and \U$57626 ( \57969 , RI986e878_26, RI9873648_192);
nor \U$57627 ( \57970 , \57968 , \57969 );
not \U$57628 ( \57971 , \57970 );
not \U$57629 ( \57972 , RI9873558_190);
and \U$57630 ( \57973 , \57971 , \57972 );
and \U$57631 ( \57974 , \57970 , RI9873558_190);
nor \U$57632 ( \57975 , \57973 , \57974 );
or \U$57633 ( \57976 , \57967 , \57975 );
not \U$57634 ( \57977 , \57975 );
not \U$57635 ( \57978 , \57967 );
or \U$57636 ( \57979 , \57977 , \57978 );
and \U$57637 ( \57980 , \14937 , RI986eb48_32);
and \U$57638 ( \57981 , RI986ea58_30, \14935 );
nor \U$57639 ( \57982 , \57980 , \57981 );
and \U$57640 ( \57983 , \57982 , \14539 );
not \U$57641 ( \57984 , \57982 );
and \U$57642 ( \57985 , \57984 , \14538 );
nor \U$57643 ( \57986 , \57983 , \57985 );
nand \U$57644 ( \57987 , \57979 , \57986 );
nand \U$57645 ( \57988 , \57976 , \57987 );
xor \U$57646 ( \57989 , \57960 , \57988 );
and \U$57647 ( \57990 , \9237 , RI9870df8_106);
and \U$57648 ( \57991 , RI9870a38_98, \9235 );
nor \U$57649 ( \57992 , \57990 , \57991 );
and \U$57650 ( \57993 , \57992 , \8836 );
not \U$57651 ( \57994 , \57992 );
and \U$57652 ( \57995 , \57994 , \9241 );
nor \U$57653 ( \57996 , \57993 , \57995 );
and \U$57654 ( \57997 , \9505 , RI9870ee8_108);
and \U$57655 ( \57998 , RI9870c18_102, \9503 );
nor \U$57656 ( \57999 , \57997 , \57998 );
and \U$57657 ( \58000 , \57999 , \9513 );
not \U$57658 ( \58001 , \57999 );
and \U$57659 ( \58002 , \58001 , \9510 );
nor \U$57660 ( \58003 , \58000 , \58002 );
or \U$57661 ( \58004 , \57996 , \58003 );
not \U$57662 ( \58005 , \58003 );
not \U$57663 ( \58006 , \57996 );
or \U$57664 ( \58007 , \58005 , \58006 );
and \U$57665 ( \58008 , \10424 , RI98710c8_112);
and \U$57666 ( \58009 , RI9870d08_104, \10422 );
nor \U$57667 ( \58010 , \58008 , \58009 );
and \U$57668 ( \58011 , \58010 , \9840 );
not \U$57669 ( \58012 , \58010 );
and \U$57670 ( \58013 , \58012 , \10428 );
nor \U$57671 ( \58014 , \58011 , \58013 );
nand \U$57672 ( \58015 , \58007 , \58014 );
nand \U$57673 ( \58016 , \58004 , \58015 );
and \U$57674 ( \58017 , \57989 , \58016 );
and \U$57675 ( \58018 , \57960 , \57988 );
nor \U$57676 ( \58019 , \58017 , \58018 );
nand \U$57677 ( \58020 , RI9870498_86, \3252 );
not \U$57678 ( \58021 , \58020 );
not \U$57679 ( \58022 , \3406 );
or \U$57680 ( \58023 , \58021 , \58022 );
or \U$57681 ( \58024 , \2935 , \58020 );
nand \U$57682 ( \58025 , \58023 , \58024 );
not \U$57683 ( \58026 , \3918 );
and \U$57684 ( \58027 , \3683 , RI9870588_88);
and \U$57685 ( \58028 , RI98703a8_84, \3681 );
nor \U$57686 ( \58029 , \58027 , \58028 );
not \U$57687 ( \58030 , \58029 );
or \U$57688 ( \58031 , \58026 , \58030 );
or \U$57689 ( \58032 , \58029 , \3918 );
nand \U$57690 ( \58033 , \58031 , \58032 );
xor \U$57691 ( \58034 , \58025 , \58033 );
xor \U$57692 ( \58035 , \57707 , \57714 );
xor \U$57693 ( \58036 , \58035 , \57723 );
and \U$57694 ( \58037 , \58034 , \58036 );
and \U$57695 ( \58038 , \58025 , \58033 );
nor \U$57696 ( \58039 , \58037 , \58038 );
or \U$57697 ( \58040 , \58019 , \58039 );
not \U$57698 ( \58041 , \58039 );
not \U$57699 ( \58042 , \58019 );
or \U$57700 ( \58043 , \58041 , \58042 );
and \U$57701 ( \58044 , \7079 , RI986ffe8_76);
and \U$57702 ( \58045 , RI986fef8_74, \7077 );
nor \U$57703 ( \58046 , \58044 , \58045 );
and \U$57704 ( \58047 , \58046 , \6709 );
not \U$57705 ( \58048 , \58046 );
and \U$57706 ( \58049 , \58048 , \6710 );
nor \U$57707 ( \58050 , \58047 , \58049 );
and \U$57708 ( \58051 , \8486 , RI9870fd8_110);
and \U$57709 ( \58052 , RI9870b28_100, \8484 );
nor \U$57710 ( \58053 , \58051 , \58052 );
and \U$57711 ( \58054 , \58053 , \8051 );
not \U$57712 ( \58055 , \58053 );
and \U$57713 ( \58056 , \58055 , \8050 );
nor \U$57714 ( \58057 , \58054 , \58056 );
or \U$57715 ( \58058 , \58050 , \58057 );
not \U$57716 ( \58059 , \58057 );
not \U$57717 ( \58060 , \58050 );
or \U$57718 ( \58061 , \58059 , \58060 );
and \U$57719 ( \58062 , \7729 , RI98700d8_78);
and \U$57720 ( \58063 , RI98701c8_80, \7727 );
nor \U$57721 ( \58064 , \58062 , \58063 );
and \U$57722 ( \58065 , \58064 , \7480 );
not \U$57723 ( \58066 , \58064 );
and \U$57724 ( \58067 , \58066 , \7733 );
nor \U$57725 ( \58068 , \58065 , \58067 );
nand \U$57726 ( \58069 , \58061 , \58068 );
nand \U$57727 ( \58070 , \58058 , \58069 );
and \U$57728 ( \58071 , \5318 , RI9870948_96);
and \U$57729 ( \58072 , RI9870858_94, \5316 );
nor \U$57730 ( \58073 , \58071 , \58072 );
and \U$57731 ( \58074 , \58073 , \5322 );
not \U$57732 ( \58075 , \58073 );
and \U$57733 ( \58076 , \58075 , \5052 );
nor \U$57734 ( \58077 , \58074 , \58076 );
and \U$57735 ( \58078 , \5881 , RI986fb38_66);
and \U$57736 ( \58079 , RI986fc28_68, \5879 );
nor \U$57737 ( \58080 , \58078 , \58079 );
and \U$57738 ( \58081 , \58080 , \5885 );
not \U$57739 ( \58082 , \58080 );
and \U$57740 ( \58083 , \58082 , \5594 );
nor \U$57741 ( \58084 , \58081 , \58083 );
or \U$57742 ( \58085 , \58077 , \58084 );
not \U$57743 ( \58086 , \58084 );
not \U$57744 ( \58087 , \58077 );
or \U$57745 ( \58088 , \58086 , \58087 );
and \U$57746 ( \58089 , \6453 , RI986fe08_72);
and \U$57747 ( \58090 , RI986fd18_70, \6451 );
nor \U$57748 ( \58091 , \58089 , \58090 );
and \U$57749 ( \58092 , \58091 , \6190 );
not \U$57750 ( \58093 , \58091 );
and \U$57751 ( \58094 , \58093 , \6705 );
nor \U$57752 ( \58095 , \58092 , \58094 );
nand \U$57753 ( \58096 , \58088 , \58095 );
nand \U$57754 ( \58097 , \58085 , \58096 );
xor \U$57755 ( \58098 , \58070 , \58097 );
and \U$57756 ( \58099 , \4203 , RI98703a8_84);
and \U$57757 ( \58100 , RI98702b8_82, \4201 );
nor \U$57758 ( \58101 , \58099 , \58100 );
and \U$57759 ( \58102 , \58101 , \4207 );
not \U$57760 ( \58103 , \58101 );
and \U$57761 ( \58104 , \58103 , \3923 );
nor \U$57762 ( \58105 , \58102 , \58104 );
not \U$57763 ( \58106 , \3918 );
and \U$57764 ( \58107 , \3683 , RI9870498_86);
and \U$57765 ( \58108 , RI9870588_88, \3681 );
nor \U$57766 ( \58109 , \58107 , \58108 );
not \U$57767 ( \58110 , \58109 );
or \U$57768 ( \58111 , \58106 , \58110 );
or \U$57769 ( \58112 , \58109 , \3918 );
nand \U$57770 ( \58113 , \58111 , \58112 );
xor \U$57771 ( \58114 , \58105 , \58113 );
not \U$57772 ( \58115 , \4521 );
and \U$57773 ( \58116 , \4710 , RI9870768_92);
and \U$57774 ( \58117 , RI9870678_90, \4708 );
nor \U$57775 ( \58118 , \58116 , \58117 );
not \U$57776 ( \58119 , \58118 );
or \U$57777 ( \58120 , \58115 , \58119 );
or \U$57778 ( \58121 , \58118 , \4519 );
nand \U$57779 ( \58122 , \58120 , \58121 );
and \U$57780 ( \58123 , \58114 , \58122 );
and \U$57781 ( \58124 , \58105 , \58113 );
or \U$57782 ( \58125 , \58123 , \58124 );
and \U$57783 ( \58126 , \58098 , \58125 );
and \U$57784 ( \58127 , \58070 , \58097 );
or \U$57785 ( \58128 , \58126 , \58127 );
nand \U$57786 ( \58129 , \58043 , \58128 );
nand \U$57787 ( \58130 , \58040 , \58129 );
nand \U$57788 ( \58131 , \57935 , \58130 );
nand \U$57789 ( \58132 , \57932 , \58131 );
xor \U$57790 ( \58133 , \57884 , \58132 );
xor \U$57791 ( \58134 , \57518 , \57598 );
xor \U$57792 ( \58135 , \58134 , \57611 );
xor \U$57793 ( \58136 , \57175 , \57194 );
xor \U$57794 ( \58137 , \58136 , \57220 );
xor \U$57795 ( \58138 , \57427 , \57432 );
xor \U$57796 ( \58139 , \58137 , \58138 );
xor \U$57797 ( \58140 , \57139 , \57141 );
xor \U$57798 ( \58141 , \58140 , \57144 );
xor \U$57799 ( \58142 , \57627 , \57634 );
xor \U$57800 ( \58143 , \58141 , \58142 );
xor \U$57801 ( \58144 , \58139 , \58143 );
xor \U$57802 ( \58145 , \58135 , \58144 );
and \U$57803 ( \58146 , \58133 , \58145 );
and \U$57804 ( \58147 , \57884 , \58132 );
or \U$57805 ( \58148 , \58146 , \58147 );
xor \U$57806 ( \58149 , \57004 , \57030 );
xor \U$57807 ( \58150 , \58149 , \57056 );
xor \U$57808 ( \58151 , \57644 , \57651 );
xor \U$57809 ( \58152 , \58150 , \58151 );
xor \U$57810 ( \58153 , \57223 , \57267 );
xor \U$57811 ( \58154 , \58153 , \57348 );
xor \U$57812 ( \58155 , \58152 , \58154 );
xor \U$57813 ( \58156 , \57437 , \57614 );
xor \U$57814 ( \58157 , \58156 , \57639 );
xor \U$57815 ( \58158 , \58155 , \58157 );
and \U$57816 ( \58159 , \58148 , \58158 );
xor \U$57817 ( \58160 , \57462 , \57489 );
xor \U$57818 ( \58161 , \58160 , \57515 );
and \U$57819 ( \58162 , \57873 , \58161 );
xor \U$57820 ( \58163 , \57462 , \57489 );
xor \U$57821 ( \58164 , \58163 , \57515 );
and \U$57822 ( \58165 , \57877 , \58164 );
and \U$57823 ( \58166 , \57873 , \57877 );
or \U$57824 ( \58167 , \58162 , \58165 , \58166 );
xor \U$57825 ( \58168 , \57755 , \57830 );
and \U$57826 ( \58169 , \58168 , \57849 );
and \U$57827 ( \58170 , \57755 , \57830 );
or \U$57828 ( \58171 , \58169 , \58170 );
xor \U$57829 ( \58172 , \58167 , \58171 );
xor \U$57830 ( \58173 , \57860 , \57862 );
and \U$57831 ( \58174 , \58173 , \57867 );
and \U$57832 ( \58175 , \57860 , \57862 );
or \U$57833 ( \58176 , \58174 , \58175 );
and \U$57834 ( \58177 , \58172 , \58176 );
and \U$57835 ( \58178 , \58167 , \58171 );
or \U$57836 ( \58179 , \58177 , \58178 );
xor \U$57837 ( \58180 , \57134 , \57136 );
xor \U$57838 ( \58181 , \58180 , \57147 );
xor \U$57839 ( \58182 , \58179 , \58181 );
xor \U$57840 ( \58183 , \57518 , \57598 );
xor \U$57841 ( \58184 , \58183 , \57611 );
and \U$57842 ( \58185 , \58139 , \58184 );
xor \U$57843 ( \58186 , \57518 , \57598 );
xor \U$57844 ( \58187 , \58186 , \57611 );
and \U$57845 ( \58188 , \58143 , \58187 );
and \U$57846 ( \58189 , \58139 , \58143 );
or \U$57847 ( \58190 , \58185 , \58188 , \58189 );
xor \U$57848 ( \58191 , \58182 , \58190 );
xor \U$57849 ( \58192 , \58152 , \58154 );
xor \U$57850 ( \58193 , \58192 , \58157 );
and \U$57851 ( \58194 , \58191 , \58193 );
and \U$57852 ( \58195 , \58148 , \58191 );
or \U$57853 ( \58196 , \58159 , \58194 , \58195 );
xor \U$57854 ( \58197 , \57673 , \58196 );
xor \U$57855 ( \58198 , \58179 , \58181 );
and \U$57856 ( \58199 , \58198 , \58190 );
and \U$57857 ( \58200 , \58179 , \58181 );
or \U$57858 ( \58201 , \58199 , \58200 );
xor \U$57859 ( \58202 , \57150 , \57351 );
xor \U$57860 ( \58203 , \58202 , \57366 );
xor \U$57861 ( \58204 , \58201 , \58203 );
xor \U$57862 ( \58205 , \58152 , \58154 );
and \U$57863 ( \58206 , \58205 , \58157 );
and \U$57864 ( \58207 , \58152 , \58154 );
or \U$57865 ( \58208 , \58206 , \58207 );
xor \U$57866 ( \58209 , \58204 , \58208 );
and \U$57867 ( \58210 , \58197 , \58209 );
and \U$57868 ( \58211 , \57673 , \58196 );
nor \U$57869 ( \58212 , \58210 , \58211 );
xnor \U$57870 ( \58213 , \57664 , \57422 );
not \U$57871 ( \58214 , \58213 );
not \U$57872 ( \58215 , \57419 );
and \U$57873 ( \58216 , \58214 , \58215 );
and \U$57874 ( \58217 , \58213 , \57419 );
nor \U$57875 ( \58218 , \58216 , \58217 );
not \U$57876 ( \58219 , \58218 );
xor \U$57877 ( \58220 , \58201 , \58203 );
and \U$57878 ( \58221 , \58220 , \58208 );
and \U$57879 ( \58222 , \58201 , \58203 );
or \U$57880 ( \58223 , \58221 , \58222 );
not \U$57881 ( \58224 , \58223 );
and \U$57882 ( \58225 , \58219 , \58224 );
and \U$57883 ( \58226 , \58218 , \58223 );
nor \U$57884 ( \58227 , \58225 , \58226 );
or \U$57885 ( \58228 , \58212 , \58227 );
xnor \U$57886 ( \58229 , \58227 , \58212 );
xor \U$57887 ( \58230 , \57673 , \58196 );
xor \U$57888 ( \58231 , \58230 , \58209 );
xor \U$57889 ( \58232 , \58152 , \58154 );
xor \U$57890 ( \58233 , \58232 , \58157 );
xor \U$57891 ( \58234 , \58148 , \58191 );
xor \U$57892 ( \58235 , \58233 , \58234 );
not \U$57893 ( \58236 , \58235 );
xor \U$57894 ( \58237 , \57884 , \58132 );
xor \U$57895 ( \58238 , \58237 , \58145 );
xor \U$57896 ( \58239 , \57905 , \57907 );
xor \U$57897 ( \58240 , \58239 , \57928 );
xnor \U$57898 ( \58241 , \57828 , \57800 );
not \U$57899 ( \58242 , \58241 );
not \U$57900 ( \58243 , \57774 );
and \U$57901 ( \58244 , \58242 , \58243 );
and \U$57902 ( \58245 , \58241 , \57774 );
nor \U$57903 ( \58246 , \58244 , \58245 );
or \U$57904 ( \58247 , \58240 , \58246 );
not \U$57905 ( \58248 , \58246 );
not \U$57906 ( \58249 , \58240 );
or \U$57907 ( \58250 , \58248 , \58249 );
xor \U$57908 ( \58251 , \57852 , \57854 );
xor \U$57909 ( \58252 , \58251 , \57857 );
xor \U$57910 ( \58253 , \57886 , \57893 );
xor \U$57911 ( \58254 , \58252 , \58253 );
nand \U$57912 ( \58255 , \58250 , \58254 );
nand \U$57913 ( \58256 , \58247 , \58255 );
xor \U$57914 ( \58257 , \57960 , \57988 );
xor \U$57915 ( \58258 , \58257 , \58016 );
xor \U$57916 ( \58259 , \58025 , \58033 );
xor \U$57917 ( \58260 , \58259 , \58036 );
xor \U$57918 ( \58261 , \58258 , \58260 );
xor \U$57919 ( \58262 , \58070 , \58097 );
xor \U$57920 ( \58263 , \58262 , \58125 );
and \U$57921 ( \58264 , \58261 , \58263 );
and \U$57922 ( \58265 , \58258 , \58260 );
or \U$57923 ( \58266 , \58264 , \58265 );
and \U$57924 ( \58267 , \4203 , RI9870588_88);
and \U$57925 ( \58268 , RI98703a8_84, \4201 );
nor \U$57926 ( \58269 , \58267 , \58268 );
and \U$57927 ( \58270 , \58269 , \3922 );
not \U$57928 ( \58271 , \58269 );
and \U$57929 ( \58272 , \58271 , \4207 );
nor \U$57930 ( \58273 , \58270 , \58272 );
not \U$57931 ( \58274 , \58273 );
and \U$57932 ( \58275 , \5318 , RI9870678_90);
and \U$57933 ( \58276 , RI9870948_96, \5316 );
nor \U$57934 ( \58277 , \58275 , \58276 );
and \U$57935 ( \58278 , \58277 , \5322 );
not \U$57936 ( \58279 , \58277 );
and \U$57937 ( \58280 , \58279 , \5052 );
nor \U$57938 ( \58281 , \58278 , \58280 );
not \U$57939 ( \58282 , \58281 );
and \U$57940 ( \58283 , \58274 , \58282 );
and \U$57941 ( \58284 , \58281 , \58273 );
and \U$57942 ( \58285 , \4710 , RI98702b8_82);
and \U$57943 ( \58286 , RI9870768_92, \4708 );
nor \U$57944 ( \58287 , \58285 , \58286 );
not \U$57945 ( \58288 , \58287 );
not \U$57946 ( \58289 , \4521 );
and \U$57947 ( \58290 , \58288 , \58289 );
and \U$57948 ( \58291 , \58287 , \4519 );
nor \U$57949 ( \58292 , \58290 , \58291 );
nor \U$57950 ( \58293 , \58284 , \58292 );
nor \U$57951 ( \58294 , \58283 , \58293 );
and \U$57952 ( \58295 , \7729 , RI986fef8_74);
and \U$57953 ( \58296 , RI98700d8_78, \7727 );
nor \U$57954 ( \58297 , \58295 , \58296 );
and \U$57955 ( \58298 , \58297 , \7733 );
not \U$57956 ( \58299 , \58297 );
and \U$57957 ( \58300 , \58299 , \7480 );
nor \U$57958 ( \58301 , \58298 , \58300 );
and \U$57959 ( \58302 , \8486 , RI98701c8_80);
and \U$57960 ( \58303 , RI9870fd8_110, \8484 );
nor \U$57961 ( \58304 , \58302 , \58303 );
and \U$57962 ( \58305 , \58304 , \8051 );
not \U$57963 ( \58306 , \58304 );
and \U$57964 ( \58307 , \58306 , \8050 );
nor \U$57965 ( \58308 , \58305 , \58307 );
or \U$57966 ( \58309 , \58301 , \58308 );
not \U$57967 ( \58310 , \58308 );
not \U$57968 ( \58311 , \58301 );
or \U$57969 ( \58312 , \58310 , \58311 );
and \U$57970 ( \58313 , \9237 , RI9870b28_100);
and \U$57971 ( \58314 , RI9870df8_106, \9235 );
nor \U$57972 ( \58315 , \58313 , \58314 );
and \U$57973 ( \58316 , \58315 , \9241 );
not \U$57974 ( \58317 , \58315 );
and \U$57975 ( \58318 , \58317 , \8836 );
nor \U$57976 ( \58319 , \58316 , \58318 );
nand \U$57977 ( \58320 , \58312 , \58319 );
nand \U$57978 ( \58321 , \58309 , \58320 );
not \U$57979 ( \58322 , \58321 );
or \U$57980 ( \58323 , \58294 , \58322 );
and \U$57981 ( \58324 , \58294 , \58322 );
and \U$57982 ( \58325 , \6453 , RI986fc28_68);
and \U$57983 ( \58326 , RI986fe08_72, \6451 );
nor \U$57984 ( \58327 , \58325 , \58326 );
and \U$57985 ( \58328 , \58327 , \6190 );
not \U$57986 ( \58329 , \58327 );
and \U$57987 ( \58330 , \58329 , \6180 );
nor \U$57988 ( \58331 , \58328 , \58330 );
and \U$57989 ( \58332 , \7079 , RI986fd18_70);
and \U$57990 ( \58333 , RI986ffe8_76, \7077 );
nor \U$57991 ( \58334 , \58332 , \58333 );
and \U$57992 ( \58335 , \58334 , \6710 );
not \U$57993 ( \58336 , \58334 );
and \U$57994 ( \58337 , \58336 , \6709 );
nor \U$57995 ( \58338 , \58335 , \58337 );
xor \U$57996 ( \58339 , \58331 , \58338 );
and \U$57997 ( \58340 , \5881 , RI9870858_94);
and \U$57998 ( \58341 , RI986fb38_66, \5879 );
nor \U$57999 ( \58342 , \58340 , \58341 );
and \U$58000 ( \58343 , \58342 , \5594 );
not \U$58001 ( \58344 , \58342 );
and \U$58002 ( \58345 , \58344 , \5885 );
nor \U$58003 ( \58346 , \58343 , \58345 );
and \U$58004 ( \58347 , \58339 , \58346 );
and \U$58005 ( \58348 , \58331 , \58338 );
nor \U$58006 ( \58349 , \58347 , \58348 );
nor \U$58007 ( \58350 , \58324 , \58349 );
not \U$58008 ( \58351 , \58350 );
nand \U$58009 ( \58352 , \58323 , \58351 );
and \U$58010 ( \58353 , \13045 , RI9871488_120);
and \U$58011 ( \58354 , RI9871758_126, \13043 );
nor \U$58012 ( \58355 , \58353 , \58354 );
and \U$58013 ( \58356 , \58355 , \12619 );
not \U$58014 ( \58357 , \58355 );
and \U$58015 ( \58358 , \58357 , \13047 );
nor \U$58016 ( \58359 , \58356 , \58358 );
and \U$58017 ( \58360 , \13882 , RI9871848_128);
and \U$58018 ( \58361 , RI9871578_122, \13880 );
nor \U$58019 ( \58362 , \58360 , \58361 );
and \U$58020 ( \58363 , \58362 , \13359 );
not \U$58021 ( \58364 , \58362 );
and \U$58022 ( \58365 , \58364 , \13358 );
nor \U$58023 ( \58366 , \58363 , \58365 );
xor \U$58024 ( \58367 , \58359 , \58366 );
and \U$58025 ( \58368 , \12293 , RI98711b8_114);
and \U$58026 ( \58369 , RI9871398_118, \12291 );
nor \U$58027 ( \58370 , \58368 , \58369 );
and \U$58028 ( \58371 , \58370 , \11686 );
not \U$58029 ( \58372 , \58370 );
and \U$58030 ( \58373 , \58372 , \11687 );
nor \U$58031 ( \58374 , \58371 , \58373 );
and \U$58032 ( \58375 , \58367 , \58374 );
and \U$58033 ( \58376 , \58359 , \58366 );
nor \U$58034 ( \58377 , \58375 , \58376 );
not \U$58035 ( \58378 , RI9873558_190);
and \U$58036 ( \58379 , \15780 , RI986ea58_30);
and \U$58037 ( \58380 , RI986e968_28, RI9873648_192);
nor \U$58038 ( \58381 , \58379 , \58380 );
not \U$58039 ( \58382 , \58381 );
or \U$58040 ( \58383 , \58378 , \58382 );
or \U$58041 ( \58384 , \58381 , RI9873558_190);
nand \U$58042 ( \58385 , \58383 , \58384 );
xor \U$58043 ( \58386 , \58385 , \3918 );
and \U$58044 ( \58387 , \14937 , RI9871668_124);
and \U$58045 ( \58388 , RI986eb48_32, \14935 );
nor \U$58046 ( \58389 , \58387 , \58388 );
and \U$58047 ( \58390 , \58389 , \14539 );
not \U$58048 ( \58391 , \58389 );
and \U$58049 ( \58392 , \58391 , \14538 );
nor \U$58050 ( \58393 , \58390 , \58392 );
and \U$58051 ( \58394 , \58386 , \58393 );
and \U$58052 ( \58395 , \58385 , \3918 );
or \U$58053 ( \58396 , \58394 , \58395 );
xor \U$58054 ( \58397 , \58377 , \58396 );
and \U$58055 ( \58398 , \9505 , RI9870a38_98);
and \U$58056 ( \58399 , RI9870ee8_108, \9503 );
nor \U$58057 ( \58400 , \58398 , \58399 );
and \U$58058 ( \58401 , \58400 , \9513 );
not \U$58059 ( \58402 , \58400 );
and \U$58060 ( \58403 , \58402 , \9510 );
nor \U$58061 ( \58404 , \58401 , \58403 );
and \U$58062 ( \58405 , \11696 , RI9870d08_104);
and \U$58063 ( \58406 , RI98712a8_116, \11694 );
nor \U$58064 ( \58407 , \58405 , \58406 );
and \U$58065 ( \58408 , \58407 , \11702 );
not \U$58066 ( \58409 , \58407 );
and \U$58067 ( \58410 , \58409 , \10965 );
nor \U$58068 ( \58411 , \58408 , \58410 );
or \U$58069 ( \58412 , \58404 , \58411 );
not \U$58070 ( \58413 , \58411 );
not \U$58071 ( \58414 , \58404 );
or \U$58072 ( \58415 , \58413 , \58414 );
and \U$58073 ( \58416 , \10424 , RI9870c18_102);
and \U$58074 ( \58417 , RI98710c8_112, \10422 );
nor \U$58075 ( \58418 , \58416 , \58417 );
and \U$58076 ( \58419 , \58418 , \9840 );
not \U$58077 ( \58420 , \58418 );
and \U$58078 ( \58421 , \58420 , \10428 );
nor \U$58079 ( \58422 , \58419 , \58421 );
nand \U$58080 ( \58423 , \58415 , \58422 );
nand \U$58081 ( \58424 , \58412 , \58423 );
and \U$58082 ( \58425 , \58397 , \58424 );
and \U$58083 ( \58426 , \58377 , \58396 );
or \U$58084 ( \58427 , \58425 , \58426 );
xor \U$58085 ( \58428 , \58352 , \58427 );
not \U$58086 ( \58429 , \58084 );
not \U$58087 ( \58430 , \58095 );
or \U$58088 ( \58431 , \58429 , \58430 );
or \U$58089 ( \58432 , \58084 , \58095 );
nand \U$58090 ( \58433 , \58431 , \58432 );
not \U$58091 ( \58434 , \58433 );
not \U$58092 ( \58435 , \58077 );
and \U$58093 ( \58436 , \58434 , \58435 );
and \U$58094 ( \58437 , \58433 , \58077 );
nor \U$58095 ( \58438 , \58436 , \58437 );
not \U$58096 ( \58439 , \58057 );
not \U$58097 ( \58440 , \58068 );
or \U$58098 ( \58441 , \58439 , \58440 );
or \U$58099 ( \58442 , \58057 , \58068 );
nand \U$58100 ( \58443 , \58441 , \58442 );
not \U$58101 ( \58444 , \58443 );
not \U$58102 ( \58445 , \58050 );
and \U$58103 ( \58446 , \58444 , \58445 );
and \U$58104 ( \58447 , \58443 , \58050 );
nor \U$58105 ( \58448 , \58446 , \58447 );
or \U$58106 ( \58449 , \58438 , \58448 );
not \U$58107 ( \58450 , \58448 );
not \U$58108 ( \58451 , \58438 );
or \U$58109 ( \58452 , \58450 , \58451 );
xor \U$58110 ( \58453 , \58105 , \58113 );
xor \U$58111 ( \58454 , \58453 , \58122 );
nand \U$58112 ( \58455 , \58452 , \58454 );
nand \U$58113 ( \58456 , \58449 , \58455 );
and \U$58114 ( \58457 , \58428 , \58456 );
and \U$58115 ( \58458 , \58352 , \58427 );
or \U$58116 ( \58459 , \58457 , \58458 );
xor \U$58117 ( \58460 , \58266 , \58459 );
not \U$58118 ( \58461 , \57975 );
not \U$58119 ( \58462 , \57986 );
or \U$58120 ( \58463 , \58461 , \58462 );
or \U$58121 ( \58464 , \57986 , \57975 );
nand \U$58122 ( \58465 , \58463 , \58464 );
not \U$58123 ( \58466 , \58465 );
not \U$58124 ( \58467 , \57967 );
and \U$58125 ( \58468 , \58466 , \58467 );
and \U$58126 ( \58469 , \58465 , \57967 );
nor \U$58127 ( \58470 , \58468 , \58469 );
not \U$58128 ( \58471 , \58003 );
not \U$58129 ( \58472 , \58014 );
or \U$58130 ( \58473 , \58471 , \58472 );
or \U$58131 ( \58474 , \58003 , \58014 );
nand \U$58132 ( \58475 , \58473 , \58474 );
not \U$58133 ( \58476 , \58475 );
not \U$58134 ( \58477 , \57996 );
and \U$58135 ( \58478 , \58476 , \58477 );
and \U$58136 ( \58479 , \58475 , \57996 );
nor \U$58137 ( \58480 , \58478 , \58479 );
or \U$58138 ( \58481 , \58470 , \58480 );
not \U$58139 ( \58482 , \58480 );
not \U$58140 ( \58483 , \58470 );
or \U$58141 ( \58484 , \58482 , \58483 );
xor \U$58142 ( \58485 , \57942 , \57949 );
xor \U$58143 ( \58486 , \58485 , \57957 );
nand \U$58144 ( \58487 , \58484 , \58486 );
nand \U$58145 ( \58488 , \58481 , \58487 );
not \U$58146 ( \58489 , \57901 );
not \U$58147 ( \58490 , \57904 );
or \U$58148 ( \58491 , \58489 , \58490 );
or \U$58149 ( \58492 , \57904 , \57901 );
nand \U$58150 ( \58493 , \58491 , \58492 );
xor \U$58151 ( \58494 , \58488 , \58493 );
not \U$58152 ( \58495 , \57910 );
xor \U$58153 ( \58496 , \57921 , \57926 );
not \U$58154 ( \58497 , \58496 );
or \U$58155 ( \58498 , \58495 , \58497 );
or \U$58156 ( \58499 , \58496 , \57910 );
nand \U$58157 ( \58500 , \58498 , \58499 );
and \U$58158 ( \58501 , \58494 , \58500 );
and \U$58159 ( \58502 , \58488 , \58493 );
or \U$58160 ( \58503 , \58501 , \58502 );
and \U$58161 ( \58504 , \58460 , \58503 );
and \U$58162 ( \58505 , \58266 , \58459 );
or \U$58163 ( \58506 , \58504 , \58505 );
xor \U$58164 ( \58507 , \58256 , \58506 );
xor \U$58165 ( \58508 , \57860 , \57862 );
xor \U$58166 ( \58509 , \58508 , \57867 );
xor \U$58167 ( \58510 , \57850 , \57879 );
xor \U$58168 ( \58511 , \58509 , \58510 );
and \U$58169 ( \58512 , \58507 , \58511 );
and \U$58170 ( \58513 , \58256 , \58506 );
or \U$58171 ( \58514 , \58512 , \58513 );
xor \U$58172 ( \58515 , \58238 , \58514 );
xor \U$58173 ( \58516 , \58167 , \58171 );
xor \U$58174 ( \58517 , \58516 , \58176 );
and \U$58175 ( \58518 , \58515 , \58517 );
and \U$58176 ( \58519 , \58238 , \58514 );
nor \U$58177 ( \58520 , \58518 , \58519 );
nor \U$58178 ( \58521 , \58236 , \58520 );
and \U$58179 ( \58522 , \58231 , \58521 );
xor \U$58180 ( \58523 , \58521 , \58231 );
xnor \U$58181 ( \58524 , \58246 , \58240 );
not \U$58182 ( \58525 , \58524 );
not \U$58183 ( \58526 , \58254 );
and \U$58184 ( \58527 , \58525 , \58526 );
and \U$58185 ( \58528 , \58524 , \58254 );
nor \U$58186 ( \58529 , \58527 , \58528 );
not \U$58187 ( \58530 , \58529 );
xor \U$58188 ( \58531 , \58266 , \58459 );
xor \U$58189 ( \58532 , \58531 , \58503 );
nand \U$58190 ( \58533 , \58530 , \58532 );
not \U$58191 ( \58534 , \58130 );
not \U$58192 ( \58535 , \57931 );
or \U$58193 ( \58536 , \58534 , \58535 );
or \U$58194 ( \58537 , \57931 , \58130 );
nand \U$58195 ( \58538 , \58536 , \58537 );
not \U$58196 ( \58539 , \58538 );
not \U$58197 ( \58540 , \57899 );
and \U$58198 ( \58541 , \58539 , \58540 );
and \U$58199 ( \58542 , \58538 , \57899 );
nor \U$58200 ( \58543 , \58541 , \58542 );
xor \U$58201 ( \58544 , \58533 , \58543 );
xor \U$58202 ( \58545 , \58352 , \58427 );
xor \U$58203 ( \58546 , \58545 , \58456 );
xor \U$58204 ( \58547 , \58258 , \58260 );
xor \U$58205 ( \58548 , \58547 , \58263 );
and \U$58206 ( \58549 , \58546 , \58548 );
xor \U$58207 ( \58550 , \58488 , \58493 );
xor \U$58208 ( \58551 , \58550 , \58500 );
xor \U$58209 ( \58552 , \58258 , \58260 );
xor \U$58210 ( \58553 , \58552 , \58263 );
and \U$58211 ( \58554 , \58551 , \58553 );
and \U$58212 ( \58555 , \58546 , \58551 );
or \U$58213 ( \58556 , \58549 , \58554 , \58555 );
not \U$58214 ( \58557 , \58556 );
not \U$58215 ( \58558 , \58557 );
not \U$58216 ( \58559 , \58019 );
not \U$58217 ( \58560 , \58128 );
or \U$58218 ( \58561 , \58559 , \58560 );
or \U$58219 ( \58562 , \58128 , \58019 );
nand \U$58220 ( \58563 , \58561 , \58562 );
not \U$58221 ( \58564 , \58563 );
not \U$58222 ( \58565 , \58039 );
and \U$58223 ( \58566 , \58564 , \58565 );
and \U$58224 ( \58567 , \58563 , \58039 );
nor \U$58225 ( \58568 , \58566 , \58567 );
not \U$58226 ( \58569 , \58568 );
and \U$58227 ( \58570 , \58558 , \58569 );
and \U$58228 ( \58571 , \58557 , \58568 );
and \U$58229 ( \58572 , \9505 , RI9870df8_106);
and \U$58230 ( \58573 , RI9870a38_98, \9503 );
nor \U$58231 ( \58574 , \58572 , \58573 );
and \U$58232 ( \58575 , \58574 , \9510 );
not \U$58233 ( \58576 , \58574 );
and \U$58234 ( \58577 , \58576 , \9513 );
nor \U$58235 ( \58578 , \58575 , \58577 );
and \U$58236 ( \58579 , \9237 , RI9870fd8_110);
and \U$58237 ( \58580 , RI9870b28_100, \9235 );
nor \U$58238 ( \58581 , \58579 , \58580 );
and \U$58239 ( \58582 , \58581 , \9241 );
not \U$58240 ( \58583 , \58581 );
and \U$58241 ( \58584 , \58583 , \8836 );
nor \U$58242 ( \58585 , \58582 , \58584 );
xor \U$58243 ( \58586 , \58578 , \58585 );
and \U$58244 ( \58587 , \10424 , RI9870ee8_108);
and \U$58245 ( \58588 , RI9870c18_102, \10422 );
nor \U$58246 ( \58589 , \58587 , \58588 );
and \U$58247 ( \58590 , \58589 , \9840 );
not \U$58248 ( \58591 , \58589 );
and \U$58249 ( \58592 , \58591 , \10428 );
nor \U$58250 ( \58593 , \58590 , \58592 );
and \U$58251 ( \58594 , \58586 , \58593 );
and \U$58252 ( \58595 , \58578 , \58585 );
or \U$58253 ( \58596 , \58594 , \58595 );
and \U$58254 ( \58597 , \13882 , RI9871758_126);
and \U$58255 ( \58598 , RI9871848_128, \13880 );
nor \U$58256 ( \58599 , \58597 , \58598 );
and \U$58257 ( \58600 , \58599 , \13358 );
not \U$58258 ( \58601 , \58599 );
and \U$58259 ( \58602 , \58601 , \13359 );
nor \U$58260 ( \58603 , \58600 , \58602 );
not \U$58261 ( \58604 , RI9873558_190);
and \U$58262 ( \58605 , \15780 , RI986eb48_32);
and \U$58263 ( \58606 , RI986ea58_30, RI9873648_192);
nor \U$58264 ( \58607 , \58605 , \58606 );
not \U$58265 ( \58608 , \58607 );
or \U$58266 ( \58609 , \58604 , \58608 );
or \U$58267 ( \58610 , \58607 , RI9873558_190);
nand \U$58268 ( \58611 , \58609 , \58610 );
xor \U$58269 ( \58612 , \58603 , \58611 );
and \U$58270 ( \58613 , \14937 , RI9871578_122);
and \U$58271 ( \58614 , RI9871668_124, \14935 );
nor \U$58272 ( \58615 , \58613 , \58614 );
and \U$58273 ( \58616 , \58615 , \14539 );
not \U$58274 ( \58617 , \58615 );
and \U$58275 ( \58618 , \58617 , \14538 );
nor \U$58276 ( \58619 , \58616 , \58618 );
and \U$58277 ( \58620 , \58612 , \58619 );
and \U$58278 ( \58621 , \58603 , \58611 );
or \U$58279 ( \58622 , \58620 , \58621 );
xor \U$58280 ( \58623 , \58596 , \58622 );
and \U$58281 ( \58624 , \11696 , RI98710c8_112);
and \U$58282 ( \58625 , RI9870d08_104, \11694 );
nor \U$58283 ( \58626 , \58624 , \58625 );
and \U$58284 ( \58627 , \58626 , \10965 );
not \U$58285 ( \58628 , \58626 );
and \U$58286 ( \58629 , \58628 , \11702 );
nor \U$58287 ( \58630 , \58627 , \58629 );
and \U$58288 ( \58631 , \12293 , RI98712a8_116);
and \U$58289 ( \58632 , RI98711b8_114, \12291 );
nor \U$58290 ( \58633 , \58631 , \58632 );
and \U$58291 ( \58634 , \58633 , \11687 );
not \U$58292 ( \58635 , \58633 );
and \U$58293 ( \58636 , \58635 , \11686 );
nor \U$58294 ( \58637 , \58634 , \58636 );
xor \U$58295 ( \58638 , \58630 , \58637 );
and \U$58296 ( \58639 , \13045 , RI9871398_118);
and \U$58297 ( \58640 , RI9871488_120, \13043 );
nor \U$58298 ( \58641 , \58639 , \58640 );
and \U$58299 ( \58642 , \58641 , \13047 );
not \U$58300 ( \58643 , \58641 );
and \U$58301 ( \58644 , \58643 , \12619 );
nor \U$58302 ( \58645 , \58642 , \58644 );
and \U$58303 ( \58646 , \58638 , \58645 );
and \U$58304 ( \58647 , \58630 , \58637 );
or \U$58305 ( \58648 , \58646 , \58647 );
and \U$58306 ( \58649 , \58623 , \58648 );
and \U$58307 ( \58650 , \58596 , \58622 );
or \U$58308 ( \58651 , \58649 , \58650 );
and \U$58309 ( \58652 , \8486 , RI98700d8_78);
and \U$58310 ( \58653 , RI98701c8_80, \8484 );
nor \U$58311 ( \58654 , \58652 , \58653 );
and \U$58312 ( \58655 , \58654 , \8050 );
not \U$58313 ( \58656 , \58654 );
and \U$58314 ( \58657 , \58656 , \8051 );
nor \U$58315 ( \58658 , \58655 , \58657 );
and \U$58316 ( \58659 , \7079 , RI986fe08_72);
and \U$58317 ( \58660 , RI986fd18_70, \7077 );
nor \U$58318 ( \58661 , \58659 , \58660 );
and \U$58319 ( \58662 , \58661 , \6710 );
not \U$58320 ( \58663 , \58661 );
and \U$58321 ( \58664 , \58663 , \6709 );
nor \U$58322 ( \58665 , \58662 , \58664 );
xor \U$58323 ( \58666 , \58658 , \58665 );
and \U$58324 ( \58667 , \7729 , RI986ffe8_76);
and \U$58325 ( \58668 , RI986fef8_74, \7727 );
nor \U$58326 ( \58669 , \58667 , \58668 );
and \U$58327 ( \58670 , \58669 , \7480 );
not \U$58328 ( \58671 , \58669 );
and \U$58329 ( \58672 , \58671 , \7733 );
nor \U$58330 ( \58673 , \58670 , \58672 );
and \U$58331 ( \58674 , \58666 , \58673 );
and \U$58332 ( \58675 , \58658 , \58665 );
or \U$58333 ( \58676 , \58674 , \58675 );
not \U$58334 ( \58677 , \4521 );
and \U$58335 ( \58678 , \4710 , RI98703a8_84);
and \U$58336 ( \58679 , RI98702b8_82, \4708 );
nor \U$58337 ( \58680 , \58678 , \58679 );
not \U$58338 ( \58681 , \58680 );
or \U$58339 ( \58682 , \58677 , \58681 );
or \U$58340 ( \58683 , \58680 , \4521 );
nand \U$58341 ( \58684 , \58682 , \58683 );
and \U$58342 ( \58685 , \4203 , RI9870498_86);
and \U$58343 ( \58686 , RI9870588_88, \4201 );
nor \U$58344 ( \58687 , \58685 , \58686 );
and \U$58345 ( \58688 , \58687 , \4207 );
not \U$58346 ( \58689 , \58687 );
and \U$58347 ( \58690 , \58689 , \3922 );
nor \U$58348 ( \58691 , \58688 , \58690 );
and \U$58349 ( \58692 , \58684 , \58691 );
xor \U$58350 ( \58693 , \58676 , \58692 );
and \U$58351 ( \58694 , \6453 , RI986fb38_66);
and \U$58352 ( \58695 , RI986fc28_68, \6451 );
nor \U$58353 ( \58696 , \58694 , \58695 );
and \U$58354 ( \58697 , \58696 , \6190 );
not \U$58355 ( \58698 , \58696 );
and \U$58356 ( \58699 , \58698 , \6705 );
nor \U$58357 ( \58700 , \58697 , \58699 );
and \U$58358 ( \58701 , \5318 , RI9870768_92);
and \U$58359 ( \58702 , RI9870678_90, \5316 );
nor \U$58360 ( \58703 , \58701 , \58702 );
and \U$58361 ( \58704 , \58703 , \5052 );
not \U$58362 ( \58705 , \58703 );
and \U$58363 ( \58706 , \58705 , \5322 );
nor \U$58364 ( \58707 , \58704 , \58706 );
xor \U$58365 ( \58708 , \58700 , \58707 );
and \U$58366 ( \58709 , \5881 , RI9870948_96);
and \U$58367 ( \58710 , RI9870858_94, \5879 );
nor \U$58368 ( \58711 , \58709 , \58710 );
and \U$58369 ( \58712 , \58711 , \5594 );
not \U$58370 ( \58713 , \58711 );
and \U$58371 ( \58714 , \58713 , \5885 );
nor \U$58372 ( \58715 , \58712 , \58714 );
and \U$58373 ( \58716 , \58708 , \58715 );
and \U$58374 ( \58717 , \58700 , \58707 );
or \U$58375 ( \58718 , \58716 , \58717 );
and \U$58376 ( \58719 , \58693 , \58718 );
and \U$58377 ( \58720 , \58676 , \58692 );
or \U$58378 ( \58721 , \58719 , \58720 );
xor \U$58379 ( \58722 , \58651 , \58721 );
xor \U$58380 ( \58723 , \58331 , \58338 );
xor \U$58381 ( \58724 , \58723 , \58346 );
nand \U$58382 ( \58725 , RI9870498_86, \3681 );
not \U$58383 ( \58726 , \58725 );
not \U$58384 ( \58727 , \3412 );
or \U$58385 ( \58728 , \58726 , \58727 );
or \U$58386 ( \58729 , \3412 , \58725 );
nand \U$58387 ( \58730 , \58728 , \58729 );
xor \U$58388 ( \58731 , \58724 , \58730 );
not \U$58389 ( \58732 , \58273 );
xor \U$58390 ( \58733 , \58292 , \58281 );
not \U$58391 ( \58734 , \58733 );
or \U$58392 ( \58735 , \58732 , \58734 );
or \U$58393 ( \58736 , \58733 , \58273 );
nand \U$58394 ( \58737 , \58735 , \58736 );
and \U$58395 ( \58738 , \58731 , \58737 );
and \U$58396 ( \58739 , \58724 , \58730 );
or \U$58397 ( \58740 , \58738 , \58739 );
and \U$58398 ( \58741 , \58722 , \58740 );
and \U$58399 ( \58742 , \58651 , \58721 );
nor \U$58400 ( \58743 , \58741 , \58742 );
not \U$58401 ( \58744 , \58743 );
not \U$58402 ( \58745 , \58321 );
not \U$58403 ( \58746 , \58349 );
or \U$58404 ( \58747 , \58745 , \58746 );
or \U$58405 ( \58748 , \58349 , \58321 );
nand \U$58406 ( \58749 , \58747 , \58748 );
not \U$58407 ( \58750 , \58749 );
not \U$58408 ( \58751 , \58294 );
and \U$58409 ( \58752 , \58750 , \58751 );
and \U$58410 ( \58753 , \58749 , \58294 );
nor \U$58411 ( \58754 , \58752 , \58753 );
not \U$58412 ( \58755 , \58754 );
xor \U$58413 ( \58756 , \58377 , \58396 );
xor \U$58414 ( \58757 , \58756 , \58424 );
nand \U$58415 ( \58758 , \58755 , \58757 );
not \U$58416 ( \58759 , \58758 );
and \U$58417 ( \58760 , \58744 , \58759 );
and \U$58418 ( \58761 , \58743 , \58758 );
not \U$58419 ( \58762 , \58486 );
not \U$58420 ( \58763 , \58470 );
or \U$58421 ( \58764 , \58762 , \58763 );
or \U$58422 ( \58765 , \58470 , \58486 );
nand \U$58423 ( \58766 , \58764 , \58765 );
not \U$58424 ( \58767 , \58766 );
not \U$58425 ( \58768 , \58480 );
and \U$58426 ( \58769 , \58767 , \58768 );
and \U$58427 ( \58770 , \58766 , \58480 );
nor \U$58428 ( \58771 , \58769 , \58770 );
not \U$58429 ( \58772 , \58771 );
not \U$58430 ( \58773 , \58308 );
not \U$58431 ( \58774 , \58319 );
or \U$58432 ( \58775 , \58773 , \58774 );
or \U$58433 ( \58776 , \58308 , \58319 );
nand \U$58434 ( \58777 , \58775 , \58776 );
not \U$58435 ( \58778 , \58777 );
not \U$58436 ( \58779 , \58301 );
and \U$58437 ( \58780 , \58778 , \58779 );
and \U$58438 ( \58781 , \58777 , \58301 );
nor \U$58439 ( \58782 , \58780 , \58781 );
not \U$58440 ( \58783 , \58782 );
not \U$58441 ( \58784 , \58411 );
not \U$58442 ( \58785 , \58422 );
or \U$58443 ( \58786 , \58784 , \58785 );
or \U$58444 ( \58787 , \58411 , \58422 );
nand \U$58445 ( \58788 , \58786 , \58787 );
not \U$58446 ( \58789 , \58788 );
not \U$58447 ( \58790 , \58404 );
and \U$58448 ( \58791 , \58789 , \58790 );
and \U$58449 ( \58792 , \58788 , \58404 );
nor \U$58450 ( \58793 , \58791 , \58792 );
not \U$58451 ( \58794 , \58793 );
and \U$58452 ( \58795 , \58783 , \58794 );
and \U$58453 ( \58796 , \58793 , \58782 );
xor \U$58454 ( \58797 , \58359 , \58366 );
xor \U$58455 ( \58798 , \58797 , \58374 );
nor \U$58456 ( \58799 , \58796 , \58798 );
nor \U$58457 ( \58800 , \58795 , \58799 );
not \U$58458 ( \58801 , \58800 );
and \U$58459 ( \58802 , \58772 , \58801 );
and \U$58460 ( \58803 , \58771 , \58800 );
not \U$58461 ( \58804 , \58438 );
not \U$58462 ( \58805 , \58454 );
or \U$58463 ( \58806 , \58804 , \58805 );
or \U$58464 ( \58807 , \58438 , \58454 );
nand \U$58465 ( \58808 , \58806 , \58807 );
not \U$58466 ( \58809 , \58808 );
not \U$58467 ( \58810 , \58448 );
and \U$58468 ( \58811 , \58809 , \58810 );
and \U$58469 ( \58812 , \58808 , \58448 );
nor \U$58470 ( \58813 , \58811 , \58812 );
nor \U$58471 ( \58814 , \58803 , \58813 );
nor \U$58472 ( \58815 , \58802 , \58814 );
nor \U$58473 ( \58816 , \58761 , \58815 );
nor \U$58474 ( \58817 , \58760 , \58816 );
nor \U$58475 ( \58818 , \58571 , \58817 );
nor \U$58476 ( \58819 , \58570 , \58818 );
and \U$58477 ( \58820 , \58544 , \58819 );
and \U$58478 ( \58821 , \58533 , \58543 );
or \U$58479 ( \58822 , \58820 , \58821 );
not \U$58480 ( \58823 , \58822 );
xor \U$58481 ( \58824 , \58238 , \58514 );
xor \U$58482 ( \58825 , \58824 , \58517 );
not \U$58483 ( \58826 , \58825 );
or \U$58484 ( \58827 , \58823 , \58826 );
or \U$58485 ( \58828 , \58825 , \58822 );
nand \U$58486 ( \58829 , \58827 , \58828 );
xor \U$58487 ( \58830 , \58256 , \58506 );
xor \U$58488 ( \58831 , \58830 , \58511 );
not \U$58489 ( \58832 , \58831 );
xor \U$58490 ( \58833 , \58533 , \58543 );
xor \U$58491 ( \58834 , \58833 , \58819 );
nor \U$58492 ( \58835 , \58832 , \58834 );
and \U$58493 ( \58836 , \58829 , \58835 );
xor \U$58494 ( \58837 , \58835 , \58829 );
not \U$58495 ( \58838 , \58834 );
not \U$58496 ( \58839 , \58831 );
and \U$58497 ( \58840 , \58838 , \58839 );
and \U$58498 ( \58841 , \58834 , \58831 );
nor \U$58499 ( \58842 , \58840 , \58841 );
not \U$58500 ( \58843 , \58532 );
not \U$58501 ( \58844 , \58529 );
or \U$58502 ( \58845 , \58843 , \58844 );
or \U$58503 ( \58846 , \58529 , \58532 );
nand \U$58504 ( \58847 , \58845 , \58846 );
xor \U$58505 ( \58848 , \58676 , \58692 );
xor \U$58506 ( \58849 , \58848 , \58718 );
xor \U$58507 ( \58850 , \58596 , \58622 );
xor \U$58508 ( \58851 , \58850 , \58648 );
and \U$58509 ( \58852 , \58849 , \58851 );
xor \U$58510 ( \58853 , \58724 , \58730 );
xor \U$58511 ( \58854 , \58853 , \58737 );
xor \U$58512 ( \58855 , \58596 , \58622 );
xor \U$58513 ( \58856 , \58855 , \58648 );
and \U$58514 ( \58857 , \58854 , \58856 );
and \U$58515 ( \58858 , \58849 , \58854 );
or \U$58516 ( \58859 , \58852 , \58857 , \58858 );
and \U$58517 ( \58860 , \7079 , RI986fc28_68);
and \U$58518 ( \58861 , RI986fe08_72, \7077 );
nor \U$58519 ( \58862 , \58860 , \58861 );
and \U$58520 ( \58863 , \58862 , \6710 );
not \U$58521 ( \58864 , \58862 );
and \U$58522 ( \58865 , \58864 , \6709 );
nor \U$58523 ( \58866 , \58863 , \58865 );
and \U$58524 ( \58867 , \5881 , RI9870678_90);
and \U$58525 ( \58868 , RI9870948_96, \5879 );
nor \U$58526 ( \58869 , \58867 , \58868 );
and \U$58527 ( \58870 , \58869 , \5594 );
not \U$58528 ( \58871 , \58869 );
and \U$58529 ( \58872 , \58871 , \5885 );
nor \U$58530 ( \58873 , \58870 , \58872 );
xor \U$58531 ( \58874 , \58866 , \58873 );
and \U$58532 ( \58875 , \6453 , RI9870858_94);
and \U$58533 ( \58876 , RI986fb38_66, \6451 );
nor \U$58534 ( \58877 , \58875 , \58876 );
and \U$58535 ( \58878 , \58877 , \6190 );
not \U$58536 ( \58879 , \58877 );
and \U$58537 ( \58880 , \58879 , \6705 );
nor \U$58538 ( \58881 , \58878 , \58880 );
and \U$58539 ( \58882 , \58874 , \58881 );
and \U$58540 ( \58883 , \58866 , \58873 );
or \U$58541 ( \58884 , \58882 , \58883 );
and \U$58542 ( \58885 , \5318 , RI98702b8_82);
and \U$58543 ( \58886 , RI9870768_92, \5316 );
nor \U$58544 ( \58887 , \58885 , \58886 );
and \U$58545 ( \58888 , \58887 , \5052 );
not \U$58546 ( \58889 , \58887 );
and \U$58547 ( \58890 , \58889 , \5322 );
nor \U$58548 ( \58891 , \58888 , \58890 );
nand \U$58549 ( \58892 , RI9870498_86, \4201 );
and \U$58550 ( \58893 , \58892 , \4207 );
not \U$58551 ( \58894 , \58892 );
and \U$58552 ( \58895 , \58894 , \3923 );
nor \U$58553 ( \58896 , \58893 , \58895 );
xor \U$58554 ( \58897 , \58891 , \58896 );
not \U$58555 ( \58898 , \4521 );
and \U$58556 ( \58899 , \4710 , RI9870588_88);
and \U$58557 ( \58900 , RI98703a8_84, \4708 );
nor \U$58558 ( \58901 , \58899 , \58900 );
not \U$58559 ( \58902 , \58901 );
or \U$58560 ( \58903 , \58898 , \58902 );
or \U$58561 ( \58904 , \58901 , \4521 );
nand \U$58562 ( \58905 , \58903 , \58904 );
and \U$58563 ( \58906 , \58897 , \58905 );
and \U$58564 ( \58907 , \58891 , \58896 );
or \U$58565 ( \58908 , \58906 , \58907 );
xor \U$58566 ( \58909 , \58884 , \58908 );
and \U$58567 ( \58910 , \9237 , RI98701c8_80);
and \U$58568 ( \58911 , RI9870fd8_110, \9235 );
nor \U$58569 ( \58912 , \58910 , \58911 );
and \U$58570 ( \58913 , \58912 , \9241 );
not \U$58571 ( \58914 , \58912 );
and \U$58572 ( \58915 , \58914 , \8836 );
nor \U$58573 ( \58916 , \58913 , \58915 );
and \U$58574 ( \58917 , \7729 , RI986fd18_70);
and \U$58575 ( \58918 , RI986ffe8_76, \7727 );
nor \U$58576 ( \58919 , \58917 , \58918 );
and \U$58577 ( \58920 , \58919 , \7480 );
not \U$58578 ( \58921 , \58919 );
and \U$58579 ( \58922 , \58921 , \7733 );
nor \U$58580 ( \58923 , \58920 , \58922 );
xor \U$58581 ( \58924 , \58916 , \58923 );
and \U$58582 ( \58925 , \8486 , RI986fef8_74);
and \U$58583 ( \58926 , RI98700d8_78, \8484 );
nor \U$58584 ( \58927 , \58925 , \58926 );
and \U$58585 ( \58928 , \58927 , \8050 );
not \U$58586 ( \58929 , \58927 );
and \U$58587 ( \58930 , \58929 , \8051 );
nor \U$58588 ( \58931 , \58928 , \58930 );
and \U$58589 ( \58932 , \58924 , \58931 );
and \U$58590 ( \58933 , \58916 , \58923 );
or \U$58591 ( \58934 , \58932 , \58933 );
and \U$58592 ( \58935 , \58909 , \58934 );
and \U$58593 ( \58936 , \58884 , \58908 );
or \U$58594 ( \58937 , \58935 , \58936 );
and \U$58595 ( \58938 , \11696 , RI9870c18_102);
and \U$58596 ( \58939 , RI98710c8_112, \11694 );
nor \U$58597 ( \58940 , \58938 , \58939 );
and \U$58598 ( \58941 , \58940 , \10965 );
not \U$58599 ( \58942 , \58940 );
and \U$58600 ( \58943 , \58942 , \11702 );
nor \U$58601 ( \58944 , \58941 , \58943 );
and \U$58602 ( \58945 , \9505 , RI9870b28_100);
and \U$58603 ( \58946 , RI9870df8_106, \9503 );
nor \U$58604 ( \58947 , \58945 , \58946 );
and \U$58605 ( \58948 , \58947 , \9510 );
not \U$58606 ( \58949 , \58947 );
and \U$58607 ( \58950 , \58949 , \9513 );
nor \U$58608 ( \58951 , \58948 , \58950 );
xor \U$58609 ( \58952 , \58944 , \58951 );
and \U$58610 ( \58953 , \10424 , RI9870a38_98);
and \U$58611 ( \58954 , RI9870ee8_108, \10422 );
nor \U$58612 ( \58955 , \58953 , \58954 );
and \U$58613 ( \58956 , \58955 , \9840 );
not \U$58614 ( \58957 , \58955 );
and \U$58615 ( \58958 , \58957 , \10428 );
nor \U$58616 ( \58959 , \58956 , \58958 );
and \U$58617 ( \58960 , \58952 , \58959 );
and \U$58618 ( \58961 , \58944 , \58951 );
or \U$58619 ( \58962 , \58960 , \58961 );
not \U$58620 ( \58963 , RI9873558_190);
and \U$58621 ( \58964 , \15780 , RI9871668_124);
and \U$58622 ( \58965 , RI986eb48_32, RI9873648_192);
nor \U$58623 ( \58966 , \58964 , \58965 );
not \U$58624 ( \58967 , \58966 );
or \U$58625 ( \58968 , \58963 , \58967 );
or \U$58626 ( \58969 , \58966 , RI9873558_190);
nand \U$58627 ( \58970 , \58968 , \58969 );
xor \U$58628 ( \58971 , \58970 , \3922 );
and \U$58629 ( \58972 , \14937 , RI9871848_128);
and \U$58630 ( \58973 , RI9871578_122, \14935 );
nor \U$58631 ( \58974 , \58972 , \58973 );
and \U$58632 ( \58975 , \58974 , \14539 );
not \U$58633 ( \58976 , \58974 );
and \U$58634 ( \58977 , \58976 , \14538 );
nor \U$58635 ( \58978 , \58975 , \58977 );
and \U$58636 ( \58979 , \58971 , \58978 );
and \U$58637 ( \58980 , \58970 , \3922 );
or \U$58638 ( \58981 , \58979 , \58980 );
xor \U$58639 ( \58982 , \58962 , \58981 );
and \U$58640 ( \58983 , \13882 , RI9871488_120);
and \U$58641 ( \58984 , RI9871758_126, \13880 );
nor \U$58642 ( \58985 , \58983 , \58984 );
and \U$58643 ( \58986 , \58985 , \13358 );
not \U$58644 ( \58987 , \58985 );
and \U$58645 ( \58988 , \58987 , \13359 );
nor \U$58646 ( \58989 , \58986 , \58988 );
and \U$58647 ( \58990 , \12293 , RI9870d08_104);
and \U$58648 ( \58991 , RI98712a8_116, \12291 );
nor \U$58649 ( \58992 , \58990 , \58991 );
and \U$58650 ( \58993 , \58992 , \11687 );
not \U$58651 ( \58994 , \58992 );
and \U$58652 ( \58995 , \58994 , \11686 );
nor \U$58653 ( \58996 , \58993 , \58995 );
xor \U$58654 ( \58997 , \58989 , \58996 );
and \U$58655 ( \58998 , \13045 , RI98711b8_114);
and \U$58656 ( \58999 , RI9871398_118, \13043 );
nor \U$58657 ( \59000 , \58998 , \58999 );
and \U$58658 ( \59001 , \59000 , \13047 );
not \U$58659 ( \59002 , \59000 );
and \U$58660 ( \59003 , \59002 , \12619 );
nor \U$58661 ( \59004 , \59001 , \59003 );
and \U$58662 ( \59005 , \58997 , \59004 );
and \U$58663 ( \59006 , \58989 , \58996 );
or \U$58664 ( \59007 , \59005 , \59006 );
and \U$58665 ( \59008 , \58982 , \59007 );
and \U$58666 ( \59009 , \58962 , \58981 );
or \U$58667 ( \59010 , \59008 , \59009 );
xor \U$58668 ( \59011 , \58937 , \59010 );
xor \U$58669 ( \59012 , \58658 , \58665 );
xor \U$58670 ( \59013 , \59012 , \58673 );
xor \U$58671 ( \59014 , \58684 , \58691 );
xor \U$58672 ( \59015 , \59013 , \59014 );
xor \U$58673 ( \59016 , \58700 , \58707 );
xor \U$58674 ( \59017 , \59016 , \58715 );
and \U$58675 ( \59018 , \59015 , \59017 );
and \U$58676 ( \59019 , \59013 , \59014 );
or \U$58677 ( \59020 , \59018 , \59019 );
and \U$58678 ( \59021 , \59011 , \59020 );
and \U$58679 ( \59022 , \58937 , \59010 );
or \U$58680 ( \59023 , \59021 , \59022 );
xor \U$58681 ( \59024 , \58859 , \59023 );
xor \U$58682 ( \59025 , \58603 , \58611 );
xor \U$58683 ( \59026 , \59025 , \58619 );
xor \U$58684 ( \59027 , \58630 , \58637 );
xor \U$58685 ( \59028 , \59027 , \58645 );
and \U$58686 ( \59029 , \59026 , \59028 );
xor \U$58687 ( \59030 , \58578 , \58585 );
xor \U$58688 ( \59031 , \59030 , \58593 );
xor \U$58689 ( \59032 , \58630 , \58637 );
xor \U$58690 ( \59033 , \59032 , \58645 );
and \U$58691 ( \59034 , \59031 , \59033 );
and \U$58692 ( \59035 , \59026 , \59031 );
or \U$58693 ( \59036 , \59029 , \59034 , \59035 );
xor \U$58694 ( \59037 , \58385 , \3918 );
xor \U$58695 ( \59038 , \59037 , \58393 );
xor \U$58696 ( \59039 , \59036 , \59038 );
not \U$58697 ( \59040 , \58793 );
xor \U$58698 ( \59041 , \58782 , \58798 );
not \U$58699 ( \59042 , \59041 );
or \U$58700 ( \59043 , \59040 , \59042 );
or \U$58701 ( \59044 , \59041 , \58793 );
nand \U$58702 ( \59045 , \59043 , \59044 );
and \U$58703 ( \59046 , \59039 , \59045 );
and \U$58704 ( \59047 , \59036 , \59038 );
or \U$58705 ( \59048 , \59046 , \59047 );
and \U$58706 ( \59049 , \59024 , \59048 );
and \U$58707 ( \59050 , \58859 , \59023 );
or \U$58708 ( \59051 , \59049 , \59050 );
xor \U$58709 ( \59052 , \58651 , \58721 );
xor \U$58710 ( \59053 , \59052 , \58740 );
not \U$58711 ( \59054 , \58757 );
not \U$58712 ( \59055 , \58754 );
or \U$58713 ( \59056 , \59054 , \59055 );
or \U$58714 ( \59057 , \58754 , \58757 );
nand \U$58715 ( \59058 , \59056 , \59057 );
xor \U$58716 ( \59059 , \59053 , \59058 );
not \U$58717 ( \59060 , \58771 );
xor \U$58718 ( \59061 , \58800 , \58813 );
not \U$58719 ( \59062 , \59061 );
or \U$58720 ( \59063 , \59060 , \59062 );
or \U$58721 ( \59064 , \59061 , \58771 );
nand \U$58722 ( \59065 , \59063 , \59064 );
and \U$58723 ( \59066 , \59059 , \59065 );
and \U$58724 ( \59067 , \59053 , \59058 );
or \U$58725 ( \59068 , \59066 , \59067 );
xor \U$58726 ( \59069 , \59051 , \59068 );
xor \U$58727 ( \59070 , \58258 , \58260 );
xor \U$58728 ( \59071 , \59070 , \58263 );
xor \U$58729 ( \59072 , \58546 , \58551 );
xor \U$58730 ( \59073 , \59071 , \59072 );
and \U$58731 ( \59074 , \59069 , \59073 );
and \U$58732 ( \59075 , \59051 , \59068 );
or \U$58733 ( \59076 , \59074 , \59075 );
xor \U$58734 ( \59077 , \58847 , \59076 );
not \U$58735 ( \59078 , \58568 );
xor \U$58736 ( \59079 , \58817 , \58557 );
not \U$58737 ( \59080 , \59079 );
or \U$58738 ( \59081 , \59078 , \59080 );
or \U$58739 ( \59082 , \59079 , \58568 );
nand \U$58740 ( \59083 , \59081 , \59082 );
and \U$58741 ( \59084 , \59077 , \59083 );
and \U$58742 ( \59085 , \58847 , \59076 );
nor \U$58743 ( \59086 , \59084 , \59085 );
or \U$58744 ( \59087 , \58842 , \59086 );
xnor \U$58745 ( \59088 , \59086 , \58842 );
xor \U$58746 ( \59089 , \58847 , \59076 );
xor \U$58747 ( \59090 , \59089 , \59083 );
not \U$58748 ( \59091 , \58758 );
xor \U$58749 ( \59092 , \58743 , \58815 );
not \U$58750 ( \59093 , \59092 );
or \U$58751 ( \59094 , \59091 , \59093 );
or \U$58752 ( \59095 , \59092 , \58758 );
nand \U$58753 ( \59096 , \59094 , \59095 );
not \U$58754 ( \59097 , \59096 );
xor \U$58755 ( \59098 , \59051 , \59068 );
xor \U$58756 ( \59099 , \59098 , \59073 );
not \U$58757 ( \59100 , \59099 );
or \U$58758 ( \59101 , \59097 , \59100 );
or \U$58759 ( \59102 , \59099 , \59096 );
xor \U$58760 ( \59103 , \58884 , \58908 );
xor \U$58761 ( \59104 , \59103 , \58934 );
xor \U$58762 ( \59105 , \59013 , \59014 );
xor \U$58763 ( \59106 , \59105 , \59017 );
and \U$58764 ( \59107 , \59104 , \59106 );
xor \U$58765 ( \59108 , \58630 , \58637 );
xor \U$58766 ( \59109 , \59108 , \58645 );
xor \U$58767 ( \59110 , \59026 , \59031 );
xor \U$58768 ( \59111 , \59109 , \59110 );
xor \U$58769 ( \59112 , \59013 , \59014 );
xor \U$58770 ( \59113 , \59112 , \59017 );
and \U$58771 ( \59114 , \59111 , \59113 );
and \U$58772 ( \59115 , \59104 , \59111 );
or \U$58773 ( \59116 , \59107 , \59114 , \59115 );
and \U$58774 ( \59117 , \7079 , RI986fb38_66);
and \U$58775 ( \59118 , RI986fc28_68, \7077 );
nor \U$58776 ( \59119 , \59117 , \59118 );
and \U$58777 ( \59120 , \59119 , \6710 );
not \U$58778 ( \59121 , \59119 );
and \U$58779 ( \59122 , \59121 , \6709 );
nor \U$58780 ( \59123 , \59120 , \59122 );
and \U$58781 ( \59124 , \7729 , RI986fe08_72);
and \U$58782 ( \59125 , RI986fd18_70, \7727 );
nor \U$58783 ( \59126 , \59124 , \59125 );
and \U$58784 ( \59127 , \59126 , \7480 );
not \U$58785 ( \59128 , \59126 );
and \U$58786 ( \59129 , \59128 , \7733 );
nor \U$58787 ( \59130 , \59127 , \59129 );
xor \U$58788 ( \59131 , \59123 , \59130 );
and \U$58789 ( \59132 , \8486 , RI986ffe8_76);
and \U$58790 ( \59133 , RI986fef8_74, \8484 );
nor \U$58791 ( \59134 , \59132 , \59133 );
and \U$58792 ( \59135 , \59134 , \8050 );
not \U$58793 ( \59136 , \59134 );
and \U$58794 ( \59137 , \59136 , \8051 );
nor \U$58795 ( \59138 , \59135 , \59137 );
and \U$58796 ( \59139 , \59131 , \59138 );
and \U$58797 ( \59140 , \59123 , \59130 );
or \U$58798 ( \59141 , \59139 , \59140 );
and \U$58799 ( \59142 , \5881 , RI9870768_92);
and \U$58800 ( \59143 , RI9870678_90, \5879 );
nor \U$58801 ( \59144 , \59142 , \59143 );
and \U$58802 ( \59145 , \59144 , \5594 );
not \U$58803 ( \59146 , \59144 );
and \U$58804 ( \59147 , \59146 , \5885 );
nor \U$58805 ( \59148 , \59145 , \59147 );
and \U$58806 ( \59149 , \5318 , RI98703a8_84);
and \U$58807 ( \59150 , RI98702b8_82, \5316 );
nor \U$58808 ( \59151 , \59149 , \59150 );
and \U$58809 ( \59152 , \59151 , \5052 );
not \U$58810 ( \59153 , \59151 );
and \U$58811 ( \59154 , \59153 , \5322 );
nor \U$58812 ( \59155 , \59152 , \59154 );
xor \U$58813 ( \59156 , \59148 , \59155 );
and \U$58814 ( \59157 , \6453 , RI9870948_96);
and \U$58815 ( \59158 , RI9870858_94, \6451 );
nor \U$58816 ( \59159 , \59157 , \59158 );
and \U$58817 ( \59160 , \59159 , \6190 );
not \U$58818 ( \59161 , \59159 );
and \U$58819 ( \59162 , \59161 , \6180 );
nor \U$58820 ( \59163 , \59160 , \59162 );
and \U$58821 ( \59164 , \59156 , \59163 );
and \U$58822 ( \59165 , \59148 , \59155 );
or \U$58823 ( \59166 , \59164 , \59165 );
xor \U$58824 ( \59167 , \59141 , \59166 );
xor \U$58825 ( \59168 , \58891 , \58896 );
xor \U$58826 ( \59169 , \59168 , \58905 );
and \U$58827 ( \59170 , \59167 , \59169 );
and \U$58828 ( \59171 , \59141 , \59166 );
or \U$58829 ( \59172 , \59170 , \59171 );
and \U$58830 ( \59173 , \10424 , RI9870df8_106);
and \U$58831 ( \59174 , RI9870a38_98, \10422 );
nor \U$58832 ( \59175 , \59173 , \59174 );
and \U$58833 ( \59176 , \59175 , \9840 );
not \U$58834 ( \59177 , \59175 );
and \U$58835 ( \59178 , \59177 , \10428 );
nor \U$58836 ( \59179 , \59176 , \59178 );
and \U$58837 ( \59180 , \9237 , RI98700d8_78);
and \U$58838 ( \59181 , RI98701c8_80, \9235 );
nor \U$58839 ( \59182 , \59180 , \59181 );
and \U$58840 ( \59183 , \59182 , \9241 );
not \U$58841 ( \59184 , \59182 );
and \U$58842 ( \59185 , \59184 , \8836 );
nor \U$58843 ( \59186 , \59183 , \59185 );
xor \U$58844 ( \59187 , \59179 , \59186 );
and \U$58845 ( \59188 , \9505 , RI9870fd8_110);
and \U$58846 ( \59189 , RI9870b28_100, \9503 );
nor \U$58847 ( \59190 , \59188 , \59189 );
and \U$58848 ( \59191 , \59190 , \9510 );
not \U$58849 ( \59192 , \59190 );
and \U$58850 ( \59193 , \59192 , \9513 );
nor \U$58851 ( \59194 , \59191 , \59193 );
and \U$58852 ( \59195 , \59187 , \59194 );
and \U$58853 ( \59196 , \59179 , \59186 );
or \U$58854 ( \59197 , \59195 , \59196 );
and \U$58855 ( \59198 , \13882 , RI9871398_118);
and \U$58856 ( \59199 , RI9871488_120, \13880 );
nor \U$58857 ( \59200 , \59198 , \59199 );
and \U$58858 ( \59201 , \59200 , \13358 );
not \U$58859 ( \59202 , \59200 );
and \U$58860 ( \59203 , \59202 , \13359 );
nor \U$58861 ( \59204 , \59201 , \59203 );
not \U$58862 ( \59205 , RI9873558_190);
and \U$58863 ( \59206 , \15780 , RI9871578_122);
and \U$58864 ( \59207 , RI9871668_124, RI9873648_192);
nor \U$58865 ( \59208 , \59206 , \59207 );
not \U$58866 ( \59209 , \59208 );
or \U$58867 ( \59210 , \59205 , \59209 );
or \U$58868 ( \59211 , \59208 , RI9873558_190);
nand \U$58869 ( \59212 , \59210 , \59211 );
xor \U$58870 ( \59213 , \59204 , \59212 );
and \U$58871 ( \59214 , \14937 , RI9871758_126);
and \U$58872 ( \59215 , RI9871848_128, \14935 );
nor \U$58873 ( \59216 , \59214 , \59215 );
and \U$58874 ( \59217 , \59216 , \14539 );
not \U$58875 ( \59218 , \59216 );
and \U$58876 ( \59219 , \59218 , \14538 );
nor \U$58877 ( \59220 , \59217 , \59219 );
and \U$58878 ( \59221 , \59213 , \59220 );
and \U$58879 ( \59222 , \59204 , \59212 );
or \U$58880 ( \59223 , \59221 , \59222 );
xor \U$58881 ( \59224 , \59197 , \59223 );
and \U$58882 ( \59225 , \13045 , RI98712a8_116);
and \U$58883 ( \59226 , RI98711b8_114, \13043 );
nor \U$58884 ( \59227 , \59225 , \59226 );
and \U$58885 ( \59228 , \59227 , \13047 );
not \U$58886 ( \59229 , \59227 );
and \U$58887 ( \59230 , \59229 , \12619 );
nor \U$58888 ( \59231 , \59228 , \59230 );
and \U$58889 ( \59232 , \11696 , RI9870ee8_108);
and \U$58890 ( \59233 , RI9870c18_102, \11694 );
nor \U$58891 ( \59234 , \59232 , \59233 );
and \U$58892 ( \59235 , \59234 , \10965 );
not \U$58893 ( \59236 , \59234 );
and \U$58894 ( \59237 , \59236 , \11702 );
nor \U$58895 ( \59238 , \59235 , \59237 );
xor \U$58896 ( \59239 , \59231 , \59238 );
and \U$58897 ( \59240 , \12293 , RI98710c8_112);
and \U$58898 ( \59241 , RI9870d08_104, \12291 );
nor \U$58899 ( \59242 , \59240 , \59241 );
and \U$58900 ( \59243 , \59242 , \11687 );
not \U$58901 ( \59244 , \59242 );
and \U$58902 ( \59245 , \59244 , \11686 );
nor \U$58903 ( \59246 , \59243 , \59245 );
and \U$58904 ( \59247 , \59239 , \59246 );
and \U$58905 ( \59248 , \59231 , \59238 );
or \U$58906 ( \59249 , \59247 , \59248 );
and \U$58907 ( \59250 , \59224 , \59249 );
and \U$58908 ( \59251 , \59197 , \59223 );
or \U$58909 ( \59252 , \59250 , \59251 );
xor \U$58910 ( \59253 , \59172 , \59252 );
xor \U$58911 ( \59254 , \58866 , \58873 );
xor \U$58912 ( \59255 , \59254 , \58881 );
xor \U$58913 ( \59256 , \58944 , \58951 );
xor \U$58914 ( \59257 , \59256 , \58959 );
and \U$58915 ( \59258 , \59255 , \59257 );
xor \U$58916 ( \59259 , \58916 , \58923 );
xor \U$58917 ( \59260 , \59259 , \58931 );
xor \U$58918 ( \59261 , \58944 , \58951 );
xor \U$58919 ( \59262 , \59261 , \58959 );
and \U$58920 ( \59263 , \59260 , \59262 );
and \U$58921 ( \59264 , \59255 , \59260 );
or \U$58922 ( \59265 , \59258 , \59263 , \59264 );
and \U$58923 ( \59266 , \59253 , \59265 );
and \U$58924 ( \59267 , \59172 , \59252 );
or \U$58925 ( \59268 , \59266 , \59267 );
xor \U$58926 ( \59269 , \59116 , \59268 );
xor \U$58927 ( \59270 , \58596 , \58622 );
xor \U$58928 ( \59271 , \59270 , \58648 );
xor \U$58929 ( \59272 , \58849 , \58854 );
xor \U$58930 ( \59273 , \59271 , \59272 );
and \U$58931 ( \59274 , \59269 , \59273 );
and \U$58932 ( \59275 , \59116 , \59268 );
or \U$58933 ( \59276 , \59274 , \59275 );
xor \U$58934 ( \59277 , \58859 , \59023 );
xor \U$58935 ( \59278 , \59277 , \59048 );
and \U$58936 ( \59279 , \59276 , \59278 );
xor \U$58937 ( \59280 , \59053 , \59058 );
xor \U$58938 ( \59281 , \59280 , \59065 );
xor \U$58939 ( \59282 , \58859 , \59023 );
xor \U$58940 ( \59283 , \59282 , \59048 );
and \U$58941 ( \59284 , \59281 , \59283 );
and \U$58942 ( \59285 , \59276 , \59281 );
or \U$58943 ( \59286 , \59279 , \59284 , \59285 );
nand \U$58944 ( \59287 , \59102 , \59286 );
nand \U$58945 ( \59288 , \59101 , \59287 );
and \U$58946 ( \59289 , \59090 , \59288 );
xor \U$58947 ( \59290 , \59288 , \59090 );
xor \U$58948 ( \59291 , \58859 , \59023 );
xor \U$58949 ( \59292 , \59291 , \59048 );
xor \U$58950 ( \59293 , \59276 , \59281 );
xor \U$58951 ( \59294 , \59292 , \59293 );
xor \U$58952 ( \59295 , \58937 , \59010 );
xor \U$58953 ( \59296 , \59295 , \59020 );
xor \U$58954 ( \59297 , \59116 , \59268 );
xor \U$58955 ( \59298 , \59297 , \59273 );
and \U$58956 ( \59299 , \59296 , \59298 );
xor \U$58957 ( \59300 , \59294 , \59299 );
and \U$58958 ( \59301 , \9505 , RI98701c8_80);
and \U$58959 ( \59302 , RI9870fd8_110, \9503 );
nor \U$58960 ( \59303 , \59301 , \59302 );
and \U$58961 ( \59304 , \59303 , \9510 );
not \U$58962 ( \59305 , \59303 );
and \U$58963 ( \59306 , \59305 , \9513 );
nor \U$58964 ( \59307 , \59304 , \59306 );
and \U$58965 ( \59308 , \10424 , RI9870b28_100);
and \U$58966 ( \59309 , RI9870df8_106, \10422 );
nor \U$58967 ( \59310 , \59308 , \59309 );
and \U$58968 ( \59311 , \59310 , \9840 );
not \U$58969 ( \59312 , \59310 );
and \U$58970 ( \59313 , \59312 , \10428 );
nor \U$58971 ( \59314 , \59311 , \59313 );
xor \U$58972 ( \59315 , \59307 , \59314 );
and \U$58973 ( \59316 , \11696 , RI9870a38_98);
and \U$58974 ( \59317 , RI9870ee8_108, \11694 );
nor \U$58975 ( \59318 , \59316 , \59317 );
and \U$58976 ( \59319 , \59318 , \10965 );
not \U$58977 ( \59320 , \59318 );
and \U$58978 ( \59321 , \59320 , \11702 );
nor \U$58979 ( \59322 , \59319 , \59321 );
and \U$58980 ( \59323 , \59315 , \59322 );
and \U$58981 ( \59324 , \59307 , \59314 );
or \U$58982 ( \59325 , \59323 , \59324 );
not \U$58983 ( \59326 , RI9873558_190);
and \U$58984 ( \59327 , \15780 , RI9871848_128);
and \U$58985 ( \59328 , RI9871578_122, RI9873648_192);
nor \U$58986 ( \59329 , \59327 , \59328 );
not \U$58987 ( \59330 , \59329 );
or \U$58988 ( \59331 , \59326 , \59330 );
or \U$58989 ( \59332 , \59329 , RI9873558_190);
nand \U$58990 ( \59333 , \59331 , \59332 );
xor \U$58991 ( \59334 , \59333 , \4521 );
and \U$58992 ( \59335 , \14937 , RI9871488_120);
and \U$58993 ( \59336 , RI9871758_126, \14935 );
nor \U$58994 ( \59337 , \59335 , \59336 );
and \U$58995 ( \59338 , \59337 , \14539 );
not \U$58996 ( \59339 , \59337 );
and \U$58997 ( \59340 , \59339 , \14538 );
nor \U$58998 ( \59341 , \59338 , \59340 );
and \U$58999 ( \59342 , \59334 , \59341 );
and \U$59000 ( \59343 , \59333 , \4521 );
or \U$59001 ( \59344 , \59342 , \59343 );
xor \U$59002 ( \59345 , \59325 , \59344 );
and \U$59003 ( \59346 , \13882 , RI98711b8_114);
and \U$59004 ( \59347 , RI9871398_118, \13880 );
nor \U$59005 ( \59348 , \59346 , \59347 );
and \U$59006 ( \59349 , \59348 , \13358 );
not \U$59007 ( \59350 , \59348 );
and \U$59008 ( \59351 , \59350 , \13359 );
nor \U$59009 ( \59352 , \59349 , \59351 );
and \U$59010 ( \59353 , \12293 , RI9870c18_102);
and \U$59011 ( \59354 , RI98710c8_112, \12291 );
nor \U$59012 ( \59355 , \59353 , \59354 );
and \U$59013 ( \59356 , \59355 , \11687 );
not \U$59014 ( \59357 , \59355 );
and \U$59015 ( \59358 , \59357 , \11686 );
nor \U$59016 ( \59359 , \59356 , \59358 );
xor \U$59017 ( \59360 , \59352 , \59359 );
and \U$59018 ( \59361 , \13045 , RI9870d08_104);
and \U$59019 ( \59362 , RI98712a8_116, \13043 );
nor \U$59020 ( \59363 , \59361 , \59362 );
and \U$59021 ( \59364 , \59363 , \13047 );
not \U$59022 ( \59365 , \59363 );
and \U$59023 ( \59366 , \59365 , \12619 );
nor \U$59024 ( \59367 , \59364 , \59366 );
and \U$59025 ( \59368 , \59360 , \59367 );
and \U$59026 ( \59369 , \59352 , \59359 );
or \U$59027 ( \59370 , \59368 , \59369 );
and \U$59028 ( \59371 , \59345 , \59370 );
and \U$59029 ( \59372 , \59325 , \59344 );
or \U$59030 ( \59373 , \59371 , \59372 );
and \U$59031 ( \59374 , \5881 , RI98702b8_82);
and \U$59032 ( \59375 , RI9870768_92, \5879 );
nor \U$59033 ( \59376 , \59374 , \59375 );
and \U$59034 ( \59377 , \59376 , \5594 );
not \U$59035 ( \59378 , \59376 );
and \U$59036 ( \59379 , \59378 , \5885 );
nor \U$59037 ( \59380 , \59377 , \59379 );
and \U$59038 ( \59381 , \6453 , RI9870678_90);
and \U$59039 ( \59382 , RI9870948_96, \6451 );
nor \U$59040 ( \59383 , \59381 , \59382 );
and \U$59041 ( \59384 , \59383 , \6190 );
not \U$59042 ( \59385 , \59383 );
and \U$59043 ( \59386 , \59385 , \6705 );
nor \U$59044 ( \59387 , \59384 , \59386 );
xor \U$59045 ( \59388 , \59380 , \59387 );
and \U$59046 ( \59389 , \7079 , RI9870858_94);
and \U$59047 ( \59390 , RI986fb38_66, \7077 );
nor \U$59048 ( \59391 , \59389 , \59390 );
and \U$59049 ( \59392 , \59391 , \6710 );
not \U$59050 ( \59393 , \59391 );
and \U$59051 ( \59394 , \59393 , \6709 );
nor \U$59052 ( \59395 , \59392 , \59394 );
and \U$59053 ( \59396 , \59388 , \59395 );
and \U$59054 ( \59397 , \59380 , \59387 );
or \U$59055 ( \59398 , \59396 , \59397 );
not \U$59056 ( \59399 , \4519 );
and \U$59057 ( \59400 , \4710 , RI9870498_86);
and \U$59058 ( \59401 , RI9870588_88, \4708 );
nor \U$59059 ( \59402 , \59400 , \59401 );
not \U$59060 ( \59403 , \59402 );
or \U$59061 ( \59404 , \59399 , \59403 );
or \U$59062 ( \59405 , \59402 , \4521 );
nand \U$59063 ( \59406 , \59404 , \59405 );
xor \U$59064 ( \59407 , \59398 , \59406 );
and \U$59065 ( \59408 , \7729 , RI986fc28_68);
and \U$59066 ( \59409 , RI986fe08_72, \7727 );
nor \U$59067 ( \59410 , \59408 , \59409 );
and \U$59068 ( \59411 , \59410 , \7480 );
not \U$59069 ( \59412 , \59410 );
and \U$59070 ( \59413 , \59412 , \7733 );
nor \U$59071 ( \59414 , \59411 , \59413 );
and \U$59072 ( \59415 , \8486 , RI986fd18_70);
and \U$59073 ( \59416 , RI986ffe8_76, \8484 );
nor \U$59074 ( \59417 , \59415 , \59416 );
and \U$59075 ( \59418 , \59417 , \8050 );
not \U$59076 ( \59419 , \59417 );
and \U$59077 ( \59420 , \59419 , \8051 );
nor \U$59078 ( \59421 , \59418 , \59420 );
xor \U$59079 ( \59422 , \59414 , \59421 );
and \U$59080 ( \59423 , \9237 , RI986fef8_74);
and \U$59081 ( \59424 , RI98700d8_78, \9235 );
nor \U$59082 ( \59425 , \59423 , \59424 );
and \U$59083 ( \59426 , \59425 , \9241 );
not \U$59084 ( \59427 , \59425 );
and \U$59085 ( \59428 , \59427 , \8836 );
nor \U$59086 ( \59429 , \59426 , \59428 );
and \U$59087 ( \59430 , \59422 , \59429 );
and \U$59088 ( \59431 , \59414 , \59421 );
or \U$59089 ( \59432 , \59430 , \59431 );
and \U$59090 ( \59433 , \59407 , \59432 );
and \U$59091 ( \59434 , \59398 , \59406 );
or \U$59092 ( \59435 , \59433 , \59434 );
xor \U$59093 ( \59436 , \59373 , \59435 );
xor \U$59094 ( \59437 , \59148 , \59155 );
xor \U$59095 ( \59438 , \59437 , \59163 );
xor \U$59096 ( \59439 , \59179 , \59186 );
xor \U$59097 ( \59440 , \59439 , \59194 );
and \U$59098 ( \59441 , \59438 , \59440 );
xor \U$59099 ( \59442 , \59123 , \59130 );
xor \U$59100 ( \59443 , \59442 , \59138 );
xor \U$59101 ( \59444 , \59179 , \59186 );
xor \U$59102 ( \59445 , \59444 , \59194 );
and \U$59103 ( \59446 , \59443 , \59445 );
and \U$59104 ( \59447 , \59438 , \59443 );
or \U$59105 ( \59448 , \59441 , \59446 , \59447 );
and \U$59106 ( \59449 , \59436 , \59448 );
and \U$59107 ( \59450 , \59373 , \59435 );
or \U$59108 ( \59451 , \59449 , \59450 );
xor \U$59109 ( \59452 , \59141 , \59166 );
xor \U$59110 ( \59453 , \59452 , \59169 );
xor \U$59111 ( \59454 , \59197 , \59223 );
xor \U$59112 ( \59455 , \59454 , \59249 );
and \U$59113 ( \59456 , \59453 , \59455 );
xor \U$59114 ( \59457 , \59451 , \59456 );
xor \U$59115 ( \59458 , \58970 , \3922 );
xor \U$59116 ( \59459 , \59458 , \58978 );
xor \U$59117 ( \59460 , \58989 , \58996 );
xor \U$59118 ( \59461 , \59460 , \59004 );
xor \U$59119 ( \59462 , \59459 , \59461 );
xor \U$59120 ( \59463 , \58944 , \58951 );
xor \U$59121 ( \59464 , \59463 , \58959 );
xor \U$59122 ( \59465 , \59255 , \59260 );
xor \U$59123 ( \59466 , \59464 , \59465 );
and \U$59124 ( \59467 , \59462 , \59466 );
and \U$59125 ( \59468 , \59459 , \59461 );
or \U$59126 ( \59469 , \59467 , \59468 );
and \U$59127 ( \59470 , \59457 , \59469 );
and \U$59128 ( \59471 , \59451 , \59456 );
or \U$59129 ( \59472 , \59470 , \59471 );
xor \U$59130 ( \59473 , \59036 , \59038 );
xor \U$59131 ( \59474 , \59473 , \59045 );
xor \U$59132 ( \59475 , \59472 , \59474 );
xor \U$59133 ( \59476 , \58962 , \58981 );
xor \U$59134 ( \59477 , \59476 , \59007 );
xor \U$59135 ( \59478 , \59172 , \59252 );
xor \U$59136 ( \59479 , \59478 , \59265 );
and \U$59137 ( \59480 , \59477 , \59479 );
xor \U$59138 ( \59481 , \59013 , \59014 );
xor \U$59139 ( \59482 , \59481 , \59017 );
xor \U$59140 ( \59483 , \59104 , \59111 );
xor \U$59141 ( \59484 , \59482 , \59483 );
xor \U$59142 ( \59485 , \59172 , \59252 );
xor \U$59143 ( \59486 , \59485 , \59265 );
and \U$59144 ( \59487 , \59484 , \59486 );
and \U$59145 ( \59488 , \59477 , \59484 );
or \U$59146 ( \59489 , \59480 , \59487 , \59488 );
and \U$59147 ( \59490 , \59475 , \59489 );
and \U$59148 ( \59491 , \59472 , \59474 );
or \U$59149 ( \59492 , \59490 , \59491 );
xor \U$59150 ( \59493 , \59300 , \59492 );
xor \U$59151 ( \59494 , \59296 , \59298 );
not \U$59152 ( \59495 , \59494 );
xor \U$59153 ( \59496 , \59472 , \59474 );
xor \U$59154 ( \59497 , \59496 , \59489 );
not \U$59155 ( \59498 , \59497 );
or \U$59156 ( \59499 , \59495 , \59498 );
or \U$59157 ( \59500 , \59497 , \59494 );
and \U$59158 ( \59501 , \9505 , RI98700d8_78);
and \U$59159 ( \59502 , RI98701c8_80, \9503 );
nor \U$59160 ( \59503 , \59501 , \59502 );
and \U$59161 ( \59504 , \59503 , \9510 );
not \U$59162 ( \59505 , \59503 );
and \U$59163 ( \59506 , \59505 , \9513 );
nor \U$59164 ( \59507 , \59504 , \59506 );
and \U$59165 ( \59508 , \9237 , RI986ffe8_76);
and \U$59166 ( \59509 , RI986fef8_74, \9235 );
nor \U$59167 ( \59510 , \59508 , \59509 );
and \U$59168 ( \59511 , \59510 , \9241 );
not \U$59169 ( \59512 , \59510 );
and \U$59170 ( \59513 , \59512 , \8836 );
nor \U$59171 ( \59514 , \59511 , \59513 );
xor \U$59172 ( \59515 , \59507 , \59514 );
and \U$59173 ( \59516 , \10424 , RI9870fd8_110);
and \U$59174 ( \59517 , RI9870b28_100, \10422 );
nor \U$59175 ( \59518 , \59516 , \59517 );
and \U$59176 ( \59519 , \59518 , \9840 );
not \U$59177 ( \59520 , \59518 );
and \U$59178 ( \59521 , \59520 , \10428 );
nor \U$59179 ( \59522 , \59519 , \59521 );
and \U$59180 ( \59523 , \59515 , \59522 );
and \U$59181 ( \59524 , \59507 , \59514 );
or \U$59182 ( \59525 , \59523 , \59524 );
and \U$59183 ( \59526 , \13882 , RI98712a8_116);
and \U$59184 ( \59527 , RI98711b8_114, \13880 );
nor \U$59185 ( \59528 , \59526 , \59527 );
and \U$59186 ( \59529 , \59528 , \13358 );
not \U$59187 ( \59530 , \59528 );
and \U$59188 ( \59531 , \59530 , \13359 );
nor \U$59189 ( \59532 , \59529 , \59531 );
not \U$59190 ( \59533 , RI9873558_190);
and \U$59191 ( \59534 , \15780 , RI9871758_126);
and \U$59192 ( \59535 , RI9871848_128, RI9873648_192);
nor \U$59193 ( \59536 , \59534 , \59535 );
not \U$59194 ( \59537 , \59536 );
or \U$59195 ( \59538 , \59533 , \59537 );
or \U$59196 ( \59539 , \59536 , RI9873558_190);
nand \U$59197 ( \59540 , \59538 , \59539 );
xor \U$59198 ( \59541 , \59532 , \59540 );
and \U$59199 ( \59542 , \14937 , RI9871398_118);
and \U$59200 ( \59543 , RI9871488_120, \14935 );
nor \U$59201 ( \59544 , \59542 , \59543 );
and \U$59202 ( \59545 , \59544 , \14539 );
not \U$59203 ( \59546 , \59544 );
and \U$59204 ( \59547 , \59546 , \14538 );
nor \U$59205 ( \59548 , \59545 , \59547 );
and \U$59206 ( \59549 , \59541 , \59548 );
and \U$59207 ( \59550 , \59532 , \59540 );
or \U$59208 ( \59551 , \59549 , \59550 );
xor \U$59209 ( \59552 , \59525 , \59551 );
and \U$59210 ( \59553 , \12293 , RI9870ee8_108);
and \U$59211 ( \59554 , RI9870c18_102, \12291 );
nor \U$59212 ( \59555 , \59553 , \59554 );
and \U$59213 ( \59556 , \59555 , \11687 );
not \U$59214 ( \59557 , \59555 );
and \U$59215 ( \59558 , \59557 , \11686 );
nor \U$59216 ( \59559 , \59556 , \59558 );
and \U$59217 ( \59560 , \11696 , RI9870df8_106);
and \U$59218 ( \59561 , RI9870a38_98, \11694 );
nor \U$59219 ( \59562 , \59560 , \59561 );
and \U$59220 ( \59563 , \59562 , \10965 );
not \U$59221 ( \59564 , \59562 );
and \U$59222 ( \59565 , \59564 , \11702 );
nor \U$59223 ( \59566 , \59563 , \59565 );
xor \U$59224 ( \59567 , \59559 , \59566 );
and \U$59225 ( \59568 , \13045 , RI98710c8_112);
and \U$59226 ( \59569 , RI9870d08_104, \13043 );
nor \U$59227 ( \59570 , \59568 , \59569 );
and \U$59228 ( \59571 , \59570 , \13047 );
not \U$59229 ( \59572 , \59570 );
and \U$59230 ( \59573 , \59572 , \12619 );
nor \U$59231 ( \59574 , \59571 , \59573 );
and \U$59232 ( \59575 , \59567 , \59574 );
and \U$59233 ( \59576 , \59559 , \59566 );
or \U$59234 ( \59577 , \59575 , \59576 );
and \U$59235 ( \59578 , \59552 , \59577 );
and \U$59236 ( \59579 , \59525 , \59551 );
or \U$59237 ( \59580 , \59578 , \59579 );
and \U$59238 ( \59581 , \5318 , RI9870498_86);
and \U$59239 ( \59582 , RI9870588_88, \5316 );
nor \U$59240 ( \59583 , \59581 , \59582 );
and \U$59241 ( \59584 , \59583 , \5052 );
not \U$59242 ( \59585 , \59583 );
and \U$59243 ( \59586 , \59585 , \5322 );
nor \U$59244 ( \59587 , \59584 , \59586 );
and \U$59245 ( \59588 , \5881 , RI98703a8_84);
and \U$59246 ( \59589 , RI98702b8_82, \5879 );
nor \U$59247 ( \59590 , \59588 , \59589 );
and \U$59248 ( \59591 , \59590 , \5594 );
not \U$59249 ( \59592 , \59590 );
and \U$59250 ( \59593 , \59592 , \5885 );
nor \U$59251 ( \59594 , \59591 , \59593 );
xor \U$59252 ( \59595 , \59587 , \59594 );
and \U$59253 ( \59596 , \6453 , RI9870768_92);
and \U$59254 ( \59597 , RI9870678_90, \6451 );
nor \U$59255 ( \59598 , \59596 , \59597 );
and \U$59256 ( \59599 , \59598 , \6190 );
not \U$59257 ( \59600 , \59598 );
and \U$59258 ( \59601 , \59600 , \6180 );
nor \U$59259 ( \59602 , \59599 , \59601 );
and \U$59260 ( \59603 , \59595 , \59602 );
and \U$59261 ( \59604 , \59587 , \59594 );
or \U$59262 ( \59605 , \59603 , \59604 );
and \U$59263 ( \59606 , \5318 , RI9870588_88);
and \U$59264 ( \59607 , RI98703a8_84, \5316 );
nor \U$59265 ( \59608 , \59606 , \59607 );
and \U$59266 ( \59609 , \59608 , \5052 );
not \U$59267 ( \59610 , \59608 );
and \U$59268 ( \59611 , \59610 , \5322 );
nor \U$59269 ( \59612 , \59609 , \59611 );
xor \U$59270 ( \59613 , \59605 , \59612 );
and \U$59271 ( \59614 , \7729 , RI986fb38_66);
and \U$59272 ( \59615 , RI986fc28_68, \7727 );
nor \U$59273 ( \59616 , \59614 , \59615 );
and \U$59274 ( \59617 , \59616 , \7480 );
not \U$59275 ( \59618 , \59616 );
and \U$59276 ( \59619 , \59618 , \7733 );
nor \U$59277 ( \59620 , \59617 , \59619 );
and \U$59278 ( \59621 , \7079 , RI9870948_96);
and \U$59279 ( \59622 , RI9870858_94, \7077 );
nor \U$59280 ( \59623 , \59621 , \59622 );
and \U$59281 ( \59624 , \59623 , \6710 );
not \U$59282 ( \59625 , \59623 );
and \U$59283 ( \59626 , \59625 , \6709 );
nor \U$59284 ( \59627 , \59624 , \59626 );
xor \U$59285 ( \59628 , \59620 , \59627 );
and \U$59286 ( \59629 , \8486 , RI986fe08_72);
and \U$59287 ( \59630 , RI986fd18_70, \8484 );
nor \U$59288 ( \59631 , \59629 , \59630 );
and \U$59289 ( \59632 , \59631 , \8050 );
not \U$59290 ( \59633 , \59631 );
and \U$59291 ( \59634 , \59633 , \8051 );
nor \U$59292 ( \59635 , \59632 , \59634 );
and \U$59293 ( \59636 , \59628 , \59635 );
and \U$59294 ( \59637 , \59620 , \59627 );
or \U$59295 ( \59638 , \59636 , \59637 );
and \U$59296 ( \59639 , \59613 , \59638 );
and \U$59297 ( \59640 , \59605 , \59612 );
or \U$59298 ( \59641 , \59639 , \59640 );
xor \U$59299 ( \59642 , \59580 , \59641 );
xor \U$59300 ( \59643 , \59414 , \59421 );
xor \U$59301 ( \59644 , \59643 , \59429 );
nand \U$59302 ( \59645 , RI9870498_86, \4708 );
not \U$59303 ( \59646 , \59645 );
not \U$59304 ( \59647 , \4519 );
or \U$59305 ( \59648 , \59646 , \59647 );
or \U$59306 ( \59649 , \4519 , \59645 );
nand \U$59307 ( \59650 , \59648 , \59649 );
xor \U$59308 ( \59651 , \59644 , \59650 );
xor \U$59309 ( \59652 , \59380 , \59387 );
xor \U$59310 ( \59653 , \59652 , \59395 );
and \U$59311 ( \59654 , \59651 , \59653 );
and \U$59312 ( \59655 , \59644 , \59650 );
or \U$59313 ( \59656 , \59654 , \59655 );
and \U$59314 ( \59657 , \59642 , \59656 );
and \U$59315 ( \59658 , \59580 , \59641 );
or \U$59316 ( \59659 , \59657 , \59658 );
xor \U$59317 ( \59660 , \59204 , \59212 );
xor \U$59318 ( \59661 , \59660 , \59220 );
xor \U$59319 ( \59662 , \59231 , \59238 );
xor \U$59320 ( \59663 , \59662 , \59246 );
and \U$59321 ( \59664 , \59661 , \59663 );
xor \U$59322 ( \59665 , \59307 , \59314 );
xor \U$59323 ( \59666 , \59665 , \59322 );
xor \U$59324 ( \59667 , \59333 , \4521 );
xor \U$59325 ( \59668 , \59667 , \59341 );
and \U$59326 ( \59669 , \59666 , \59668 );
xor \U$59327 ( \59670 , \59352 , \59359 );
xor \U$59328 ( \59671 , \59670 , \59367 );
xor \U$59329 ( \59672 , \59333 , \4521 );
xor \U$59330 ( \59673 , \59672 , \59341 );
and \U$59331 ( \59674 , \59671 , \59673 );
and \U$59332 ( \59675 , \59666 , \59671 );
or \U$59333 ( \59676 , \59669 , \59674 , \59675 );
xor \U$59334 ( \59677 , \59231 , \59238 );
xor \U$59335 ( \59678 , \59677 , \59246 );
and \U$59336 ( \59679 , \59676 , \59678 );
and \U$59337 ( \59680 , \59661 , \59676 );
or \U$59338 ( \59681 , \59664 , \59679 , \59680 );
xor \U$59339 ( \59682 , \59659 , \59681 );
xor \U$59340 ( \59683 , \59398 , \59406 );
xor \U$59341 ( \59684 , \59683 , \59432 );
xor \U$59342 ( \59685 , \59325 , \59344 );
xor \U$59343 ( \59686 , \59685 , \59370 );
and \U$59344 ( \59687 , \59684 , \59686 );
xor \U$59345 ( \59688 , \59179 , \59186 );
xor \U$59346 ( \59689 , \59688 , \59194 );
xor \U$59347 ( \59690 , \59438 , \59443 );
xor \U$59348 ( \59691 , \59689 , \59690 );
xor \U$59349 ( \59692 , \59325 , \59344 );
xor \U$59350 ( \59693 , \59692 , \59370 );
and \U$59351 ( \59694 , \59691 , \59693 );
and \U$59352 ( \59695 , \59684 , \59691 );
or \U$59353 ( \59696 , \59687 , \59694 , \59695 );
and \U$59354 ( \59697 , \59682 , \59696 );
and \U$59355 ( \59698 , \59659 , \59681 );
or \U$59356 ( \59699 , \59697 , \59698 );
xor \U$59357 ( \59700 , \59453 , \59455 );
xor \U$59358 ( \59701 , \59459 , \59461 );
xor \U$59359 ( \59702 , \59701 , \59466 );
and \U$59360 ( \59703 , \59700 , \59702 );
xor \U$59361 ( \59704 , \59373 , \59435 );
xor \U$59362 ( \59705 , \59704 , \59448 );
xor \U$59363 ( \59706 , \59459 , \59461 );
xor \U$59364 ( \59707 , \59706 , \59466 );
and \U$59365 ( \59708 , \59705 , \59707 );
and \U$59366 ( \59709 , \59700 , \59705 );
or \U$59367 ( \59710 , \59703 , \59708 , \59709 );
xor \U$59368 ( \59711 , \59699 , \59710 );
xor \U$59369 ( \59712 , \59172 , \59252 );
xor \U$59370 ( \59713 , \59712 , \59265 );
xor \U$59371 ( \59714 , \59477 , \59484 );
xor \U$59372 ( \59715 , \59713 , \59714 );
and \U$59373 ( \59716 , \59711 , \59715 );
and \U$59374 ( \59717 , \59699 , \59710 );
or \U$59375 ( \59718 , \59716 , \59717 );
nand \U$59376 ( \59719 , \59500 , \59718 );
nand \U$59377 ( \59720 , \59499 , \59719 );
and \U$59378 ( \59721 , \59493 , \59720 );
xor \U$59379 ( \59722 , \59493 , \59720 );
xnor \U$59380 ( \59723 , \59718 , \59497 );
not \U$59381 ( \59724 , \59723 );
not \U$59382 ( \59725 , \59494 );
and \U$59383 ( \59726 , \59724 , \59725 );
and \U$59384 ( \59727 , \59723 , \59494 );
nor \U$59385 ( \59728 , \59726 , \59727 );
xor \U$59386 ( \59729 , \59699 , \59710 );
xor \U$59387 ( \59730 , \59729 , \59715 );
xor \U$59388 ( \59731 , \59605 , \59612 );
xor \U$59389 ( \59732 , \59731 , \59638 );
xor \U$59390 ( \59733 , \59644 , \59650 );
xor \U$59391 ( \59734 , \59733 , \59653 );
and \U$59392 ( \59735 , \59732 , \59734 );
xor \U$59393 ( \59736 , \59333 , \4521 );
xor \U$59394 ( \59737 , \59736 , \59341 );
xor \U$59395 ( \59738 , \59666 , \59671 );
xor \U$59396 ( \59739 , \59737 , \59738 );
xor \U$59397 ( \59740 , \59644 , \59650 );
xor \U$59398 ( \59741 , \59740 , \59653 );
and \U$59399 ( \59742 , \59739 , \59741 );
and \U$59400 ( \59743 , \59732 , \59739 );
or \U$59401 ( \59744 , \59735 , \59742 , \59743 );
and \U$59402 ( \59745 , \7079 , RI9870678_90);
and \U$59403 ( \59746 , RI9870948_96, \7077 );
nor \U$59404 ( \59747 , \59745 , \59746 );
and \U$59405 ( \59748 , \59747 , \6710 );
not \U$59406 ( \59749 , \59747 );
and \U$59407 ( \59750 , \59749 , \6709 );
nor \U$59408 ( \59751 , \59748 , \59750 );
and \U$59409 ( \59752 , \5881 , RI9870588_88);
and \U$59410 ( \59753 , RI98703a8_84, \5879 );
nor \U$59411 ( \59754 , \59752 , \59753 );
and \U$59412 ( \59755 , \59754 , \5594 );
not \U$59413 ( \59756 , \59754 );
and \U$59414 ( \59757 , \59756 , \5885 );
nor \U$59415 ( \59758 , \59755 , \59757 );
xor \U$59416 ( \59759 , \59751 , \59758 );
and \U$59417 ( \59760 , \6453 , RI98702b8_82);
and \U$59418 ( \59761 , RI9870768_92, \6451 );
nor \U$59419 ( \59762 , \59760 , \59761 );
and \U$59420 ( \59763 , \59762 , \6190 );
not \U$59421 ( \59764 , \59762 );
and \U$59422 ( \59765 , \59764 , \6705 );
nor \U$59423 ( \59766 , \59763 , \59765 );
and \U$59424 ( \59767 , \59759 , \59766 );
and \U$59425 ( \59768 , \59751 , \59758 );
or \U$59426 ( \59769 , \59767 , \59768 );
and \U$59427 ( \59770 , \8486 , RI986fc28_68);
and \U$59428 ( \59771 , RI986fe08_72, \8484 );
nor \U$59429 ( \59772 , \59770 , \59771 );
and \U$59430 ( \59773 , \59772 , \8050 );
not \U$59431 ( \59774 , \59772 );
and \U$59432 ( \59775 , \59774 , \8051 );
nor \U$59433 ( \59776 , \59773 , \59775 );
and \U$59434 ( \59777 , \7729 , RI9870858_94);
and \U$59435 ( \59778 , RI986fb38_66, \7727 );
nor \U$59436 ( \59779 , \59777 , \59778 );
and \U$59437 ( \59780 , \59779 , \7480 );
not \U$59438 ( \59781 , \59779 );
and \U$59439 ( \59782 , \59781 , \7733 );
nor \U$59440 ( \59783 , \59780 , \59782 );
xor \U$59441 ( \59784 , \59776 , \59783 );
and \U$59442 ( \59785 , \9237 , RI986fd18_70);
and \U$59443 ( \59786 , RI986ffe8_76, \9235 );
nor \U$59444 ( \59787 , \59785 , \59786 );
and \U$59445 ( \59788 , \59787 , \9241 );
not \U$59446 ( \59789 , \59787 );
and \U$59447 ( \59790 , \59789 , \8836 );
nor \U$59448 ( \59791 , \59788 , \59790 );
and \U$59449 ( \59792 , \59784 , \59791 );
and \U$59450 ( \59793 , \59776 , \59783 );
or \U$59451 ( \59794 , \59792 , \59793 );
xor \U$59452 ( \59795 , \59769 , \59794 );
xor \U$59453 ( \59796 , \59587 , \59594 );
xor \U$59454 ( \59797 , \59796 , \59602 );
and \U$59455 ( \59798 , \59795 , \59797 );
and \U$59456 ( \59799 , \59769 , \59794 );
or \U$59457 ( \59800 , \59798 , \59799 );
and \U$59458 ( \59801 , \13882 , RI9870d08_104);
and \U$59459 ( \59802 , RI98712a8_116, \13880 );
nor \U$59460 ( \59803 , \59801 , \59802 );
and \U$59461 ( \59804 , \59803 , \13358 );
not \U$59462 ( \59805 , \59803 );
and \U$59463 ( \59806 , \59805 , \13359 );
nor \U$59464 ( \59807 , \59804 , \59806 );
and \U$59465 ( \59808 , \12293 , RI9870a38_98);
and \U$59466 ( \59809 , RI9870ee8_108, \12291 );
nor \U$59467 ( \59810 , \59808 , \59809 );
and \U$59468 ( \59811 , \59810 , \11687 );
not \U$59469 ( \59812 , \59810 );
and \U$59470 ( \59813 , \59812 , \11686 );
nor \U$59471 ( \59814 , \59811 , \59813 );
xor \U$59472 ( \59815 , \59807 , \59814 );
and \U$59473 ( \59816 , \13045 , RI9870c18_102);
and \U$59474 ( \59817 , RI98710c8_112, \13043 );
nor \U$59475 ( \59818 , \59816 , \59817 );
and \U$59476 ( \59819 , \59818 , \13047 );
not \U$59477 ( \59820 , \59818 );
and \U$59478 ( \59821 , \59820 , \12619 );
nor \U$59479 ( \59822 , \59819 , \59821 );
and \U$59480 ( \59823 , \59815 , \59822 );
and \U$59481 ( \59824 , \59807 , \59814 );
or \U$59482 ( \59825 , \59823 , \59824 );
not \U$59483 ( \59826 , RI9873558_190);
and \U$59484 ( \59827 , \15780 , RI9871488_120);
and \U$59485 ( \59828 , RI9871758_126, RI9873648_192);
nor \U$59486 ( \59829 , \59827 , \59828 );
not \U$59487 ( \59830 , \59829 );
or \U$59488 ( \59831 , \59826 , \59830 );
or \U$59489 ( \59832 , \59829 , RI9873558_190);
nand \U$59490 ( \59833 , \59831 , \59832 );
xor \U$59491 ( \59834 , \59833 , \5322 );
and \U$59492 ( \59835 , \14937 , RI98711b8_114);
and \U$59493 ( \59836 , RI9871398_118, \14935 );
nor \U$59494 ( \59837 , \59835 , \59836 );
and \U$59495 ( \59838 , \59837 , \14539 );
not \U$59496 ( \59839 , \59837 );
and \U$59497 ( \59840 , \59839 , \14538 );
nor \U$59498 ( \59841 , \59838 , \59840 );
and \U$59499 ( \59842 , \59834 , \59841 );
and \U$59500 ( \59843 , \59833 , \5322 );
or \U$59501 ( \59844 , \59842 , \59843 );
xor \U$59502 ( \59845 , \59825 , \59844 );
and \U$59503 ( \59846 , \9505 , RI986fef8_74);
and \U$59504 ( \59847 , RI98700d8_78, \9503 );
nor \U$59505 ( \59848 , \59846 , \59847 );
and \U$59506 ( \59849 , \59848 , \9510 );
not \U$59507 ( \59850 , \59848 );
and \U$59508 ( \59851 , \59850 , \9513 );
nor \U$59509 ( \59852 , \59849 , \59851 );
and \U$59510 ( \59853 , \10424 , RI98701c8_80);
and \U$59511 ( \59854 , RI9870fd8_110, \10422 );
nor \U$59512 ( \59855 , \59853 , \59854 );
and \U$59513 ( \59856 , \59855 , \9840 );
not \U$59514 ( \59857 , \59855 );
and \U$59515 ( \59858 , \59857 , \10428 );
nor \U$59516 ( \59859 , \59856 , \59858 );
xor \U$59517 ( \59860 , \59852 , \59859 );
and \U$59518 ( \59861 , \11696 , RI9870b28_100);
and \U$59519 ( \59862 , RI9870df8_106, \11694 );
nor \U$59520 ( \59863 , \59861 , \59862 );
and \U$59521 ( \59864 , \59863 , \10965 );
not \U$59522 ( \59865 , \59863 );
and \U$59523 ( \59866 , \59865 , \11702 );
nor \U$59524 ( \59867 , \59864 , \59866 );
and \U$59525 ( \59868 , \59860 , \59867 );
and \U$59526 ( \59869 , \59852 , \59859 );
or \U$59527 ( \59870 , \59868 , \59869 );
and \U$59528 ( \59871 , \59845 , \59870 );
and \U$59529 ( \59872 , \59825 , \59844 );
or \U$59530 ( \59873 , \59871 , \59872 );
xor \U$59531 ( \59874 , \59800 , \59873 );
xor \U$59532 ( \59875 , \59620 , \59627 );
xor \U$59533 ( \59876 , \59875 , \59635 );
xor \U$59534 ( \59877 , \59507 , \59514 );
xor \U$59535 ( \59878 , \59877 , \59522 );
and \U$59536 ( \59879 , \59876 , \59878 );
xor \U$59537 ( \59880 , \59559 , \59566 );
xor \U$59538 ( \59881 , \59880 , \59574 );
xor \U$59539 ( \59882 , \59507 , \59514 );
xor \U$59540 ( \59883 , \59882 , \59522 );
and \U$59541 ( \59884 , \59881 , \59883 );
and \U$59542 ( \59885 , \59876 , \59881 );
or \U$59543 ( \59886 , \59879 , \59884 , \59885 );
and \U$59544 ( \59887 , \59874 , \59886 );
and \U$59545 ( \59888 , \59800 , \59873 );
or \U$59546 ( \59889 , \59887 , \59888 );
xor \U$59547 ( \59890 , \59744 , \59889 );
xor \U$59548 ( \59891 , \59325 , \59344 );
xor \U$59549 ( \59892 , \59891 , \59370 );
xor \U$59550 ( \59893 , \59684 , \59691 );
xor \U$59551 ( \59894 , \59892 , \59893 );
and \U$59552 ( \59895 , \59890 , \59894 );
and \U$59553 ( \59896 , \59744 , \59889 );
or \U$59554 ( \59897 , \59895 , \59896 );
xor \U$59555 ( \59898 , \59580 , \59641 );
xor \U$59556 ( \59899 , \59898 , \59656 );
xor \U$59557 ( \59900 , \59231 , \59238 );
xor \U$59558 ( \59901 , \59900 , \59246 );
xor \U$59559 ( \59902 , \59661 , \59676 );
xor \U$59560 ( \59903 , \59901 , \59902 );
and \U$59561 ( \59904 , \59899 , \59903 );
xor \U$59562 ( \59905 , \59897 , \59904 );
xor \U$59563 ( \59906 , \59459 , \59461 );
xor \U$59564 ( \59907 , \59906 , \59466 );
xor \U$59565 ( \59908 , \59700 , \59705 );
xor \U$59566 ( \59909 , \59907 , \59908 );
and \U$59567 ( \59910 , \59905 , \59909 );
and \U$59568 ( \59911 , \59897 , \59904 );
or \U$59569 ( \59912 , \59910 , \59911 );
xor \U$59570 ( \59913 , \59730 , \59912 );
xor \U$59571 ( \59914 , \59451 , \59456 );
xor \U$59572 ( \59915 , \59914 , \59469 );
and \U$59573 ( \59916 , \59913 , \59915 );
and \U$59574 ( \59917 , \59730 , \59912 );
nor \U$59575 ( \59918 , \59916 , \59917 );
or \U$59576 ( \59919 , \59728 , \59918 );
xnor \U$59577 ( \59920 , \59918 , \59728 );
and \U$59578 ( \59921 , \7079 , RI9870768_92);
and \U$59579 ( \59922 , RI9870678_90, \7077 );
nor \U$59580 ( \59923 , \59921 , \59922 );
and \U$59581 ( \59924 , \59923 , \6710 );
not \U$59582 ( \59925 , \59923 );
and \U$59583 ( \59926 , \59925 , \6709 );
nor \U$59584 ( \59927 , \59924 , \59926 );
and \U$59585 ( \59928 , \7729 , RI9870948_96);
and \U$59586 ( \59929 , RI9870858_94, \7727 );
nor \U$59587 ( \59930 , \59928 , \59929 );
and \U$59588 ( \59931 , \59930 , \7480 );
not \U$59589 ( \59932 , \59930 );
and \U$59590 ( \59933 , \59932 , \7733 );
nor \U$59591 ( \59934 , \59931 , \59933 );
xor \U$59592 ( \59935 , \59927 , \59934 );
and \U$59593 ( \59936 , \8486 , RI986fb38_66);
and \U$59594 ( \59937 , RI986fc28_68, \8484 );
nor \U$59595 ( \59938 , \59936 , \59937 );
and \U$59596 ( \59939 , \59938 , \8050 );
not \U$59597 ( \59940 , \59938 );
and \U$59598 ( \59941 , \59940 , \8051 );
nor \U$59599 ( \59942 , \59939 , \59941 );
and \U$59600 ( \59943 , \59935 , \59942 );
and \U$59601 ( \59944 , \59927 , \59934 );
or \U$59602 ( \59945 , \59943 , \59944 );
nand \U$59603 ( \59946 , RI9870498_86, \5316 );
and \U$59604 ( \59947 , \59946 , \5052 );
not \U$59605 ( \59948 , \59946 );
and \U$59606 ( \59949 , \59948 , \5322 );
nor \U$59607 ( \59950 , \59947 , \59949 );
xor \U$59608 ( \59951 , \59945 , \59950 );
xor \U$59609 ( \59952 , \59751 , \59758 );
xor \U$59610 ( \59953 , \59952 , \59766 );
and \U$59611 ( \59954 , \59951 , \59953 );
and \U$59612 ( \59955 , \59945 , \59950 );
or \U$59613 ( \59956 , \59954 , \59955 );
and \U$59614 ( \59957 , \9237 , RI986fe08_72);
and \U$59615 ( \59958 , RI986fd18_70, \9235 );
nor \U$59616 ( \59959 , \59957 , \59958 );
and \U$59617 ( \59960 , \59959 , \9241 );
not \U$59618 ( \59961 , \59959 );
and \U$59619 ( \59962 , \59961 , \8836 );
nor \U$59620 ( \59963 , \59960 , \59962 );
and \U$59621 ( \59964 , \9505 , RI986ffe8_76);
and \U$59622 ( \59965 , RI986fef8_74, \9503 );
nor \U$59623 ( \59966 , \59964 , \59965 );
and \U$59624 ( \59967 , \59966 , \9510 );
not \U$59625 ( \59968 , \59966 );
and \U$59626 ( \59969 , \59968 , \9513 );
nor \U$59627 ( \59970 , \59967 , \59969 );
xor \U$59628 ( \59971 , \59963 , \59970 );
and \U$59629 ( \59972 , \10424 , RI98700d8_78);
and \U$59630 ( \59973 , RI98701c8_80, \10422 );
nor \U$59631 ( \59974 , \59972 , \59973 );
and \U$59632 ( \59975 , \59974 , \9840 );
not \U$59633 ( \59976 , \59974 );
and \U$59634 ( \59977 , \59976 , \10428 );
nor \U$59635 ( \59978 , \59975 , \59977 );
and \U$59636 ( \59979 , \59971 , \59978 );
and \U$59637 ( \59980 , \59963 , \59970 );
or \U$59638 ( \59981 , \59979 , \59980 );
and \U$59639 ( \59982 , \13882 , RI98710c8_112);
and \U$59640 ( \59983 , RI9870d08_104, \13880 );
nor \U$59641 ( \59984 , \59982 , \59983 );
and \U$59642 ( \59985 , \59984 , \13358 );
not \U$59643 ( \59986 , \59984 );
and \U$59644 ( \59987 , \59986 , \13359 );
nor \U$59645 ( \59988 , \59985 , \59987 );
not \U$59646 ( \59989 , RI9873558_190);
and \U$59647 ( \59990 , \15780 , RI9871398_118);
and \U$59648 ( \59991 , RI9871488_120, RI9873648_192);
nor \U$59649 ( \59992 , \59990 , \59991 );
not \U$59650 ( \59993 , \59992 );
or \U$59651 ( \59994 , \59989 , \59993 );
or \U$59652 ( \59995 , \59992 , RI9873558_190);
nand \U$59653 ( \59996 , \59994 , \59995 );
xor \U$59654 ( \59997 , \59988 , \59996 );
and \U$59655 ( \59998 , \14937 , RI98712a8_116);
and \U$59656 ( \59999 , RI98711b8_114, \14935 );
nor \U$59657 ( \60000 , \59998 , \59999 );
and \U$59658 ( \60001 , \60000 , \14539 );
not \U$59659 ( \60002 , \60000 );
and \U$59660 ( \60003 , \60002 , \14538 );
nor \U$59661 ( \60004 , \60001 , \60003 );
and \U$59662 ( \60005 , \59997 , \60004 );
and \U$59663 ( \60006 , \59988 , \59996 );
or \U$59664 ( \60007 , \60005 , \60006 );
xor \U$59665 ( \60008 , \59981 , \60007 );
and \U$59666 ( \60009 , \12293 , RI9870df8_106);
and \U$59667 ( \60010 , RI9870a38_98, \12291 );
nor \U$59668 ( \60011 , \60009 , \60010 );
and \U$59669 ( \60012 , \60011 , \11687 );
not \U$59670 ( \60013 , \60011 );
and \U$59671 ( \60014 , \60013 , \11686 );
nor \U$59672 ( \60015 , \60012 , \60014 );
and \U$59673 ( \60016 , \11696 , RI9870fd8_110);
and \U$59674 ( \60017 , RI9870b28_100, \11694 );
nor \U$59675 ( \60018 , \60016 , \60017 );
and \U$59676 ( \60019 , \60018 , \10965 );
not \U$59677 ( \60020 , \60018 );
and \U$59678 ( \60021 , \60020 , \11702 );
nor \U$59679 ( \60022 , \60019 , \60021 );
xor \U$59680 ( \60023 , \60015 , \60022 );
and \U$59681 ( \60024 , \13045 , RI9870ee8_108);
and \U$59682 ( \60025 , RI9870c18_102, \13043 );
nor \U$59683 ( \60026 , \60024 , \60025 );
and \U$59684 ( \60027 , \60026 , \13047 );
not \U$59685 ( \60028 , \60026 );
and \U$59686 ( \60029 , \60028 , \12619 );
nor \U$59687 ( \60030 , \60027 , \60029 );
and \U$59688 ( \60031 , \60023 , \60030 );
and \U$59689 ( \60032 , \60015 , \60022 );
or \U$59690 ( \60033 , \60031 , \60032 );
and \U$59691 ( \60034 , \60008 , \60033 );
and \U$59692 ( \60035 , \59981 , \60007 );
or \U$59693 ( \60036 , \60034 , \60035 );
xor \U$59694 ( \60037 , \59956 , \60036 );
xor \U$59695 ( \60038 , \59852 , \59859 );
xor \U$59696 ( \60039 , \60038 , \59867 );
xor \U$59697 ( \60040 , \59776 , \59783 );
xor \U$59698 ( \60041 , \60040 , \59791 );
and \U$59699 ( \60042 , \60039 , \60041 );
xor \U$59700 ( \60043 , \59807 , \59814 );
xor \U$59701 ( \60044 , \60043 , \59822 );
xor \U$59702 ( \60045 , \59776 , \59783 );
xor \U$59703 ( \60046 , \60045 , \59791 );
and \U$59704 ( \60047 , \60044 , \60046 );
and \U$59705 ( \60048 , \60039 , \60044 );
or \U$59706 ( \60049 , \60042 , \60047 , \60048 );
xor \U$59707 ( \60050 , \60037 , \60049 );
xor \U$59708 ( \60051 , \59769 , \59794 );
xor \U$59709 ( \60052 , \60051 , \59797 );
xor \U$59710 ( \60053 , \59532 , \59540 );
xor \U$59711 ( \60054 , \60053 , \59548 );
xor \U$59712 ( \60055 , \59507 , \59514 );
xor \U$59713 ( \60056 , \60055 , \59522 );
xor \U$59714 ( \60057 , \59876 , \59881 );
xor \U$59715 ( \60058 , \60056 , \60057 );
xor \U$59716 ( \60059 , \60054 , \60058 );
xor \U$59717 ( \60060 , \60052 , \60059 );
and \U$59718 ( \60061 , \60050 , \60060 );
xor \U$59719 ( \60062 , \59644 , \59650 );
xor \U$59720 ( \60063 , \60062 , \59653 );
xor \U$59721 ( \60064 , \59732 , \59739 );
xor \U$59722 ( \60065 , \60063 , \60064 );
xor \U$59723 ( \60066 , \60061 , \60065 );
and \U$59724 ( \60067 , \9505 , RI986fd18_70);
and \U$59725 ( \60068 , RI986ffe8_76, \9503 );
nor \U$59726 ( \60069 , \60067 , \60068 );
and \U$59727 ( \60070 , \60069 , \9510 );
not \U$59728 ( \60071 , \60069 );
and \U$59729 ( \60072 , \60071 , \9513 );
nor \U$59730 ( \60073 , \60070 , \60072 );
and \U$59731 ( \60074 , \10424 , RI986fef8_74);
and \U$59732 ( \60075 , RI98700d8_78, \10422 );
nor \U$59733 ( \60076 , \60074 , \60075 );
and \U$59734 ( \60077 , \60076 , \9840 );
not \U$59735 ( \60078 , \60076 );
and \U$59736 ( \60079 , \60078 , \10428 );
nor \U$59737 ( \60080 , \60077 , \60079 );
xor \U$59738 ( \60081 , \60073 , \60080 );
and \U$59739 ( \60082 , \11696 , RI98701c8_80);
and \U$59740 ( \60083 , RI9870fd8_110, \11694 );
nor \U$59741 ( \60084 , \60082 , \60083 );
and \U$59742 ( \60085 , \60084 , \10965 );
not \U$59743 ( \60086 , \60084 );
and \U$59744 ( \60087 , \60086 , \11702 );
nor \U$59745 ( \60088 , \60085 , \60087 );
and \U$59746 ( \60089 , \60081 , \60088 );
and \U$59747 ( \60090 , \60073 , \60080 );
or \U$59748 ( \60091 , \60089 , \60090 );
not \U$59749 ( \60092 , RI9873558_190);
and \U$59750 ( \60093 , \15780 , RI98711b8_114);
and \U$59751 ( \60094 , RI9871398_118, RI9873648_192);
nor \U$59752 ( \60095 , \60093 , \60094 );
not \U$59753 ( \60096 , \60095 );
or \U$59754 ( \60097 , \60092 , \60096 );
or \U$59755 ( \60098 , \60095 , RI9873558_190);
nand \U$59756 ( \60099 , \60097 , \60098 );
xor \U$59757 ( \60100 , \60099 , \5885 );
and \U$59758 ( \60101 , \14937 , RI9870d08_104);
and \U$59759 ( \60102 , RI98712a8_116, \14935 );
nor \U$59760 ( \60103 , \60101 , \60102 );
and \U$59761 ( \60104 , \60103 , \14539 );
not \U$59762 ( \60105 , \60103 );
and \U$59763 ( \60106 , \60105 , \14538 );
nor \U$59764 ( \60107 , \60104 , \60106 );
and \U$59765 ( \60108 , \60100 , \60107 );
and \U$59766 ( \60109 , \60099 , \5885 );
or \U$59767 ( \60110 , \60108 , \60109 );
xor \U$59768 ( \60111 , \60091 , \60110 );
and \U$59769 ( \60112 , \12293 , RI9870b28_100);
and \U$59770 ( \60113 , RI9870df8_106, \12291 );
nor \U$59771 ( \60114 , \60112 , \60113 );
and \U$59772 ( \60115 , \60114 , \11687 );
not \U$59773 ( \60116 , \60114 );
and \U$59774 ( \60117 , \60116 , \11686 );
nor \U$59775 ( \60118 , \60115 , \60117 );
and \U$59776 ( \60119 , \13045 , RI9870a38_98);
and \U$59777 ( \60120 , RI9870ee8_108, \13043 );
nor \U$59778 ( \60121 , \60119 , \60120 );
and \U$59779 ( \60122 , \60121 , \13047 );
not \U$59780 ( \60123 , \60121 );
and \U$59781 ( \60124 , \60123 , \12619 );
nor \U$59782 ( \60125 , \60122 , \60124 );
xor \U$59783 ( \60126 , \60118 , \60125 );
and \U$59784 ( \60127 , \13882 , RI9870c18_102);
and \U$59785 ( \60128 , RI98710c8_112, \13880 );
nor \U$59786 ( \60129 , \60127 , \60128 );
and \U$59787 ( \60130 , \60129 , \13358 );
not \U$59788 ( \60131 , \60129 );
and \U$59789 ( \60132 , \60131 , \13359 );
nor \U$59790 ( \60133 , \60130 , \60132 );
and \U$59791 ( \60134 , \60126 , \60133 );
and \U$59792 ( \60135 , \60118 , \60125 );
or \U$59793 ( \60136 , \60134 , \60135 );
and \U$59794 ( \60137 , \60111 , \60136 );
and \U$59795 ( \60138 , \60091 , \60110 );
or \U$59796 ( \60139 , \60137 , \60138 );
and \U$59797 ( \60140 , \7079 , RI98702b8_82);
and \U$59798 ( \60141 , RI9870768_92, \7077 );
nor \U$59799 ( \60142 , \60140 , \60141 );
and \U$59800 ( \60143 , \60142 , \6710 );
not \U$59801 ( \60144 , \60142 );
and \U$59802 ( \60145 , \60144 , \6709 );
nor \U$59803 ( \60146 , \60143 , \60145 );
nand \U$59804 ( \60147 , RI9870498_86, \5879 );
and \U$59805 ( \60148 , \60147 , \5594 );
not \U$59806 ( \60149 , \60147 );
and \U$59807 ( \60150 , \60149 , \5885 );
nor \U$59808 ( \60151 , \60148 , \60150 );
xor \U$59809 ( \60152 , \60146 , \60151 );
and \U$59810 ( \60153 , \6453 , RI9870588_88);
and \U$59811 ( \60154 , RI98703a8_84, \6451 );
nor \U$59812 ( \60155 , \60153 , \60154 );
and \U$59813 ( \60156 , \60155 , \6190 );
not \U$59814 ( \60157 , \60155 );
and \U$59815 ( \60158 , \60157 , \6705 );
nor \U$59816 ( \60159 , \60156 , \60158 );
and \U$59817 ( \60160 , \60152 , \60159 );
and \U$59818 ( \60161 , \60146 , \60151 );
or \U$59819 ( \60162 , \60160 , \60161 );
and \U$59820 ( \60163 , \6453 , RI98703a8_84);
and \U$59821 ( \60164 , RI98702b8_82, \6451 );
nor \U$59822 ( \60165 , \60163 , \60164 );
and \U$59823 ( \60166 , \60165 , \6190 );
not \U$59824 ( \60167 , \60165 );
and \U$59825 ( \60168 , \60167 , \6705 );
nor \U$59826 ( \60169 , \60166 , \60168 );
xor \U$59827 ( \60170 , \60162 , \60169 );
and \U$59828 ( \60171 , \8486 , RI9870858_94);
and \U$59829 ( \60172 , RI986fb38_66, \8484 );
nor \U$59830 ( \60173 , \60171 , \60172 );
and \U$59831 ( \60174 , \60173 , \8050 );
not \U$59832 ( \60175 , \60173 );
and \U$59833 ( \60176 , \60175 , \8051 );
nor \U$59834 ( \60177 , \60174 , \60176 );
and \U$59835 ( \60178 , \7729 , RI9870678_90);
and \U$59836 ( \60179 , RI9870948_96, \7727 );
nor \U$59837 ( \60180 , \60178 , \60179 );
and \U$59838 ( \60181 , \60180 , \7480 );
not \U$59839 ( \60182 , \60180 );
and \U$59840 ( \60183 , \60182 , \7733 );
nor \U$59841 ( \60184 , \60181 , \60183 );
xor \U$59842 ( \60185 , \60177 , \60184 );
and \U$59843 ( \60186 , \9237 , RI986fc28_68);
and \U$59844 ( \60187 , RI986fe08_72, \9235 );
nor \U$59845 ( \60188 , \60186 , \60187 );
and \U$59846 ( \60189 , \60188 , \9241 );
not \U$59847 ( \60190 , \60188 );
and \U$59848 ( \60191 , \60190 , \8836 );
nor \U$59849 ( \60192 , \60189 , \60191 );
and \U$59850 ( \60193 , \60185 , \60192 );
and \U$59851 ( \60194 , \60177 , \60184 );
or \U$59852 ( \60195 , \60193 , \60194 );
and \U$59853 ( \60196 , \60170 , \60195 );
and \U$59854 ( \60197 , \60162 , \60169 );
or \U$59855 ( \60198 , \60196 , \60197 );
xor \U$59856 ( \60199 , \60139 , \60198 );
and \U$59857 ( \60200 , \5881 , RI9870498_86);
and \U$59858 ( \60201 , RI9870588_88, \5879 );
nor \U$59859 ( \60202 , \60200 , \60201 );
and \U$59860 ( \60203 , \60202 , \5594 );
not \U$59861 ( \60204 , \60202 );
and \U$59862 ( \60205 , \60204 , \5885 );
nor \U$59863 ( \60206 , \60203 , \60205 );
xor \U$59864 ( \60207 , \59927 , \59934 );
xor \U$59865 ( \60208 , \60207 , \59942 );
and \U$59866 ( \60209 , \60206 , \60208 );
xor \U$59867 ( \60210 , \59963 , \59970 );
xor \U$59868 ( \60211 , \60210 , \59978 );
xor \U$59869 ( \60212 , \59927 , \59934 );
xor \U$59870 ( \60213 , \60212 , \59942 );
and \U$59871 ( \60214 , \60211 , \60213 );
and \U$59872 ( \60215 , \60206 , \60211 );
or \U$59873 ( \60216 , \60209 , \60214 , \60215 );
and \U$59874 ( \60217 , \60199 , \60216 );
and \U$59875 ( \60218 , \60139 , \60198 );
or \U$59876 ( \60219 , \60217 , \60218 );
xor \U$59877 ( \60220 , \59825 , \59844 );
xor \U$59878 ( \60221 , \60220 , \59870 );
xor \U$59879 ( \60222 , \60219 , \60221 );
xor \U$59880 ( \60223 , \59833 , \5322 );
xor \U$59881 ( \60224 , \60223 , \59841 );
xor \U$59882 ( \60225 , \59945 , \59950 );
xor \U$59883 ( \60226 , \60225 , \59953 );
and \U$59884 ( \60227 , \60224 , \60226 );
xor \U$59885 ( \60228 , \59776 , \59783 );
xor \U$59886 ( \60229 , \60228 , \59791 );
xor \U$59887 ( \60230 , \60039 , \60044 );
xor \U$59888 ( \60231 , \60229 , \60230 );
xor \U$59889 ( \60232 , \59945 , \59950 );
xor \U$59890 ( \60233 , \60232 , \59953 );
and \U$59891 ( \60234 , \60231 , \60233 );
and \U$59892 ( \60235 , \60224 , \60231 );
or \U$59893 ( \60236 , \60227 , \60234 , \60235 );
and \U$59894 ( \60237 , \60222 , \60236 );
and \U$59895 ( \60238 , \60219 , \60221 );
or \U$59896 ( \60239 , \60237 , \60238 );
and \U$59897 ( \60240 , \60066 , \60239 );
and \U$59898 ( \60241 , \60061 , \60065 );
or \U$59899 ( \60242 , \60240 , \60241 );
xor \U$59900 ( \60243 , \59800 , \59873 );
xor \U$59901 ( \60244 , \60243 , \59886 );
xor \U$59902 ( \60245 , \59956 , \60036 );
and \U$59903 ( \60246 , \60245 , \60049 );
and \U$59904 ( \60247 , \59956 , \60036 );
or \U$59905 ( \60248 , \60246 , \60247 );
xor \U$59906 ( \60249 , \59525 , \59551 );
xor \U$59907 ( \60250 , \60249 , \59577 );
xor \U$59908 ( \60251 , \60248 , \60250 );
xor \U$59909 ( \60252 , \59769 , \59794 );
xor \U$59910 ( \60253 , \60252 , \59797 );
and \U$59911 ( \60254 , \60054 , \60253 );
xor \U$59912 ( \60255 , \59769 , \59794 );
xor \U$59913 ( \60256 , \60255 , \59797 );
and \U$59914 ( \60257 , \60058 , \60256 );
and \U$59915 ( \60258 , \60054 , \60058 );
or \U$59916 ( \60259 , \60254 , \60257 , \60258 );
xor \U$59917 ( \60260 , \60251 , \60259 );
and \U$59918 ( \60261 , \60244 , \60260 );
xor \U$59919 ( \60262 , \60242 , \60261 );
xor \U$59920 ( \60263 , \60248 , \60250 );
and \U$59921 ( \60264 , \60263 , \60259 );
and \U$59922 ( \60265 , \60248 , \60250 );
or \U$59923 ( \60266 , \60264 , \60265 );
xor \U$59924 ( \60267 , \59899 , \59903 );
xor \U$59925 ( \60268 , \60266 , \60267 );
xor \U$59926 ( \60269 , \59744 , \59889 );
xor \U$59927 ( \60270 , \60269 , \59894 );
xor \U$59928 ( \60271 , \60268 , \60270 );
and \U$59929 ( \60272 , \60262 , \60271 );
and \U$59930 ( \60273 , \60242 , \60261 );
nor \U$59931 ( \60274 , \60272 , \60273 );
xor \U$59932 ( \60275 , \59659 , \59681 );
xor \U$59933 ( \60276 , \60275 , \59696 );
xor \U$59934 ( \60277 , \60266 , \60267 );
and \U$59935 ( \60278 , \60277 , \60270 );
and \U$59936 ( \60279 , \60266 , \60267 );
or \U$59937 ( \60280 , \60278 , \60279 );
xnor \U$59938 ( \60281 , \60276 , \60280 );
not \U$59939 ( \60282 , \60281 );
xor \U$59940 ( \60283 , \59897 , \59904 );
xor \U$59941 ( \60284 , \60283 , \59909 );
not \U$59942 ( \60285 , \60284 );
and \U$59943 ( \60286 , \60282 , \60285 );
and \U$59944 ( \60287 , \60281 , \60284 );
nor \U$59945 ( \60288 , \60286 , \60287 );
or \U$59946 ( \60289 , \60274 , \60288 );
xnor \U$59947 ( \60290 , \60288 , \60274 );
xor \U$59948 ( \60291 , \60242 , \60261 );
xor \U$59949 ( \60292 , \60291 , \60271 );
xor \U$59950 ( \60293 , \60244 , \60260 );
not \U$59951 ( \60294 , \60293 );
xor \U$59952 ( \60295 , \60061 , \60065 );
xor \U$59953 ( \60296 , \60295 , \60239 );
not \U$59954 ( \60297 , \60296 );
or \U$59955 ( \60298 , \60294 , \60297 );
or \U$59956 ( \60299 , \60296 , \60293 );
xor \U$59957 ( \60300 , \60050 , \60060 );
xor \U$59958 ( \60301 , \60015 , \60022 );
xor \U$59959 ( \60302 , \60301 , \60030 );
xor \U$59960 ( \60303 , \59988 , \59996 );
xor \U$59961 ( \60304 , \60303 , \60004 );
xor \U$59962 ( \60305 , \60302 , \60304 );
xor \U$59963 ( \60306 , \59927 , \59934 );
xor \U$59964 ( \60307 , \60306 , \59942 );
xor \U$59965 ( \60308 , \60206 , \60211 );
xor \U$59966 ( \60309 , \60307 , \60308 );
and \U$59967 ( \60310 , \60305 , \60309 );
and \U$59968 ( \60311 , \60302 , \60304 );
or \U$59969 ( \60312 , \60310 , \60311 );
xor \U$59970 ( \60313 , \59981 , \60007 );
xor \U$59971 ( \60314 , \60313 , \60033 );
xor \U$59972 ( \60315 , \60312 , \60314 );
xor \U$59973 ( \60316 , \60146 , \60151 );
xor \U$59974 ( \60317 , \60316 , \60159 );
and \U$59975 ( \60318 , \7079 , RI98703a8_84);
and \U$59976 ( \60319 , RI98702b8_82, \7077 );
nor \U$59977 ( \60320 , \60318 , \60319 );
and \U$59978 ( \60321 , \60320 , \6709 );
not \U$59979 ( \60322 , \60320 );
and \U$59980 ( \60323 , \60322 , \6710 );
nor \U$59981 ( \60324 , \60321 , \60323 );
and \U$59982 ( \60325 , \7729 , RI9870768_92);
and \U$59983 ( \60326 , RI9870678_90, \7727 );
nor \U$59984 ( \60327 , \60325 , \60326 );
and \U$59985 ( \60328 , \60327 , \7733 );
not \U$59986 ( \60329 , \60327 );
and \U$59987 ( \60330 , \60329 , \7480 );
nor \U$59988 ( \60331 , \60328 , \60330 );
or \U$59989 ( \60332 , \60324 , \60331 );
not \U$59990 ( \60333 , \60331 );
not \U$59991 ( \60334 , \60324 );
or \U$59992 ( \60335 , \60333 , \60334 );
and \U$59993 ( \60336 , \8486 , RI9870948_96);
and \U$59994 ( \60337 , RI9870858_94, \8484 );
nor \U$59995 ( \60338 , \60336 , \60337 );
and \U$59996 ( \60339 , \60338 , \8050 );
not \U$59997 ( \60340 , \60338 );
and \U$59998 ( \60341 , \60340 , \8051 );
nor \U$59999 ( \60342 , \60339 , \60341 );
nand \U$60000 ( \60343 , \60335 , \60342 );
nand \U$60001 ( \60344 , \60332 , \60343 );
xor \U$60002 ( \60345 , \60317 , \60344 );
xor \U$60003 ( \60346 , \60177 , \60184 );
xor \U$60004 ( \60347 , \60346 , \60192 );
and \U$60005 ( \60348 , \60345 , \60347 );
and \U$60006 ( \60349 , \60317 , \60344 );
or \U$60007 ( \60350 , \60348 , \60349 );
and \U$60008 ( \60351 , \13045 , RI9870df8_106);
and \U$60009 ( \60352 , RI9870a38_98, \13043 );
nor \U$60010 ( \60353 , \60351 , \60352 );
and \U$60011 ( \60354 , \60353 , \13047 );
not \U$60012 ( \60355 , \60353 );
and \U$60013 ( \60356 , \60355 , \12619 );
nor \U$60014 ( \60357 , \60354 , \60356 );
and \U$60015 ( \60358 , \11696 , RI98700d8_78);
and \U$60016 ( \60359 , RI98701c8_80, \11694 );
nor \U$60017 ( \60360 , \60358 , \60359 );
and \U$60018 ( \60361 , \60360 , \10965 );
not \U$60019 ( \60362 , \60360 );
and \U$60020 ( \60363 , \60362 , \11702 );
nor \U$60021 ( \60364 , \60361 , \60363 );
xor \U$60022 ( \60365 , \60357 , \60364 );
and \U$60023 ( \60366 , \12293 , RI9870fd8_110);
and \U$60024 ( \60367 , RI9870b28_100, \12291 );
nor \U$60025 ( \60368 , \60366 , \60367 );
and \U$60026 ( \60369 , \60368 , \11687 );
not \U$60027 ( \60370 , \60368 );
and \U$60028 ( \60371 , \60370 , \11686 );
nor \U$60029 ( \60372 , \60369 , \60371 );
and \U$60030 ( \60373 , \60365 , \60372 );
and \U$60031 ( \60374 , \60357 , \60364 );
or \U$60032 ( \60375 , \60373 , \60374 );
and \U$60033 ( \60376 , \13882 , RI9870ee8_108);
and \U$60034 ( \60377 , RI9870c18_102, \13880 );
nor \U$60035 ( \60378 , \60376 , \60377 );
and \U$60036 ( \60379 , \60378 , \13359 );
not \U$60037 ( \60380 , \60378 );
and \U$60038 ( \60381 , \60380 , \13358 );
nor \U$60039 ( \60382 , \60379 , \60381 );
and \U$60040 ( \60383 , \15780 , RI98712a8_116);
and \U$60041 ( \60384 , RI98711b8_114, RI9873648_192);
nor \U$60042 ( \60385 , \60383 , \60384 );
not \U$60043 ( \60386 , \60385 );
not \U$60044 ( \60387 , RI9873558_190);
and \U$60045 ( \60388 , \60386 , \60387 );
and \U$60046 ( \60389 , \60385 , RI9873558_190);
nor \U$60047 ( \60390 , \60388 , \60389 );
or \U$60048 ( \60391 , \60382 , \60390 );
not \U$60049 ( \60392 , \60390 );
not \U$60050 ( \60393 , \60382 );
or \U$60051 ( \60394 , \60392 , \60393 );
and \U$60052 ( \60395 , \14937 , RI98710c8_112);
and \U$60053 ( \60396 , RI9870d08_104, \14935 );
nor \U$60054 ( \60397 , \60395 , \60396 );
and \U$60055 ( \60398 , \60397 , \14539 );
not \U$60056 ( \60399 , \60397 );
and \U$60057 ( \60400 , \60399 , \14538 );
nor \U$60058 ( \60401 , \60398 , \60400 );
nand \U$60059 ( \60402 , \60394 , \60401 );
nand \U$60060 ( \60403 , \60391 , \60402 );
xor \U$60061 ( \60404 , \60375 , \60403 );
and \U$60062 ( \60405 , \9237 , RI986fb38_66);
and \U$60063 ( \60406 , RI986fc28_68, \9235 );
nor \U$60064 ( \60407 , \60405 , \60406 );
and \U$60065 ( \60408 , \60407 , \8836 );
not \U$60066 ( \60409 , \60407 );
and \U$60067 ( \60410 , \60409 , \9241 );
nor \U$60068 ( \60411 , \60408 , \60410 );
and \U$60069 ( \60412 , \9505 , RI986fe08_72);
and \U$60070 ( \60413 , RI986fd18_70, \9503 );
nor \U$60071 ( \60414 , \60412 , \60413 );
and \U$60072 ( \60415 , \60414 , \9513 );
not \U$60073 ( \60416 , \60414 );
and \U$60074 ( \60417 , \60416 , \9510 );
nor \U$60075 ( \60418 , \60415 , \60417 );
or \U$60076 ( \60419 , \60411 , \60418 );
not \U$60077 ( \60420 , \60418 );
not \U$60078 ( \60421 , \60411 );
or \U$60079 ( \60422 , \60420 , \60421 );
and \U$60080 ( \60423 , \10424 , RI986ffe8_76);
and \U$60081 ( \60424 , RI986fef8_74, \10422 );
nor \U$60082 ( \60425 , \60423 , \60424 );
and \U$60083 ( \60426 , \60425 , \9840 );
not \U$60084 ( \60427 , \60425 );
and \U$60085 ( \60428 , \60427 , \10428 );
nor \U$60086 ( \60429 , \60426 , \60428 );
nand \U$60087 ( \60430 , \60422 , \60429 );
nand \U$60088 ( \60431 , \60419 , \60430 );
and \U$60089 ( \60432 , \60404 , \60431 );
and \U$60090 ( \60433 , \60375 , \60403 );
or \U$60091 ( \60434 , \60432 , \60433 );
xor \U$60092 ( \60435 , \60350 , \60434 );
xor \U$60093 ( \60436 , \60073 , \60080 );
xor \U$60094 ( \60437 , \60436 , \60088 );
xor \U$60095 ( \60438 , \60118 , \60125 );
xor \U$60096 ( \60439 , \60438 , \60133 );
and \U$60097 ( \60440 , \60437 , \60439 );
xor \U$60098 ( \60441 , \60099 , \5885 );
xor \U$60099 ( \60442 , \60441 , \60107 );
xor \U$60100 ( \60443 , \60118 , \60125 );
xor \U$60101 ( \60444 , \60443 , \60133 );
and \U$60102 ( \60445 , \60442 , \60444 );
and \U$60103 ( \60446 , \60437 , \60442 );
or \U$60104 ( \60447 , \60440 , \60445 , \60446 );
and \U$60105 ( \60448 , \60435 , \60447 );
and \U$60106 ( \60449 , \60350 , \60434 );
or \U$60107 ( \60450 , \60448 , \60449 );
and \U$60108 ( \60451 , \60315 , \60450 );
and \U$60109 ( \60452 , \60312 , \60314 );
or \U$60110 ( \60453 , \60451 , \60452 );
xor \U$60111 ( \60454 , \60300 , \60453 );
xor \U$60112 ( \60455 , \60219 , \60221 );
xor \U$60113 ( \60456 , \60455 , \60236 );
and \U$60114 ( \60457 , \60454 , \60456 );
and \U$60115 ( \60458 , \60300 , \60453 );
or \U$60116 ( \60459 , \60457 , \60458 );
nand \U$60117 ( \60460 , \60299 , \60459 );
nand \U$60118 ( \60461 , \60298 , \60460 );
and \U$60119 ( \60462 , \60292 , \60461 );
xor \U$60120 ( \60463 , \60461 , \60292 );
and \U$60121 ( \60464 , \9237 , RI9870858_94);
and \U$60122 ( \60465 , RI986fb38_66, \9235 );
nor \U$60123 ( \60466 , \60464 , \60465 );
and \U$60124 ( \60467 , \60466 , \9241 );
not \U$60125 ( \60468 , \60466 );
and \U$60126 ( \60469 , \60468 , \8836 );
nor \U$60127 ( \60470 , \60467 , \60469 );
and \U$60128 ( \60471 , \7729 , RI98702b8_82);
and \U$60129 ( \60472 , RI9870768_92, \7727 );
nor \U$60130 ( \60473 , \60471 , \60472 );
and \U$60131 ( \60474 , \60473 , \7480 );
not \U$60132 ( \60475 , \60473 );
and \U$60133 ( \60476 , \60475 , \7733 );
nor \U$60134 ( \60477 , \60474 , \60476 );
xor \U$60135 ( \60478 , \60470 , \60477 );
and \U$60136 ( \60479 , \8486 , RI9870678_90);
and \U$60137 ( \60480 , RI9870948_96, \8484 );
nor \U$60138 ( \60481 , \60479 , \60480 );
and \U$60139 ( \60482 , \60481 , \8050 );
not \U$60140 ( \60483 , \60481 );
and \U$60141 ( \60484 , \60483 , \8051 );
nor \U$60142 ( \60485 , \60482 , \60484 );
and \U$60143 ( \60486 , \60478 , \60485 );
and \U$60144 ( \60487 , \60470 , \60477 );
or \U$60145 ( \60488 , \60486 , \60487 );
nand \U$60146 ( \60489 , RI9870498_86, \6451 );
and \U$60147 ( \60490 , \60489 , \6190 );
not \U$60148 ( \60491 , \60489 );
and \U$60149 ( \60492 , \60491 , \6705 );
nor \U$60150 ( \60493 , \60490 , \60492 );
and \U$60151 ( \60494 , \7079 , RI9870588_88);
and \U$60152 ( \60495 , RI98703a8_84, \7077 );
nor \U$60153 ( \60496 , \60494 , \60495 );
and \U$60154 ( \60497 , \60496 , \6710 );
not \U$60155 ( \60498 , \60496 );
and \U$60156 ( \60499 , \60498 , \6709 );
nor \U$60157 ( \60500 , \60497 , \60499 );
and \U$60158 ( \60501 , \60493 , \60500 );
xnor \U$60159 ( \60502 , \60488 , \60501 );
not \U$60160 ( \60503 , \60502 );
and \U$60161 ( \60504 , \6453 , RI9870498_86);
and \U$60162 ( \60505 , RI9870588_88, \6451 );
nor \U$60163 ( \60506 , \60504 , \60505 );
and \U$60164 ( \60507 , \60506 , \6190 );
not \U$60165 ( \60508 , \60506 );
and \U$60166 ( \60509 , \60508 , \6705 );
nor \U$60167 ( \60510 , \60507 , \60509 );
not \U$60168 ( \60511 , \60510 );
and \U$60169 ( \60512 , \60503 , \60511 );
and \U$60170 ( \60513 , \60502 , \60510 );
nor \U$60171 ( \60514 , \60512 , \60513 );
not \U$60172 ( \60515 , \60390 );
not \U$60173 ( \60516 , \60401 );
or \U$60174 ( \60517 , \60515 , \60516 );
or \U$60175 ( \60518 , \60401 , \60390 );
nand \U$60176 ( \60519 , \60517 , \60518 );
not \U$60177 ( \60520 , \60519 );
not \U$60178 ( \60521 , \60382 );
and \U$60179 ( \60522 , \60520 , \60521 );
and \U$60180 ( \60523 , \60519 , \60382 );
nor \U$60181 ( \60524 , \60522 , \60523 );
xor \U$60182 ( \60525 , \60514 , \60524 );
not \U$60183 ( \60526 , \60331 );
not \U$60184 ( \60527 , \60342 );
or \U$60185 ( \60528 , \60526 , \60527 );
or \U$60186 ( \60529 , \60331 , \60342 );
nand \U$60187 ( \60530 , \60528 , \60529 );
not \U$60188 ( \60531 , \60530 );
not \U$60189 ( \60532 , \60324 );
and \U$60190 ( \60533 , \60531 , \60532 );
and \U$60191 ( \60534 , \60530 , \60324 );
nor \U$60192 ( \60535 , \60533 , \60534 );
not \U$60193 ( \60536 , \60535 );
xor \U$60194 ( \60537 , \60357 , \60364 );
xor \U$60195 ( \60538 , \60537 , \60372 );
not \U$60196 ( \60539 , \60538 );
or \U$60197 ( \60540 , \60536 , \60539 );
or \U$60198 ( \60541 , \60535 , \60538 );
nand \U$60199 ( \60542 , \60540 , \60541 );
not \U$60200 ( \60543 , \60542 );
not \U$60201 ( \60544 , \60418 );
not \U$60202 ( \60545 , \60429 );
or \U$60203 ( \60546 , \60544 , \60545 );
or \U$60204 ( \60547 , \60418 , \60429 );
nand \U$60205 ( \60548 , \60546 , \60547 );
not \U$60206 ( \60549 , \60548 );
not \U$60207 ( \60550 , \60411 );
and \U$60208 ( \60551 , \60549 , \60550 );
and \U$60209 ( \60552 , \60548 , \60411 );
nor \U$60210 ( \60553 , \60551 , \60552 );
not \U$60211 ( \60554 , \60553 );
and \U$60212 ( \60555 , \60543 , \60554 );
and \U$60213 ( \60556 , \60542 , \60553 );
nor \U$60214 ( \60557 , \60555 , \60556 );
and \U$60215 ( \60558 , \60525 , \60557 );
and \U$60216 ( \60559 , \60514 , \60524 );
or \U$60217 ( \60560 , \60558 , \60559 );
and \U$60218 ( \60561 , \12293 , RI98701c8_80);
and \U$60219 ( \60562 , RI9870fd8_110, \12291 );
nor \U$60220 ( \60563 , \60561 , \60562 );
and \U$60221 ( \60564 , \60563 , \11687 );
not \U$60222 ( \60565 , \60563 );
and \U$60223 ( \60566 , \60565 , \11686 );
nor \U$60224 ( \60567 , \60564 , \60566 );
and \U$60225 ( \60568 , \13045 , RI9870b28_100);
and \U$60226 ( \60569 , RI9870df8_106, \13043 );
nor \U$60227 ( \60570 , \60568 , \60569 );
and \U$60228 ( \60571 , \60570 , \13047 );
not \U$60229 ( \60572 , \60570 );
and \U$60230 ( \60573 , \60572 , \12619 );
nor \U$60231 ( \60574 , \60571 , \60573 );
xor \U$60232 ( \60575 , \60567 , \60574 );
and \U$60233 ( \60576 , \13882 , RI9870a38_98);
and \U$60234 ( \60577 , RI9870ee8_108, \13880 );
nor \U$60235 ( \60578 , \60576 , \60577 );
and \U$60236 ( \60579 , \60578 , \13358 );
not \U$60237 ( \60580 , \60578 );
and \U$60238 ( \60581 , \60580 , \13359 );
nor \U$60239 ( \60582 , \60579 , \60581 );
xor \U$60240 ( \60583 , \60575 , \60582 );
and \U$60241 ( \60584 , \11696 , RI986fef8_74);
and \U$60242 ( \60585 , RI98700d8_78, \11694 );
nor \U$60243 ( \60586 , \60584 , \60585 );
and \U$60244 ( \60587 , \60586 , \10965 );
not \U$60245 ( \60588 , \60586 );
and \U$60246 ( \60589 , \60588 , \11702 );
nor \U$60247 ( \60590 , \60587 , \60589 );
and \U$60248 ( \60591 , \9505 , RI986fc28_68);
and \U$60249 ( \60592 , RI986fe08_72, \9503 );
nor \U$60250 ( \60593 , \60591 , \60592 );
and \U$60251 ( \60594 , \60593 , \9510 );
not \U$60252 ( \60595 , \60593 );
and \U$60253 ( \60596 , \60595 , \9513 );
nor \U$60254 ( \60597 , \60594 , \60596 );
xor \U$60255 ( \60598 , \60590 , \60597 );
and \U$60256 ( \60599 , \10424 , RI986fd18_70);
and \U$60257 ( \60600 , RI986ffe8_76, \10422 );
nor \U$60258 ( \60601 , \60599 , \60600 );
and \U$60259 ( \60602 , \60601 , \9840 );
not \U$60260 ( \60603 , \60601 );
and \U$60261 ( \60604 , \60603 , \10428 );
nor \U$60262 ( \60605 , \60602 , \60604 );
xor \U$60263 ( \60606 , \60598 , \60605 );
and \U$60264 ( \60607 , \60583 , \60606 );
not \U$60265 ( \60608 , RI9873558_190);
and \U$60266 ( \60609 , \15780 , RI9870d08_104);
and \U$60267 ( \60610 , RI98712a8_116, RI9873648_192);
nor \U$60268 ( \60611 , \60609 , \60610 );
not \U$60269 ( \60612 , \60611 );
or \U$60270 ( \60613 , \60608 , \60612 );
or \U$60271 ( \60614 , \60611 , RI9873558_190);
nand \U$60272 ( \60615 , \60613 , \60614 );
xor \U$60273 ( \60616 , \60615 , \6180 );
and \U$60274 ( \60617 , \14937 , RI9870c18_102);
and \U$60275 ( \60618 , RI98710c8_112, \14935 );
nor \U$60276 ( \60619 , \60617 , \60618 );
and \U$60277 ( \60620 , \60619 , \14539 );
not \U$60278 ( \60621 , \60619 );
and \U$60279 ( \60622 , \60621 , \14538 );
nor \U$60280 ( \60623 , \60620 , \60622 );
xor \U$60281 ( \60624 , \60616 , \60623 );
xor \U$60282 ( \60625 , \60590 , \60597 );
xor \U$60283 ( \60626 , \60625 , \60605 );
and \U$60284 ( \60627 , \60624 , \60626 );
and \U$60285 ( \60628 , \60583 , \60624 );
or \U$60286 ( \60629 , \60607 , \60627 , \60628 );
and \U$60287 ( \60630 , \10424 , RI986fe08_72);
and \U$60288 ( \60631 , RI986fd18_70, \10422 );
nor \U$60289 ( \60632 , \60630 , \60631 );
and \U$60290 ( \60633 , \60632 , \9840 );
not \U$60291 ( \60634 , \60632 );
and \U$60292 ( \60635 , \60634 , \10428 );
nor \U$60293 ( \60636 , \60633 , \60635 );
and \U$60294 ( \60637 , \9237 , RI9870948_96);
and \U$60295 ( \60638 , RI9870858_94, \9235 );
nor \U$60296 ( \60639 , \60637 , \60638 );
and \U$60297 ( \60640 , \60639 , \9241 );
not \U$60298 ( \60641 , \60639 );
and \U$60299 ( \60642 , \60641 , \8836 );
nor \U$60300 ( \60643 , \60640 , \60642 );
xor \U$60301 ( \60644 , \60636 , \60643 );
and \U$60302 ( \60645 , \9505 , RI986fb38_66);
and \U$60303 ( \60646 , RI986fc28_68, \9503 );
nor \U$60304 ( \60647 , \60645 , \60646 );
and \U$60305 ( \60648 , \60647 , \9510 );
not \U$60306 ( \60649 , \60647 );
and \U$60307 ( \60650 , \60649 , \9513 );
nor \U$60308 ( \60651 , \60648 , \60650 );
and \U$60309 ( \60652 , \60644 , \60651 );
and \U$60310 ( \60653 , \60636 , \60643 );
or \U$60311 ( \60654 , \60652 , \60653 );
and \U$60312 ( \60655 , \14937 , RI9870ee8_108);
and \U$60313 ( \60656 , RI9870c18_102, \14935 );
nor \U$60314 ( \60657 , \60655 , \60656 );
and \U$60315 ( \60658 , \60657 , \14539 );
not \U$60316 ( \60659 , \60657 );
and \U$60317 ( \60660 , \60659 , \14538 );
nor \U$60318 ( \60661 , \60658 , \60660 );
not \U$60319 ( \60662 , RI9873558_190);
and \U$60320 ( \60663 , \15780 , RI98710c8_112);
and \U$60321 ( \60664 , RI9870d08_104, RI9873648_192);
nor \U$60322 ( \60665 , \60663 , \60664 );
not \U$60323 ( \60666 , \60665 );
or \U$60324 ( \60667 , \60662 , \60666 );
or \U$60325 ( \60668 , \60665 , RI9873558_190);
nand \U$60326 ( \60669 , \60667 , \60668 );
xor \U$60327 ( \60670 , \60661 , \60669 );
and \U$60328 ( \60671 , \13882 , RI9870df8_106);
and \U$60329 ( \60672 , RI9870a38_98, \13880 );
nor \U$60330 ( \60673 , \60671 , \60672 );
and \U$60331 ( \60674 , \60673 , \13358 );
not \U$60332 ( \60675 , \60673 );
and \U$60333 ( \60676 , \60675 , \13359 );
nor \U$60334 ( \60677 , \60674 , \60676 );
and \U$60335 ( \60678 , \60670 , \60677 );
and \U$60336 ( \60679 , \60661 , \60669 );
or \U$60337 ( \60680 , \60678 , \60679 );
xor \U$60338 ( \60681 , \60654 , \60680 );
and \U$60339 ( \60682 , \13045 , RI9870fd8_110);
and \U$60340 ( \60683 , RI9870b28_100, \13043 );
nor \U$60341 ( \60684 , \60682 , \60683 );
and \U$60342 ( \60685 , \60684 , \13047 );
not \U$60343 ( \60686 , \60684 );
and \U$60344 ( \60687 , \60686 , \12619 );
nor \U$60345 ( \60688 , \60685 , \60687 );
and \U$60346 ( \60689 , \11696 , RI986ffe8_76);
and \U$60347 ( \60690 , RI986fef8_74, \11694 );
nor \U$60348 ( \60691 , \60689 , \60690 );
and \U$60349 ( \60692 , \60691 , \10965 );
not \U$60350 ( \60693 , \60691 );
and \U$60351 ( \60694 , \60693 , \11702 );
nor \U$60352 ( \60695 , \60692 , \60694 );
xor \U$60353 ( \60696 , \60688 , \60695 );
and \U$60354 ( \60697 , \12293 , RI98700d8_78);
and \U$60355 ( \60698 , RI98701c8_80, \12291 );
nor \U$60356 ( \60699 , \60697 , \60698 );
and \U$60357 ( \60700 , \60699 , \11687 );
not \U$60358 ( \60701 , \60699 );
and \U$60359 ( \60702 , \60701 , \11686 );
nor \U$60360 ( \60703 , \60700 , \60702 );
and \U$60361 ( \60704 , \60696 , \60703 );
and \U$60362 ( \60705 , \60688 , \60695 );
or \U$60363 ( \60706 , \60704 , \60705 );
and \U$60364 ( \60707 , \60681 , \60706 );
and \U$60365 ( \60708 , \60654 , \60680 );
or \U$60366 ( \60709 , \60707 , \60708 );
xor \U$60367 ( \60710 , \60629 , \60709 );
and \U$60368 ( \60711 , \7079 , RI9870498_86);
and \U$60369 ( \60712 , RI9870588_88, \7077 );
nor \U$60370 ( \60713 , \60711 , \60712 );
and \U$60371 ( \60714 , \60713 , \6710 );
not \U$60372 ( \60715 , \60713 );
and \U$60373 ( \60716 , \60715 , \6709 );
nor \U$60374 ( \60717 , \60714 , \60716 );
and \U$60375 ( \60718 , \7729 , RI98703a8_84);
and \U$60376 ( \60719 , RI98702b8_82, \7727 );
nor \U$60377 ( \60720 , \60718 , \60719 );
and \U$60378 ( \60721 , \60720 , \7480 );
not \U$60379 ( \60722 , \60720 );
and \U$60380 ( \60723 , \60722 , \7733 );
nor \U$60381 ( \60724 , \60721 , \60723 );
xor \U$60382 ( \60725 , \60717 , \60724 );
and \U$60383 ( \60726 , \8486 , RI9870768_92);
and \U$60384 ( \60727 , RI9870678_90, \8484 );
nor \U$60385 ( \60728 , \60726 , \60727 );
and \U$60386 ( \60729 , \60728 , \8050 );
not \U$60387 ( \60730 , \60728 );
and \U$60388 ( \60731 , \60730 , \8051 );
nor \U$60389 ( \60732 , \60729 , \60731 );
and \U$60390 ( \60733 , \60725 , \60732 );
and \U$60391 ( \60734 , \60717 , \60724 );
or \U$60392 ( \60735 , \60733 , \60734 );
xor \U$60393 ( \60736 , \60493 , \60500 );
xor \U$60394 ( \60737 , \60735 , \60736 );
xor \U$60395 ( \60738 , \60470 , \60477 );
xor \U$60396 ( \60739 , \60738 , \60485 );
and \U$60397 ( \60740 , \60737 , \60739 );
and \U$60398 ( \60741 , \60735 , \60736 );
or \U$60399 ( \60742 , \60740 , \60741 );
and \U$60400 ( \60743 , \60710 , \60742 );
and \U$60401 ( \60744 , \60629 , \60709 );
nor \U$60402 ( \60745 , \60743 , \60744 );
or \U$60403 ( \60746 , \60560 , \60745 );
not \U$60404 ( \60747 , \60745 );
not \U$60405 ( \60748 , \60560 );
or \U$60406 ( \60749 , \60747 , \60748 );
xor \U$60407 ( \60750 , \60317 , \60344 );
xor \U$60408 ( \60751 , \60750 , \60347 );
xor \U$60409 ( \60752 , \60375 , \60403 );
xor \U$60410 ( \60753 , \60752 , \60431 );
xor \U$60411 ( \60754 , \60118 , \60125 );
xor \U$60412 ( \60755 , \60754 , \60133 );
xor \U$60413 ( \60756 , \60437 , \60442 );
xor \U$60414 ( \60757 , \60755 , \60756 );
xor \U$60415 ( \60758 , \60753 , \60757 );
xor \U$60416 ( \60759 , \60751 , \60758 );
nand \U$60417 ( \60760 , \60749 , \60759 );
nand \U$60418 ( \60761 , \60746 , \60760 );
xor \U$60419 ( \60762 , \60567 , \60574 );
and \U$60420 ( \60763 , \60762 , \60582 );
and \U$60421 ( \60764 , \60567 , \60574 );
or \U$60422 ( \60765 , \60763 , \60764 );
xor \U$60423 ( \60766 , \60615 , \6180 );
and \U$60424 ( \60767 , \60766 , \60623 );
and \U$60425 ( \60768 , \60615 , \6180 );
or \U$60426 ( \60769 , \60767 , \60768 );
xor \U$60427 ( \60770 , \60765 , \60769 );
xor \U$60428 ( \60771 , \60590 , \60597 );
and \U$60429 ( \60772 , \60771 , \60605 );
and \U$60430 ( \60773 , \60590 , \60597 );
or \U$60431 ( \60774 , \60772 , \60773 );
and \U$60432 ( \60775 , \60770 , \60774 );
and \U$60433 ( \60776 , \60765 , \60769 );
or \U$60434 ( \60777 , \60775 , \60776 );
not \U$60435 ( \60778 , \60510 );
not \U$60436 ( \60779 , \60501 );
or \U$60437 ( \60780 , \60778 , \60779 );
or \U$60438 ( \60781 , \60501 , \60510 );
nand \U$60439 ( \60782 , \60781 , \60488 );
nand \U$60440 ( \60783 , \60780 , \60782 );
xor \U$60441 ( \60784 , \60777 , \60783 );
or \U$60442 ( \60785 , \60535 , \60553 );
not \U$60443 ( \60786 , \60553 );
not \U$60444 ( \60787 , \60535 );
or \U$60445 ( \60788 , \60786 , \60787 );
nand \U$60446 ( \60789 , \60788 , \60538 );
nand \U$60447 ( \60790 , \60785 , \60789 );
and \U$60448 ( \60791 , \60784 , \60790 );
and \U$60449 ( \60792 , \60777 , \60783 );
or \U$60450 ( \60793 , \60791 , \60792 );
xor \U$60451 ( \60794 , \60162 , \60169 );
xor \U$60452 ( \60795 , \60794 , \60195 );
xor \U$60453 ( \60796 , \60793 , \60795 );
xor \U$60454 ( \60797 , \60317 , \60344 );
xor \U$60455 ( \60798 , \60797 , \60347 );
and \U$60456 ( \60799 , \60753 , \60798 );
xor \U$60457 ( \60800 , \60317 , \60344 );
xor \U$60458 ( \60801 , \60800 , \60347 );
and \U$60459 ( \60802 , \60757 , \60801 );
and \U$60460 ( \60803 , \60753 , \60757 );
or \U$60461 ( \60804 , \60799 , \60802 , \60803 );
xor \U$60462 ( \60805 , \60796 , \60804 );
and \U$60463 ( \60806 , \60761 , \60805 );
xor \U$60464 ( \60807 , \60302 , \60304 );
xor \U$60465 ( \60808 , \60807 , \60309 );
xor \U$60466 ( \60809 , \60091 , \60110 );
xor \U$60467 ( \60810 , \60809 , \60136 );
xor \U$60468 ( \60811 , \60350 , \60434 );
xor \U$60469 ( \60812 , \60811 , \60447 );
xor \U$60470 ( \60813 , \60810 , \60812 );
xor \U$60471 ( \60814 , \60808 , \60813 );
xor \U$60472 ( \60815 , \60793 , \60795 );
xor \U$60473 ( \60816 , \60815 , \60804 );
and \U$60474 ( \60817 , \60814 , \60816 );
and \U$60475 ( \60818 , \60761 , \60814 );
or \U$60476 ( \60819 , \60806 , \60817 , \60818 );
not \U$60477 ( \60820 , \60819 );
xor \U$60478 ( \60821 , \60302 , \60304 );
xor \U$60479 ( \60822 , \60821 , \60309 );
and \U$60480 ( \60823 , \60810 , \60822 );
xor \U$60481 ( \60824 , \60302 , \60304 );
xor \U$60482 ( \60825 , \60824 , \60309 );
and \U$60483 ( \60826 , \60812 , \60825 );
and \U$60484 ( \60827 , \60810 , \60812 );
or \U$60485 ( \60828 , \60823 , \60826 , \60827 );
xor \U$60486 ( \60829 , \60793 , \60795 );
and \U$60487 ( \60830 , \60829 , \60804 );
and \U$60488 ( \60831 , \60793 , \60795 );
or \U$60489 ( \60832 , \60830 , \60831 );
xnor \U$60490 ( \60833 , \60828 , \60832 );
not \U$60491 ( \60834 , \60833 );
xor \U$60492 ( \60835 , \59945 , \59950 );
xor \U$60493 ( \60836 , \60835 , \59953 );
xor \U$60494 ( \60837 , \60224 , \60231 );
xor \U$60495 ( \60838 , \60836 , \60837 );
not \U$60496 ( \60839 , \60838 );
and \U$60497 ( \60840 , \60834 , \60839 );
and \U$60498 ( \60841 , \60833 , \60838 );
nor \U$60499 ( \60842 , \60840 , \60841 );
not \U$60500 ( \60843 , \60842 );
and \U$60501 ( \60844 , \60820 , \60843 );
and \U$60502 ( \60845 , \60819 , \60842 );
nor \U$60503 ( \60846 , \60844 , \60845 );
not \U$60504 ( \60847 , \60846 );
xor \U$60505 ( \60848 , \60139 , \60198 );
xor \U$60506 ( \60849 , \60848 , \60216 );
xor \U$60507 ( \60850 , \60312 , \60314 );
xor \U$60508 ( \60851 , \60850 , \60450 );
xor \U$60509 ( \60852 , \60849 , \60851 );
not \U$60510 ( \60853 , \60852 );
and \U$60511 ( \60854 , \60847 , \60853 );
and \U$60512 ( \60855 , \60846 , \60852 );
nor \U$60513 ( \60856 , \60854 , \60855 );
xor \U$60514 ( \60857 , \60777 , \60783 );
xor \U$60515 ( \60858 , \60857 , \60790 );
not \U$60516 ( \60859 , \60858 );
xor \U$60517 ( \60860 , \60514 , \60524 );
xor \U$60518 ( \60861 , \60860 , \60557 );
not \U$60519 ( \60862 , \60861 );
xor \U$60520 ( \60863 , \60629 , \60709 );
xor \U$60521 ( \60864 , \60863 , \60742 );
nand \U$60522 ( \60865 , \60862 , \60864 );
nand \U$60523 ( \60866 , \60859 , \60865 );
and \U$60524 ( \60867 , \13045 , RI98701c8_80);
and \U$60525 ( \60868 , RI9870fd8_110, \13043 );
nor \U$60526 ( \60869 , \60867 , \60868 );
and \U$60527 ( \60870 , \60869 , \12619 );
not \U$60528 ( \60871 , \60869 );
and \U$60529 ( \60872 , \60871 , \13047 );
nor \U$60530 ( \60873 , \60870 , \60872 );
and \U$60531 ( \60874 , \13882 , RI9870b28_100);
and \U$60532 ( \60875 , RI9870df8_106, \13880 );
nor \U$60533 ( \60876 , \60874 , \60875 );
and \U$60534 ( \60877 , \60876 , \13359 );
not \U$60535 ( \60878 , \60876 );
and \U$60536 ( \60879 , \60878 , \13358 );
nor \U$60537 ( \60880 , \60877 , \60879 );
xor \U$60538 ( \60881 , \60873 , \60880 );
and \U$60539 ( \60882 , \12293 , RI986fef8_74);
and \U$60540 ( \60883 , RI98700d8_78, \12291 );
nor \U$60541 ( \60884 , \60882 , \60883 );
and \U$60542 ( \60885 , \60884 , \11686 );
not \U$60543 ( \60886 , \60884 );
and \U$60544 ( \60887 , \60886 , \11687 );
nor \U$60545 ( \60888 , \60885 , \60887 );
and \U$60546 ( \60889 , \60881 , \60888 );
and \U$60547 ( \60890 , \60873 , \60880 );
nor \U$60548 ( \60891 , \60889 , \60890 );
not \U$60549 ( \60892 , RI9873558_190);
and \U$60550 ( \60893 , \15780 , RI9870c18_102);
and \U$60551 ( \60894 , RI98710c8_112, RI9873648_192);
nor \U$60552 ( \60895 , \60893 , \60894 );
not \U$60553 ( \60896 , \60895 );
or \U$60554 ( \60897 , \60892 , \60896 );
or \U$60555 ( \60898 , \60895 , RI9873558_190);
nand \U$60556 ( \60899 , \60897 , \60898 );
xor \U$60557 ( \60900 , \60899 , \6709 );
and \U$60558 ( \60901 , \14937 , RI9870a38_98);
and \U$60559 ( \60902 , RI9870ee8_108, \14935 );
nor \U$60560 ( \60903 , \60901 , \60902 );
and \U$60561 ( \60904 , \60903 , \14539 );
not \U$60562 ( \60905 , \60903 );
and \U$60563 ( \60906 , \60905 , \14538 );
nor \U$60564 ( \60907 , \60904 , \60906 );
and \U$60565 ( \60908 , \60900 , \60907 );
and \U$60566 ( \60909 , \60899 , \6709 );
or \U$60567 ( \60910 , \60908 , \60909 );
xor \U$60568 ( \60911 , \60891 , \60910 );
and \U$60569 ( \60912 , \11696 , RI986fd18_70);
and \U$60570 ( \60913 , RI986ffe8_76, \11694 );
nor \U$60571 ( \60914 , \60912 , \60913 );
and \U$60572 ( \60915 , \60914 , \10965 );
not \U$60573 ( \60916 , \60914 );
and \U$60574 ( \60917 , \60916 , \11702 );
nor \U$60575 ( \60918 , \60915 , \60917 );
and \U$60576 ( \60919 , \9505 , RI9870858_94);
and \U$60577 ( \60920 , RI986fb38_66, \9503 );
nor \U$60578 ( \60921 , \60919 , \60920 );
and \U$60579 ( \60922 , \60921 , \9510 );
not \U$60580 ( \60923 , \60921 );
and \U$60581 ( \60924 , \60923 , \9513 );
nor \U$60582 ( \60925 , \60922 , \60924 );
xor \U$60583 ( \60926 , \60918 , \60925 );
and \U$60584 ( \60927 , \10424 , RI986fc28_68);
and \U$60585 ( \60928 , RI986fe08_72, \10422 );
nor \U$60586 ( \60929 , \60927 , \60928 );
and \U$60587 ( \60930 , \60929 , \9840 );
not \U$60588 ( \60931 , \60929 );
and \U$60589 ( \60932 , \60931 , \10428 );
nor \U$60590 ( \60933 , \60930 , \60932 );
and \U$60591 ( \60934 , \60926 , \60933 );
and \U$60592 ( \60935 , \60918 , \60925 );
or \U$60593 ( \60936 , \60934 , \60935 );
and \U$60594 ( \60937 , \60911 , \60936 );
and \U$60595 ( \60938 , \60891 , \60910 );
or \U$60596 ( \60939 , \60937 , \60938 );
xor \U$60597 ( \60940 , \60688 , \60695 );
xor \U$60598 ( \60941 , \60940 , \60703 );
xor \U$60599 ( \60942 , \60661 , \60669 );
xor \U$60600 ( \60943 , \60942 , \60677 );
and \U$60601 ( \60944 , \60941 , \60943 );
xor \U$60602 ( \60945 , \60939 , \60944 );
and \U$60603 ( \60946 , \7729 , RI9870588_88);
and \U$60604 ( \60947 , RI98703a8_84, \7727 );
nor \U$60605 ( \60948 , \60946 , \60947 );
and \U$60606 ( \60949 , \60948 , \7480 );
not \U$60607 ( \60950 , \60948 );
and \U$60608 ( \60951 , \60950 , \7733 );
nor \U$60609 ( \60952 , \60949 , \60951 );
and \U$60610 ( \60953 , \8486 , RI98702b8_82);
and \U$60611 ( \60954 , RI9870768_92, \8484 );
nor \U$60612 ( \60955 , \60953 , \60954 );
and \U$60613 ( \60956 , \60955 , \8050 );
not \U$60614 ( \60957 , \60955 );
and \U$60615 ( \60958 , \60957 , \8051 );
nor \U$60616 ( \60959 , \60956 , \60958 );
xor \U$60617 ( \60960 , \60952 , \60959 );
and \U$60618 ( \60961 , \9237 , RI9870678_90);
and \U$60619 ( \60962 , RI9870948_96, \9235 );
nor \U$60620 ( \60963 , \60961 , \60962 );
and \U$60621 ( \60964 , \60963 , \9241 );
not \U$60622 ( \60965 , \60963 );
and \U$60623 ( \60966 , \60965 , \8836 );
nor \U$60624 ( \60967 , \60964 , \60966 );
and \U$60625 ( \60968 , \60960 , \60967 );
and \U$60626 ( \60969 , \60952 , \60959 );
or \U$60627 ( \60970 , \60968 , \60969 );
xor \U$60628 ( \60971 , \60717 , \60724 );
xor \U$60629 ( \60972 , \60971 , \60732 );
and \U$60630 ( \60973 , \60970 , \60972 );
xor \U$60631 ( \60974 , \60636 , \60643 );
xor \U$60632 ( \60975 , \60974 , \60651 );
xor \U$60633 ( \60976 , \60717 , \60724 );
xor \U$60634 ( \60977 , \60976 , \60732 );
and \U$60635 ( \60978 , \60975 , \60977 );
and \U$60636 ( \60979 , \60970 , \60975 );
or \U$60637 ( \60980 , \60973 , \60978 , \60979 );
and \U$60638 ( \60981 , \60945 , \60980 );
and \U$60639 ( \60982 , \60939 , \60944 );
or \U$60640 ( \60983 , \60981 , \60982 );
xor \U$60641 ( \60984 , \60765 , \60769 );
xor \U$60642 ( \60985 , \60984 , \60774 );
xor \U$60643 ( \60986 , \60983 , \60985 );
xor \U$60644 ( \60987 , \60654 , \60680 );
xor \U$60645 ( \60988 , \60987 , \60706 );
xor \U$60646 ( \60989 , \60735 , \60736 );
xor \U$60647 ( \60990 , \60989 , \60739 );
and \U$60648 ( \60991 , \60988 , \60990 );
xor \U$60649 ( \60992 , \60590 , \60597 );
xor \U$60650 ( \60993 , \60992 , \60605 );
xor \U$60651 ( \60994 , \60583 , \60624 );
xor \U$60652 ( \60995 , \60993 , \60994 );
xor \U$60653 ( \60996 , \60735 , \60736 );
xor \U$60654 ( \60997 , \60996 , \60739 );
and \U$60655 ( \60998 , \60995 , \60997 );
and \U$60656 ( \60999 , \60988 , \60995 );
or \U$60657 ( \61000 , \60991 , \60998 , \60999 );
and \U$60658 ( \61001 , \60986 , \61000 );
and \U$60659 ( \61002 , \60983 , \60985 );
or \U$60660 ( \61003 , \61001 , \61002 );
and \U$60661 ( \61004 , \60866 , \61003 );
not \U$60662 ( \61005 , \60865 );
and \U$60663 ( \61006 , \60858 , \61005 );
nor \U$60664 ( \61007 , \61004 , \61006 );
not \U$60665 ( \61008 , \61007 );
xor \U$60666 ( \61009 , \60793 , \60795 );
xor \U$60667 ( \61010 , \61009 , \60804 );
xor \U$60668 ( \61011 , \60761 , \60814 );
xor \U$60669 ( \61012 , \61010 , \61011 );
nand \U$60670 ( \61013 , \61008 , \61012 );
or \U$60671 ( \61014 , \60856 , \61013 );
xnor \U$60672 ( \61015 , \61013 , \60856 );
not \U$60673 ( \61016 , \61007 );
not \U$60674 ( \61017 , \61012 );
or \U$60675 ( \61018 , \61016 , \61017 );
or \U$60676 ( \61019 , \61012 , \61007 );
nand \U$60677 ( \61020 , \61018 , \61019 );
not \U$60678 ( \61021 , \60858 );
not \U$60679 ( \61022 , \61003 );
not \U$60680 ( \61023 , \60865 );
and \U$60681 ( \61024 , \61022 , \61023 );
and \U$60682 ( \61025 , \61003 , \60865 );
nor \U$60683 ( \61026 , \61024 , \61025 );
not \U$60684 ( \61027 , \61026 );
or \U$60685 ( \61028 , \61021 , \61027 );
or \U$60686 ( \61029 , \61026 , \60858 );
nand \U$60687 ( \61030 , \61028 , \61029 );
not \U$60688 ( \61031 , \61030 );
xnor \U$60689 ( \61032 , \60745 , \60560 );
not \U$60690 ( \61033 , \61032 );
not \U$60691 ( \61034 , \60759 );
and \U$60692 ( \61035 , \61033 , \61034 );
and \U$60693 ( \61036 , \61032 , \60759 );
nor \U$60694 ( \61037 , \61035 , \61036 );
nor \U$60695 ( \61038 , \61031 , \61037 );
and \U$60696 ( \61039 , \61020 , \61038 );
xor \U$60697 ( \61040 , \61038 , \61020 );
not \U$60698 ( \61041 , \61030 );
not \U$60699 ( \61042 , \61037 );
and \U$60700 ( \61043 , \61041 , \61042 );
and \U$60701 ( \61044 , \61030 , \61037 );
nor \U$60702 ( \61045 , \61043 , \61044 );
xor \U$60703 ( \61046 , \60983 , \60985 );
xor \U$60704 ( \61047 , \61046 , \61000 );
not \U$60705 ( \61048 , \60861 );
not \U$60706 ( \61049 , \60864 );
or \U$60707 ( \61050 , \61048 , \61049 );
or \U$60708 ( \61051 , \60864 , \60861 );
nand \U$60709 ( \61052 , \61050 , \61051 );
and \U$60710 ( \61053 , \61047 , \61052 );
not \U$60711 ( \61054 , \61047 );
not \U$60712 ( \61055 , \61052 );
and \U$60713 ( \61056 , \61054 , \61055 );
xor \U$60714 ( \61057 , \60941 , \60943 );
xor \U$60715 ( \61058 , \60891 , \60910 );
xor \U$60716 ( \61059 , \61058 , \60936 );
and \U$60717 ( \61060 , \61057 , \61059 );
xor \U$60718 ( \61061 , \60717 , \60724 );
xor \U$60719 ( \61062 , \61061 , \60732 );
xor \U$60720 ( \61063 , \60970 , \60975 );
xor \U$60721 ( \61064 , \61062 , \61063 );
xor \U$60722 ( \61065 , \60891 , \60910 );
xor \U$60723 ( \61066 , \61065 , \60936 );
and \U$60724 ( \61067 , \61064 , \61066 );
and \U$60725 ( \61068 , \61057 , \61064 );
or \U$60726 ( \61069 , \61060 , \61067 , \61068 );
and \U$60727 ( \61070 , \14937 , RI9870df8_106);
and \U$60728 ( \61071 , RI9870a38_98, \14935 );
nor \U$60729 ( \61072 , \61070 , \61071 );
and \U$60730 ( \61073 , \61072 , \14539 );
not \U$60731 ( \61074 , \61072 );
and \U$60732 ( \61075 , \61074 , \14538 );
nor \U$60733 ( \61076 , \61073 , \61075 );
not \U$60734 ( \61077 , RI9873558_190);
and \U$60735 ( \61078 , \15780 , RI9870ee8_108);
and \U$60736 ( \61079 , RI9870c18_102, RI9873648_192);
nor \U$60737 ( \61080 , \61078 , \61079 );
not \U$60738 ( \61081 , \61080 );
or \U$60739 ( \61082 , \61077 , \61081 );
or \U$60740 ( \61083 , \61080 , RI9873558_190);
nand \U$60741 ( \61084 , \61082 , \61083 );
xor \U$60742 ( \61085 , \61076 , \61084 );
and \U$60743 ( \61086 , \13882 , RI9870fd8_110);
and \U$60744 ( \61087 , RI9870b28_100, \13880 );
nor \U$60745 ( \61088 , \61086 , \61087 );
and \U$60746 ( \61089 , \61088 , \13358 );
not \U$60747 ( \61090 , \61088 );
and \U$60748 ( \61091 , \61090 , \13359 );
nor \U$60749 ( \61092 , \61089 , \61091 );
and \U$60750 ( \61093 , \61085 , \61092 );
and \U$60751 ( \61094 , \61076 , \61084 );
nor \U$60752 ( \61095 , \61093 , \61094 );
and \U$60753 ( \61096 , \9505 , RI9870948_96);
and \U$60754 ( \61097 , RI9870858_94, \9503 );
nor \U$60755 ( \61098 , \61096 , \61097 );
and \U$60756 ( \61099 , \61098 , \9513 );
not \U$60757 ( \61100 , \61098 );
and \U$60758 ( \61101 , \61100 , \9510 );
nor \U$60759 ( \61102 , \61099 , \61101 );
and \U$60760 ( \61103 , \9237 , RI9870768_92);
and \U$60761 ( \61104 , RI9870678_90, \9235 );
nor \U$60762 ( \61105 , \61103 , \61104 );
and \U$60763 ( \61106 , \61105 , \8836 );
not \U$60764 ( \61107 , \61105 );
and \U$60765 ( \61108 , \61107 , \9241 );
nor \U$60766 ( \61109 , \61106 , \61108 );
xor \U$60767 ( \61110 , \61102 , \61109 );
and \U$60768 ( \61111 , \10424 , RI986fb38_66);
and \U$60769 ( \61112 , RI986fc28_68, \10422 );
nor \U$60770 ( \61113 , \61111 , \61112 );
and \U$60771 ( \61114 , \61113 , \10428 );
not \U$60772 ( \61115 , \61113 );
and \U$60773 ( \61116 , \61115 , \9840 );
nor \U$60774 ( \61117 , \61114 , \61116 );
and \U$60775 ( \61118 , \61110 , \61117 );
and \U$60776 ( \61119 , \61102 , \61109 );
or \U$60777 ( \61120 , \61118 , \61119 );
xor \U$60778 ( \61121 , \61095 , \61120 );
and \U$60779 ( \61122 , \11696 , RI986fe08_72);
and \U$60780 ( \61123 , RI986fd18_70, \11694 );
nor \U$60781 ( \61124 , \61122 , \61123 );
and \U$60782 ( \61125 , \61124 , \11702 );
not \U$60783 ( \61126 , \61124 );
and \U$60784 ( \61127 , \61126 , \10965 );
nor \U$60785 ( \61128 , \61125 , \61127 );
and \U$60786 ( \61129 , \12293 , RI986ffe8_76);
and \U$60787 ( \61130 , RI986fef8_74, \12291 );
nor \U$60788 ( \61131 , \61129 , \61130 );
and \U$60789 ( \61132 , \61131 , \11686 );
not \U$60790 ( \61133 , \61131 );
and \U$60791 ( \61134 , \61133 , \11687 );
nor \U$60792 ( \61135 , \61132 , \61134 );
xor \U$60793 ( \61136 , \61128 , \61135 );
and \U$60794 ( \61137 , \13045 , RI98700d8_78);
and \U$60795 ( \61138 , RI98701c8_80, \13043 );
nor \U$60796 ( \61139 , \61137 , \61138 );
and \U$60797 ( \61140 , \61139 , \12619 );
not \U$60798 ( \61141 , \61139 );
and \U$60799 ( \61142 , \61141 , \13047 );
nor \U$60800 ( \61143 , \61140 , \61142 );
and \U$60801 ( \61144 , \61136 , \61143 );
and \U$60802 ( \61145 , \61128 , \61135 );
or \U$60803 ( \61146 , \61144 , \61145 );
and \U$60804 ( \61147 , \61121 , \61146 );
and \U$60805 ( \61148 , \61095 , \61120 );
nor \U$60806 ( \61149 , \61147 , \61148 );
xor \U$60807 ( \61150 , \60899 , \6709 );
xor \U$60808 ( \61151 , \61150 , \60907 );
not \U$60809 ( \61152 , \61151 );
xor \U$60810 ( \61153 , \60873 , \60880 );
xor \U$60811 ( \61154 , \61153 , \60888 );
nor \U$60812 ( \61155 , \61152 , \61154 );
xor \U$60813 ( \61156 , \61149 , \61155 );
nand \U$60814 ( \61157 , RI9870498_86, \7077 );
and \U$60815 ( \61158 , \61157 , \6710 );
not \U$60816 ( \61159 , \61157 );
and \U$60817 ( \61160 , \61159 , \6709 );
nor \U$60818 ( \61161 , \61158 , \61160 );
xor \U$60819 ( \61162 , \60918 , \60925 );
xor \U$60820 ( \61163 , \61162 , \60933 );
and \U$60821 ( \61164 , \61161 , \61163 );
xor \U$60822 ( \61165 , \60952 , \60959 );
xor \U$60823 ( \61166 , \61165 , \60967 );
xor \U$60824 ( \61167 , \60918 , \60925 );
xor \U$60825 ( \61168 , \61167 , \60933 );
and \U$60826 ( \61169 , \61166 , \61168 );
and \U$60827 ( \61170 , \61161 , \61166 );
or \U$60828 ( \61171 , \61164 , \61169 , \61170 );
and \U$60829 ( \61172 , \61156 , \61171 );
and \U$60830 ( \61173 , \61149 , \61155 );
or \U$60831 ( \61174 , \61172 , \61173 );
xor \U$60832 ( \61175 , \61069 , \61174 );
xor \U$60833 ( \61176 , \60735 , \60736 );
xor \U$60834 ( \61177 , \61176 , \60739 );
xor \U$60835 ( \61178 , \60988 , \60995 );
xor \U$60836 ( \61179 , \61177 , \61178 );
and \U$60837 ( \61180 , \61175 , \61179 );
and \U$60838 ( \61181 , \61069 , \61174 );
nor \U$60839 ( \61182 , \61180 , \61181 );
nor \U$60840 ( \61183 , \61056 , \61182 );
nor \U$60841 ( \61184 , \61053 , \61183 );
or \U$60842 ( \61185 , \61045 , \61184 );
xnor \U$60843 ( \61186 , \61184 , \61045 );
not \U$60844 ( \61187 , \61182 );
not \U$60845 ( \61188 , \61047 );
or \U$60846 ( \61189 , \61187 , \61188 );
or \U$60847 ( \61190 , \61047 , \61182 );
nand \U$60848 ( \61191 , \61189 , \61190 );
xor \U$60849 ( \61192 , \61052 , \61191 );
xor \U$60850 ( \61193 , \60939 , \60944 );
xor \U$60851 ( \61194 , \61193 , \60980 );
not \U$60852 ( \61195 , \61194 );
xor \U$60853 ( \61196 , \61069 , \61174 );
xor \U$60854 ( \61197 , \61196 , \61179 );
not \U$60855 ( \61198 , \61197 );
or \U$60856 ( \61199 , \61195 , \61198 );
or \U$60857 ( \61200 , \61197 , \61194 );
xor \U$60858 ( \61201 , \61095 , \61120 );
xor \U$60859 ( \61202 , \61201 , \61146 );
not \U$60860 ( \61203 , \61151 );
not \U$60861 ( \61204 , \61154 );
and \U$60862 ( \61205 , \61203 , \61204 );
and \U$60863 ( \61206 , \61151 , \61154 );
nor \U$60864 ( \61207 , \61205 , \61206 );
or \U$60865 ( \61208 , \61202 , \61207 );
not \U$60866 ( \61209 , \61207 );
not \U$60867 ( \61210 , \61202 );
or \U$60868 ( \61211 , \61209 , \61210 );
xor \U$60869 ( \61212 , \60918 , \60925 );
xor \U$60870 ( \61213 , \61212 , \60933 );
xor \U$60871 ( \61214 , \61161 , \61166 );
xor \U$60872 ( \61215 , \61213 , \61214 );
nand \U$60873 ( \61216 , \61211 , \61215 );
nand \U$60874 ( \61217 , \61208 , \61216 );
and \U$60875 ( \61218 , \12293 , RI986fd18_70);
and \U$60876 ( \61219 , RI986ffe8_76, \12291 );
nor \U$60877 ( \61220 , \61218 , \61219 );
and \U$60878 ( \61221 , \61220 , \11687 );
not \U$60879 ( \61222 , \61220 );
and \U$60880 ( \61223 , \61222 , \11686 );
nor \U$60881 ( \61224 , \61221 , \61223 );
and \U$60882 ( \61225 , \13045 , RI986fef8_74);
and \U$60883 ( \61226 , RI98700d8_78, \13043 );
nor \U$60884 ( \61227 , \61225 , \61226 );
and \U$60885 ( \61228 , \61227 , \13047 );
not \U$60886 ( \61229 , \61227 );
and \U$60887 ( \61230 , \61229 , \12619 );
nor \U$60888 ( \61231 , \61228 , \61230 );
xor \U$60889 ( \61232 , \61224 , \61231 );
and \U$60890 ( \61233 , \13882 , RI98701c8_80);
and \U$60891 ( \61234 , RI9870fd8_110, \13880 );
nor \U$60892 ( \61235 , \61233 , \61234 );
and \U$60893 ( \61236 , \61235 , \13358 );
not \U$60894 ( \61237 , \61235 );
and \U$60895 ( \61238 , \61237 , \13359 );
nor \U$60896 ( \61239 , \61236 , \61238 );
and \U$60897 ( \61240 , \61232 , \61239 );
and \U$60898 ( \61241 , \61224 , \61231 );
or \U$60899 ( \61242 , \61240 , \61241 );
not \U$60900 ( \61243 , RI9873558_190);
and \U$60901 ( \61244 , \15780 , RI9870a38_98);
and \U$60902 ( \61245 , RI9870ee8_108, RI9873648_192);
nor \U$60903 ( \61246 , \61244 , \61245 );
not \U$60904 ( \61247 , \61246 );
or \U$60905 ( \61248 , \61243 , \61247 );
or \U$60906 ( \61249 , \61246 , RI9873558_190);
nand \U$60907 ( \61250 , \61248 , \61249 );
xor \U$60908 ( \61251 , \61250 , \7733 );
and \U$60909 ( \61252 , \14937 , RI9870b28_100);
and \U$60910 ( \61253 , RI9870df8_106, \14935 );
nor \U$60911 ( \61254 , \61252 , \61253 );
and \U$60912 ( \61255 , \61254 , \14539 );
not \U$60913 ( \61256 , \61254 );
and \U$60914 ( \61257 , \61256 , \14538 );
nor \U$60915 ( \61258 , \61255 , \61257 );
and \U$60916 ( \61259 , \61251 , \61258 );
and \U$60917 ( \61260 , \61250 , \7733 );
or \U$60918 ( \61261 , \61259 , \61260 );
xor \U$60919 ( \61262 , \61242 , \61261 );
and \U$60920 ( \61263 , \11696 , RI986fc28_68);
and \U$60921 ( \61264 , RI986fe08_72, \11694 );
nor \U$60922 ( \61265 , \61263 , \61264 );
and \U$60923 ( \61266 , \61265 , \10965 );
not \U$60924 ( \61267 , \61265 );
and \U$60925 ( \61268 , \61267 , \11702 );
nor \U$60926 ( \61269 , \61266 , \61268 );
and \U$60927 ( \61270 , \9505 , RI9870678_90);
and \U$60928 ( \61271 , RI9870948_96, \9503 );
nor \U$60929 ( \61272 , \61270 , \61271 );
and \U$60930 ( \61273 , \61272 , \9510 );
not \U$60931 ( \61274 , \61272 );
and \U$60932 ( \61275 , \61274 , \9513 );
nor \U$60933 ( \61276 , \61273 , \61275 );
xor \U$60934 ( \61277 , \61269 , \61276 );
and \U$60935 ( \61278 , \10424 , RI9870858_94);
and \U$60936 ( \61279 , RI986fb38_66, \10422 );
nor \U$60937 ( \61280 , \61278 , \61279 );
and \U$60938 ( \61281 , \61280 , \9840 );
not \U$60939 ( \61282 , \61280 );
and \U$60940 ( \61283 , \61282 , \10428 );
nor \U$60941 ( \61284 , \61281 , \61283 );
and \U$60942 ( \61285 , \61277 , \61284 );
and \U$60943 ( \61286 , \61269 , \61276 );
or \U$60944 ( \61287 , \61285 , \61286 );
and \U$60945 ( \61288 , \61262 , \61287 );
and \U$60946 ( \61289 , \61242 , \61261 );
nor \U$60947 ( \61290 , \61288 , \61289 );
and \U$60948 ( \61291 , \7729 , RI9870498_86);
and \U$60949 ( \61292 , RI9870588_88, \7727 );
nor \U$60950 ( \61293 , \61291 , \61292 );
and \U$60951 ( \61294 , \61293 , \7733 );
not \U$60952 ( \61295 , \61293 );
and \U$60953 ( \61296 , \61295 , \7480 );
nor \U$60954 ( \61297 , \61294 , \61296 );
not \U$60955 ( \61298 , \61297 );
and \U$60956 ( \61299 , \8486 , RI98703a8_84);
and \U$60957 ( \61300 , RI98702b8_82, \8484 );
nor \U$60958 ( \61301 , \61299 , \61300 );
and \U$60959 ( \61302 , \61301 , \8051 );
not \U$60960 ( \61303 , \61301 );
and \U$60961 ( \61304 , \61303 , \8050 );
nor \U$60962 ( \61305 , \61302 , \61304 );
not \U$60963 ( \61306 , \61305 );
and \U$60964 ( \61307 , \61298 , \61306 );
and \U$60965 ( \61308 , \61305 , \61297 );
and \U$60966 ( \61309 , \9237 , RI98702b8_82);
and \U$60967 ( \61310 , RI9870768_92, \9235 );
nor \U$60968 ( \61311 , \61309 , \61310 );
and \U$60969 ( \61312 , \61311 , \9241 );
not \U$60970 ( \61313 , \61311 );
and \U$60971 ( \61314 , \61313 , \8836 );
nor \U$60972 ( \61315 , \61312 , \61314 );
nand \U$60973 ( \61316 , RI9870498_86, \7727 );
and \U$60974 ( \61317 , \61316 , \7480 );
not \U$60975 ( \61318 , \61316 );
and \U$60976 ( \61319 , \61318 , \7733 );
nor \U$60977 ( \61320 , \61317 , \61319 );
xor \U$60978 ( \61321 , \61315 , \61320 );
and \U$60979 ( \61322 , \8486 , RI9870588_88);
and \U$60980 ( \61323 , RI98703a8_84, \8484 );
nor \U$60981 ( \61324 , \61322 , \61323 );
and \U$60982 ( \61325 , \61324 , \8050 );
not \U$60983 ( \61326 , \61324 );
and \U$60984 ( \61327 , \61326 , \8051 );
nor \U$60985 ( \61328 , \61325 , \61327 );
and \U$60986 ( \61329 , \61321 , \61328 );
and \U$60987 ( \61330 , \61315 , \61320 );
or \U$60988 ( \61331 , \61329 , \61330 );
not \U$60989 ( \61332 , \61331 );
nor \U$60990 ( \61333 , \61308 , \61332 );
nor \U$60991 ( \61334 , \61307 , \61333 );
or \U$60992 ( \61335 , \61290 , \61334 );
not \U$60993 ( \61336 , \61334 );
not \U$60994 ( \61337 , \61290 );
or \U$60995 ( \61338 , \61336 , \61337 );
xor \U$60996 ( \61339 , \61102 , \61109 );
xor \U$60997 ( \61340 , \61339 , \61117 );
xor \U$60998 ( \61341 , \61128 , \61135 );
xor \U$60999 ( \61342 , \61341 , \61143 );
or \U$61000 ( \61343 , \61340 , \61342 );
not \U$61001 ( \61344 , \61342 );
not \U$61002 ( \61345 , \61340 );
or \U$61003 ( \61346 , \61344 , \61345 );
xor \U$61004 ( \61347 , \61076 , \61084 );
xor \U$61005 ( \61348 , \61347 , \61092 );
nand \U$61006 ( \61349 , \61346 , \61348 );
nand \U$61007 ( \61350 , \61343 , \61349 );
nand \U$61008 ( \61351 , \61338 , \61350 );
nand \U$61009 ( \61352 , \61335 , \61351 );
xor \U$61010 ( \61353 , \61217 , \61352 );
xor \U$61011 ( \61354 , \60891 , \60910 );
xor \U$61012 ( \61355 , \61354 , \60936 );
xor \U$61013 ( \61356 , \61057 , \61064 );
xor \U$61014 ( \61357 , \61355 , \61356 );
and \U$61015 ( \61358 , \61353 , \61357 );
and \U$61016 ( \61359 , \61217 , \61352 );
or \U$61017 ( \61360 , \61358 , \61359 );
nand \U$61018 ( \61361 , \61200 , \61360 );
nand \U$61019 ( \61362 , \61199 , \61361 );
and \U$61020 ( \61363 , \61192 , \61362 );
xor \U$61021 ( \61364 , \61362 , \61192 );
and \U$61022 ( \61365 , \9237 , RI98703a8_84);
and \U$61023 ( \61366 , RI98702b8_82, \9235 );
nor \U$61024 ( \61367 , \61365 , \61366 );
and \U$61025 ( \61368 , \61367 , \9241 );
not \U$61026 ( \61369 , \61367 );
and \U$61027 ( \61370 , \61369 , \8836 );
nor \U$61028 ( \61371 , \61368 , \61370 );
and \U$61029 ( \61372 , \9505 , RI9870768_92);
and \U$61030 ( \61373 , RI9870678_90, \9503 );
nor \U$61031 ( \61374 , \61372 , \61373 );
and \U$61032 ( \61375 , \61374 , \9510 );
not \U$61033 ( \61376 , \61374 );
and \U$61034 ( \61377 , \61376 , \9513 );
nor \U$61035 ( \61378 , \61375 , \61377 );
xor \U$61036 ( \61379 , \61371 , \61378 );
and \U$61037 ( \61380 , \10424 , RI9870948_96);
and \U$61038 ( \61381 , RI9870858_94, \10422 );
nor \U$61039 ( \61382 , \61380 , \61381 );
and \U$61040 ( \61383 , \61382 , \9840 );
not \U$61041 ( \61384 , \61382 );
and \U$61042 ( \61385 , \61384 , \10428 );
nor \U$61043 ( \61386 , \61383 , \61385 );
and \U$61044 ( \61387 , \61379 , \61386 );
and \U$61045 ( \61388 , \61371 , \61378 );
or \U$61046 ( \61389 , \61387 , \61388 );
and \U$61047 ( \61390 , \14937 , RI9870fd8_110);
and \U$61048 ( \61391 , RI9870b28_100, \14935 );
nor \U$61049 ( \61392 , \61390 , \61391 );
and \U$61050 ( \61393 , \61392 , \14539 );
not \U$61051 ( \61394 , \61392 );
and \U$61052 ( \61395 , \61394 , \14538 );
nor \U$61053 ( \61396 , \61393 , \61395 );
not \U$61054 ( \61397 , RI9873558_190);
and \U$61055 ( \61398 , \15780 , RI9870df8_106);
and \U$61056 ( \61399 , RI9870a38_98, RI9873648_192);
nor \U$61057 ( \61400 , \61398 , \61399 );
not \U$61058 ( \61401 , \61400 );
or \U$61059 ( \61402 , \61397 , \61401 );
or \U$61060 ( \61403 , \61400 , RI9873558_190);
nand \U$61061 ( \61404 , \61402 , \61403 );
xor \U$61062 ( \61405 , \61396 , \61404 );
and \U$61063 ( \61406 , \13882 , RI98700d8_78);
and \U$61064 ( \61407 , RI98701c8_80, \13880 );
nor \U$61065 ( \61408 , \61406 , \61407 );
and \U$61066 ( \61409 , \61408 , \13358 );
not \U$61067 ( \61410 , \61408 );
and \U$61068 ( \61411 , \61410 , \13359 );
nor \U$61069 ( \61412 , \61409 , \61411 );
and \U$61070 ( \61413 , \61405 , \61412 );
and \U$61071 ( \61414 , \61396 , \61404 );
or \U$61072 ( \61415 , \61413 , \61414 );
xor \U$61073 ( \61416 , \61389 , \61415 );
and \U$61074 ( \61417 , \12293 , RI986fe08_72);
and \U$61075 ( \61418 , RI986fd18_70, \12291 );
nor \U$61076 ( \61419 , \61417 , \61418 );
and \U$61077 ( \61420 , \61419 , \11687 );
not \U$61078 ( \61421 , \61419 );
and \U$61079 ( \61422 , \61421 , \11686 );
nor \U$61080 ( \61423 , \61420 , \61422 );
and \U$61081 ( \61424 , \11696 , RI986fb38_66);
and \U$61082 ( \61425 , RI986fc28_68, \11694 );
nor \U$61083 ( \61426 , \61424 , \61425 );
and \U$61084 ( \61427 , \61426 , \10965 );
not \U$61085 ( \61428 , \61426 );
and \U$61086 ( \61429 , \61428 , \11702 );
nor \U$61087 ( \61430 , \61427 , \61429 );
xor \U$61088 ( \61431 , \61423 , \61430 );
and \U$61089 ( \61432 , \13045 , RI986ffe8_76);
and \U$61090 ( \61433 , RI986fef8_74, \13043 );
nor \U$61091 ( \61434 , \61432 , \61433 );
and \U$61092 ( \61435 , \61434 , \13047 );
not \U$61093 ( \61436 , \61434 );
and \U$61094 ( \61437 , \61436 , \12619 );
nor \U$61095 ( \61438 , \61435 , \61437 );
and \U$61096 ( \61439 , \61431 , \61438 );
and \U$61097 ( \61440 , \61423 , \61430 );
or \U$61098 ( \61441 , \61439 , \61440 );
and \U$61099 ( \61442 , \61416 , \61441 );
and \U$61100 ( \61443 , \61389 , \61415 );
nor \U$61101 ( \61444 , \61442 , \61443 );
not \U$61102 ( \61445 , \61444 );
xor \U$61103 ( \61446 , \61315 , \61320 );
xor \U$61104 ( \61447 , \61446 , \61328 );
xor \U$61105 ( \61448 , \61269 , \61276 );
xor \U$61106 ( \61449 , \61448 , \61284 );
and \U$61107 ( \61450 , \61447 , \61449 );
xor \U$61108 ( \61451 , \61224 , \61231 );
xor \U$61109 ( \61452 , \61451 , \61239 );
xor \U$61110 ( \61453 , \61269 , \61276 );
xor \U$61111 ( \61454 , \61453 , \61284 );
and \U$61112 ( \61455 , \61452 , \61454 );
and \U$61113 ( \61456 , \61447 , \61452 );
or \U$61114 ( \61457 , \61450 , \61455 , \61456 );
not \U$61115 ( \61458 , \61457 );
or \U$61116 ( \61459 , \61445 , \61458 );
or \U$61117 ( \61460 , \61457 , \61444 );
nand \U$61118 ( \61461 , \61459 , \61460 );
not \U$61119 ( \61462 , \61461 );
not \U$61120 ( \61463 , \61340 );
not \U$61121 ( \61464 , \61348 );
or \U$61122 ( \61465 , \61463 , \61464 );
or \U$61123 ( \61466 , \61348 , \61340 );
nand \U$61124 ( \61467 , \61465 , \61466 );
not \U$61125 ( \61468 , \61467 );
not \U$61126 ( \61469 , \61342 );
and \U$61127 ( \61470 , \61468 , \61469 );
and \U$61128 ( \61471 , \61467 , \61342 );
nor \U$61129 ( \61472 , \61470 , \61471 );
not \U$61130 ( \61473 , \61472 );
and \U$61131 ( \61474 , \61462 , \61473 );
and \U$61132 ( \61475 , \61461 , \61472 );
nor \U$61133 ( \61476 , \61474 , \61475 );
not \U$61134 ( \61477 , \61476 );
xor \U$61135 ( \61478 , \61242 , \61261 );
xor \U$61136 ( \61479 , \61478 , \61287 );
nand \U$61137 ( \61480 , \61477 , \61479 );
not \U$61138 ( \61481 , \61480 );
xor \U$61139 ( \61482 , \61389 , \61415 );
xor \U$61140 ( \61483 , \61482 , \61441 );
xor \U$61141 ( \61484 , \61269 , \61276 );
xor \U$61142 ( \61485 , \61484 , \61284 );
xor \U$61143 ( \61486 , \61447 , \61452 );
xor \U$61144 ( \61487 , \61485 , \61486 );
and \U$61145 ( \61488 , \61483 , \61487 );
not \U$61146 ( \61489 , \61297 );
not \U$61147 ( \61490 , \61305 );
not \U$61148 ( \61491 , \61331 );
or \U$61149 ( \61492 , \61490 , \61491 );
or \U$61150 ( \61493 , \61331 , \61305 );
nand \U$61151 ( \61494 , \61492 , \61493 );
not \U$61152 ( \61495 , \61494 );
or \U$61153 ( \61496 , \61489 , \61495 );
or \U$61154 ( \61497 , \61494 , \61297 );
nand \U$61155 ( \61498 , \61496 , \61497 );
xor \U$61156 ( \61499 , \61488 , \61498 );
and \U$61157 ( \61500 , \10424 , RI9870678_90);
and \U$61158 ( \61501 , RI9870948_96, \10422 );
nor \U$61159 ( \61502 , \61500 , \61501 );
and \U$61160 ( \61503 , \61502 , \9840 );
not \U$61161 ( \61504 , \61502 );
and \U$61162 ( \61505 , \61504 , \10428 );
nor \U$61163 ( \61506 , \61503 , \61505 );
and \U$61164 ( \61507 , \9505 , RI98702b8_82);
and \U$61165 ( \61508 , RI9870768_92, \9503 );
nor \U$61166 ( \61509 , \61507 , \61508 );
and \U$61167 ( \61510 , \61509 , \9510 );
not \U$61168 ( \61511 , \61509 );
and \U$61169 ( \61512 , \61511 , \9513 );
nor \U$61170 ( \61513 , \61510 , \61512 );
xor \U$61171 ( \61514 , \61506 , \61513 );
and \U$61172 ( \61515 , \11696 , RI9870858_94);
and \U$61173 ( \61516 , RI986fb38_66, \11694 );
nor \U$61174 ( \61517 , \61515 , \61516 );
and \U$61175 ( \61518 , \61517 , \10965 );
not \U$61176 ( \61519 , \61517 );
and \U$61177 ( \61520 , \61519 , \11702 );
nor \U$61178 ( \61521 , \61518 , \61520 );
and \U$61179 ( \61522 , \61514 , \61521 );
and \U$61180 ( \61523 , \61506 , \61513 );
or \U$61181 ( \61524 , \61522 , \61523 );
not \U$61182 ( \61525 , RI9873558_190);
and \U$61183 ( \61526 , \15780 , RI9870b28_100);
and \U$61184 ( \61527 , RI9870df8_106, RI9873648_192);
nor \U$61185 ( \61528 , \61526 , \61527 );
not \U$61186 ( \61529 , \61528 );
or \U$61187 ( \61530 , \61525 , \61529 );
or \U$61188 ( \61531 , \61528 , RI9873558_190);
nand \U$61189 ( \61532 , \61530 , \61531 );
xor \U$61190 ( \61533 , \61532 , \8051 );
and \U$61191 ( \61534 , \14937 , RI98701c8_80);
and \U$61192 ( \61535 , RI9870fd8_110, \14935 );
nor \U$61193 ( \61536 , \61534 , \61535 );
and \U$61194 ( \61537 , \61536 , \14539 );
not \U$61195 ( \61538 , \61536 );
and \U$61196 ( \61539 , \61538 , \14538 );
nor \U$61197 ( \61540 , \61537 , \61539 );
and \U$61198 ( \61541 , \61533 , \61540 );
and \U$61199 ( \61542 , \61532 , \8051 );
or \U$61200 ( \61543 , \61541 , \61542 );
xor \U$61201 ( \61544 , \61524 , \61543 );
and \U$61202 ( \61545 , \13882 , RI986fef8_74);
and \U$61203 ( \61546 , RI98700d8_78, \13880 );
nor \U$61204 ( \61547 , \61545 , \61546 );
and \U$61205 ( \61548 , \61547 , \13358 );
not \U$61206 ( \61549 , \61547 );
and \U$61207 ( \61550 , \61549 , \13359 );
nor \U$61208 ( \61551 , \61548 , \61550 );
and \U$61209 ( \61552 , \12293 , RI986fc28_68);
and \U$61210 ( \61553 , RI986fe08_72, \12291 );
nor \U$61211 ( \61554 , \61552 , \61553 );
and \U$61212 ( \61555 , \61554 , \11687 );
not \U$61213 ( \61556 , \61554 );
and \U$61214 ( \61557 , \61556 , \11686 );
nor \U$61215 ( \61558 , \61555 , \61557 );
xor \U$61216 ( \61559 , \61551 , \61558 );
and \U$61217 ( \61560 , \13045 , RI986fd18_70);
and \U$61218 ( \61561 , RI986ffe8_76, \13043 );
nor \U$61219 ( \61562 , \61560 , \61561 );
and \U$61220 ( \61563 , \61562 , \13047 );
not \U$61221 ( \61564 , \61562 );
and \U$61222 ( \61565 , \61564 , \12619 );
nor \U$61223 ( \61566 , \61563 , \61565 );
and \U$61224 ( \61567 , \61559 , \61566 );
and \U$61225 ( \61568 , \61551 , \61558 );
or \U$61226 ( \61569 , \61567 , \61568 );
and \U$61227 ( \61570 , \61544 , \61569 );
and \U$61228 ( \61571 , \61524 , \61543 );
or \U$61229 ( \61572 , \61570 , \61571 );
xor \U$61230 ( \61573 , \61250 , \7733 );
xor \U$61231 ( \61574 , \61573 , \61258 );
xor \U$61232 ( \61575 , \61572 , \61574 );
and \U$61233 ( \61576 , \8486 , RI9870498_86);
and \U$61234 ( \61577 , RI9870588_88, \8484 );
nor \U$61235 ( \61578 , \61576 , \61577 );
and \U$61236 ( \61579 , \61578 , \8050 );
not \U$61237 ( \61580 , \61578 );
and \U$61238 ( \61581 , \61580 , \8051 );
nor \U$61239 ( \61582 , \61579 , \61581 );
xor \U$61240 ( \61583 , \61371 , \61378 );
xor \U$61241 ( \61584 , \61583 , \61386 );
and \U$61242 ( \61585 , \61582 , \61584 );
xor \U$61243 ( \61586 , \61423 , \61430 );
xor \U$61244 ( \61587 , \61586 , \61438 );
xor \U$61245 ( \61588 , \61371 , \61378 );
xor \U$61246 ( \61589 , \61588 , \61386 );
and \U$61247 ( \61590 , \61587 , \61589 );
and \U$61248 ( \61591 , \61582 , \61587 );
or \U$61249 ( \61592 , \61585 , \61590 , \61591 );
and \U$61250 ( \61593 , \61575 , \61592 );
and \U$61251 ( \61594 , \61572 , \61574 );
or \U$61252 ( \61595 , \61593 , \61594 );
and \U$61253 ( \61596 , \61499 , \61595 );
and \U$61254 ( \61597 , \61488 , \61498 );
or \U$61255 ( \61598 , \61596 , \61597 );
not \U$61256 ( \61599 , \61598 );
or \U$61257 ( \61600 , \61481 , \61599 );
or \U$61258 ( \61601 , \61598 , \61480 );
nand \U$61259 ( \61602 , \61600 , \61601 );
not \U$61260 ( \61603 , \61602 );
xnor \U$61261 ( \61604 , \61334 , \61290 );
not \U$61262 ( \61605 , \61604 );
not \U$61263 ( \61606 , \61350 );
and \U$61264 ( \61607 , \61605 , \61606 );
and \U$61265 ( \61608 , \61604 , \61350 );
nor \U$61266 ( \61609 , \61607 , \61608 );
not \U$61267 ( \61610 , \61609 );
or \U$61268 ( \61611 , \61472 , \61444 );
not \U$61269 ( \61612 , \61444 );
not \U$61270 ( \61613 , \61472 );
or \U$61271 ( \61614 , \61612 , \61613 );
nand \U$61272 ( \61615 , \61614 , \61457 );
nand \U$61273 ( \61616 , \61611 , \61615 );
not \U$61274 ( \61617 , \61616 );
or \U$61275 ( \61618 , \61610 , \61617 );
or \U$61276 ( \61619 , \61616 , \61609 );
nand \U$61277 ( \61620 , \61618 , \61619 );
not \U$61278 ( \61621 , \61620 );
not \U$61279 ( \61622 , \61202 );
not \U$61280 ( \61623 , \61215 );
or \U$61281 ( \61624 , \61622 , \61623 );
or \U$61282 ( \61625 , \61215 , \61202 );
nand \U$61283 ( \61626 , \61624 , \61625 );
not \U$61284 ( \61627 , \61626 );
not \U$61285 ( \61628 , \61207 );
and \U$61286 ( \61629 , \61627 , \61628 );
and \U$61287 ( \61630 , \61626 , \61207 );
nor \U$61288 ( \61631 , \61629 , \61630 );
not \U$61289 ( \61632 , \61631 );
and \U$61290 ( \61633 , \61621 , \61632 );
and \U$61291 ( \61634 , \61620 , \61631 );
nor \U$61292 ( \61635 , \61633 , \61634 );
not \U$61293 ( \61636 , \61635 );
and \U$61294 ( \61637 , \61603 , \61636 );
and \U$61295 ( \61638 , \61602 , \61635 );
nor \U$61296 ( \61639 , \61637 , \61638 );
not \U$61297 ( \61640 , \61479 );
not \U$61298 ( \61641 , \61476 );
or \U$61299 ( \61642 , \61640 , \61641 );
or \U$61300 ( \61643 , \61476 , \61479 );
nand \U$61301 ( \61644 , \61642 , \61643 );
xor \U$61302 ( \61645 , \61483 , \61487 );
and \U$61303 ( \61646 , \9237 , RI9870588_88);
and \U$61304 ( \61647 , RI98703a8_84, \9235 );
nor \U$61305 ( \61648 , \61646 , \61647 );
and \U$61306 ( \61649 , \61648 , \9241 );
not \U$61307 ( \61650 , \61648 );
and \U$61308 ( \61651 , \61650 , \8836 );
nor \U$61309 ( \61652 , \61649 , \61651 );
nand \U$61310 ( \61653 , RI9870498_86, \8484 );
and \U$61311 ( \61654 , \61653 , \8050 );
not \U$61312 ( \61655 , \61653 );
and \U$61313 ( \61656 , \61655 , \8051 );
nor \U$61314 ( \61657 , \61654 , \61656 );
xor \U$61315 ( \61658 , \61652 , \61657 );
xor \U$61316 ( \61659 , \61506 , \61513 );
xor \U$61317 ( \61660 , \61659 , \61521 );
and \U$61318 ( \61661 , \61658 , \61660 );
and \U$61319 ( \61662 , \61652 , \61657 );
or \U$61320 ( \61663 , \61661 , \61662 );
xor \U$61321 ( \61664 , \61396 , \61404 );
xor \U$61322 ( \61665 , \61664 , \61412 );
xor \U$61323 ( \61666 , \61663 , \61665 );
and \U$61324 ( \61667 , \13045 , RI986fe08_72);
and \U$61325 ( \61668 , RI986fd18_70, \13043 );
nor \U$61326 ( \61669 , \61667 , \61668 );
and \U$61327 ( \61670 , \61669 , \13047 );
not \U$61328 ( \61671 , \61669 );
and \U$61329 ( \61672 , \61671 , \12619 );
nor \U$61330 ( \61673 , \61670 , \61672 );
and \U$61331 ( \61674 , \11696 , RI9870948_96);
and \U$61332 ( \61675 , RI9870858_94, \11694 );
nor \U$61333 ( \61676 , \61674 , \61675 );
and \U$61334 ( \61677 , \61676 , \10965 );
not \U$61335 ( \61678 , \61676 );
and \U$61336 ( \61679 , \61678 , \11702 );
nor \U$61337 ( \61680 , \61677 , \61679 );
xor \U$61338 ( \61681 , \61673 , \61680 );
and \U$61339 ( \61682 , \12293 , RI986fb38_66);
and \U$61340 ( \61683 , RI986fc28_68, \12291 );
nor \U$61341 ( \61684 , \61682 , \61683 );
and \U$61342 ( \61685 , \61684 , \11687 );
not \U$61343 ( \61686 , \61684 );
and \U$61344 ( \61687 , \61686 , \11686 );
nor \U$61345 ( \61688 , \61685 , \61687 );
and \U$61346 ( \61689 , \61681 , \61688 );
and \U$61347 ( \61690 , \61673 , \61680 );
or \U$61348 ( \61691 , \61689 , \61690 );
and \U$61349 ( \61692 , \13882 , RI986ffe8_76);
and \U$61350 ( \61693 , RI986fef8_74, \13880 );
nor \U$61351 ( \61694 , \61692 , \61693 );
and \U$61352 ( \61695 , \61694 , \13359 );
not \U$61353 ( \61696 , \61694 );
and \U$61354 ( \61697 , \61696 , \13358 );
nor \U$61355 ( \61698 , \61695 , \61697 );
and \U$61356 ( \61699 , \15780 , RI9870fd8_110);
and \U$61357 ( \61700 , RI9870b28_100, RI9873648_192);
nor \U$61358 ( \61701 , \61699 , \61700 );
not \U$61359 ( \61702 , \61701 );
not \U$61360 ( \61703 , RI9873558_190);
and \U$61361 ( \61704 , \61702 , \61703 );
and \U$61362 ( \61705 , \61701 , RI9873558_190);
nor \U$61363 ( \61706 , \61704 , \61705 );
or \U$61364 ( \61707 , \61698 , \61706 );
not \U$61365 ( \61708 , \61706 );
not \U$61366 ( \61709 , \61698 );
or \U$61367 ( \61710 , \61708 , \61709 );
and \U$61368 ( \61711 , \14937 , RI98700d8_78);
and \U$61369 ( \61712 , RI98701c8_80, \14935 );
nor \U$61370 ( \61713 , \61711 , \61712 );
and \U$61371 ( \61714 , \61713 , \14539 );
not \U$61372 ( \61715 , \61713 );
and \U$61373 ( \61716 , \61715 , \14538 );
nor \U$61374 ( \61717 , \61714 , \61716 );
nand \U$61375 ( \61718 , \61710 , \61717 );
nand \U$61376 ( \61719 , \61707 , \61718 );
xor \U$61377 ( \61720 , \61691 , \61719 );
and \U$61378 ( \61721 , \9237 , RI9870498_86);
and \U$61379 ( \61722 , RI9870588_88, \9235 );
nor \U$61380 ( \61723 , \61721 , \61722 );
and \U$61381 ( \61724 , \61723 , \8836 );
not \U$61382 ( \61725 , \61723 );
and \U$61383 ( \61726 , \61725 , \9241 );
nor \U$61384 ( \61727 , \61724 , \61726 );
and \U$61385 ( \61728 , \9505 , RI98703a8_84);
and \U$61386 ( \61729 , RI98702b8_82, \9503 );
nor \U$61387 ( \61730 , \61728 , \61729 );
and \U$61388 ( \61731 , \61730 , \9513 );
not \U$61389 ( \61732 , \61730 );
and \U$61390 ( \61733 , \61732 , \9510 );
nor \U$61391 ( \61734 , \61731 , \61733 );
or \U$61392 ( \61735 , \61727 , \61734 );
not \U$61393 ( \61736 , \61734 );
not \U$61394 ( \61737 , \61727 );
or \U$61395 ( \61738 , \61736 , \61737 );
and \U$61396 ( \61739 , \10424 , RI9870768_92);
and \U$61397 ( \61740 , RI9870678_90, \10422 );
nor \U$61398 ( \61741 , \61739 , \61740 );
and \U$61399 ( \61742 , \61741 , \9840 );
not \U$61400 ( \61743 , \61741 );
and \U$61401 ( \61744 , \61743 , \10428 );
nor \U$61402 ( \61745 , \61742 , \61744 );
nand \U$61403 ( \61746 , \61738 , \61745 );
nand \U$61404 ( \61747 , \61735 , \61746 );
and \U$61405 ( \61748 , \61720 , \61747 );
and \U$61406 ( \61749 , \61691 , \61719 );
or \U$61407 ( \61750 , \61748 , \61749 );
and \U$61408 ( \61751 , \61666 , \61750 );
and \U$61409 ( \61752 , \61663 , \61665 );
or \U$61410 ( \61753 , \61751 , \61752 );
xor \U$61411 ( \61754 , \61645 , \61753 );
xor \U$61412 ( \61755 , \61572 , \61574 );
xor \U$61413 ( \61756 , \61755 , \61592 );
and \U$61414 ( \61757 , \61754 , \61756 );
and \U$61415 ( \61758 , \61645 , \61753 );
or \U$61416 ( \61759 , \61757 , \61758 );
xor \U$61417 ( \61760 , \61644 , \61759 );
xor \U$61418 ( \61761 , \61488 , \61498 );
xor \U$61419 ( \61762 , \61761 , \61595 );
and \U$61420 ( \61763 , \61760 , \61762 );
and \U$61421 ( \61764 , \61644 , \61759 );
nor \U$61422 ( \61765 , \61763 , \61764 );
or \U$61423 ( \61766 , \61639 , \61765 );
xnor \U$61424 ( \61767 , \61765 , \61639 );
xor \U$61425 ( \61768 , \61524 , \61543 );
xor \U$61426 ( \61769 , \61768 , \61569 );
xor \U$61427 ( \61770 , \61663 , \61665 );
xor \U$61428 ( \61771 , \61770 , \61750 );
xor \U$61429 ( \61772 , \61769 , \61771 );
and \U$61430 ( \61773 , \13045 , RI986fc28_68);
and \U$61431 ( \61774 , RI986fe08_72, \13043 );
nor \U$61432 ( \61775 , \61773 , \61774 );
and \U$61433 ( \61776 , \61775 , \13047 );
not \U$61434 ( \61777 , \61775 );
and \U$61435 ( \61778 , \61777 , \12619 );
nor \U$61436 ( \61779 , \61776 , \61778 );
and \U$61437 ( \61780 , \12293 , RI9870858_94);
and \U$61438 ( \61781 , RI986fb38_66, \12291 );
nor \U$61439 ( \61782 , \61780 , \61781 );
and \U$61440 ( \61783 , \61782 , \11687 );
not \U$61441 ( \61784 , \61782 );
and \U$61442 ( \61785 , \61784 , \11686 );
nor \U$61443 ( \61786 , \61783 , \61785 );
xor \U$61444 ( \61787 , \61779 , \61786 );
and \U$61445 ( \61788 , \13882 , RI986fd18_70);
and \U$61446 ( \61789 , RI986ffe8_76, \13880 );
nor \U$61447 ( \61790 , \61788 , \61789 );
and \U$61448 ( \61791 , \61790 , \13358 );
not \U$61449 ( \61792 , \61790 );
and \U$61450 ( \61793 , \61792 , \13359 );
nor \U$61451 ( \61794 , \61791 , \61793 );
and \U$61452 ( \61795 , \61787 , \61794 );
and \U$61453 ( \61796 , \61779 , \61786 );
or \U$61454 ( \61797 , \61795 , \61796 );
not \U$61455 ( \61798 , RI9873558_190);
and \U$61456 ( \61799 , \15780 , RI98701c8_80);
and \U$61457 ( \61800 , RI9870fd8_110, RI9873648_192);
nor \U$61458 ( \61801 , \61799 , \61800 );
not \U$61459 ( \61802 , \61801 );
or \U$61460 ( \61803 , \61798 , \61802 );
or \U$61461 ( \61804 , \61801 , RI9873558_190);
nand \U$61462 ( \61805 , \61803 , \61804 );
xor \U$61463 ( \61806 , \61805 , \8836 );
and \U$61464 ( \61807 , \14937 , RI986fef8_74);
and \U$61465 ( \61808 , RI98700d8_78, \14935 );
nor \U$61466 ( \61809 , \61807 , \61808 );
and \U$61467 ( \61810 , \61809 , \14539 );
not \U$61468 ( \61811 , \61809 );
and \U$61469 ( \61812 , \61811 , \14538 );
nor \U$61470 ( \61813 , \61810 , \61812 );
and \U$61471 ( \61814 , \61806 , \61813 );
and \U$61472 ( \61815 , \61805 , \8836 );
or \U$61473 ( \61816 , \61814 , \61815 );
xor \U$61474 ( \61817 , \61797 , \61816 );
and \U$61475 ( \61818 , \11696 , RI9870678_90);
and \U$61476 ( \61819 , RI9870948_96, \11694 );
nor \U$61477 ( \61820 , \61818 , \61819 );
and \U$61478 ( \61821 , \61820 , \10965 );
not \U$61479 ( \61822 , \61820 );
and \U$61480 ( \61823 , \61822 , \11702 );
nor \U$61481 ( \61824 , \61821 , \61823 );
and \U$61482 ( \61825 , \9505 , RI9870588_88);
and \U$61483 ( \61826 , RI98703a8_84, \9503 );
nor \U$61484 ( \61827 , \61825 , \61826 );
and \U$61485 ( \61828 , \61827 , \9510 );
not \U$61486 ( \61829 , \61827 );
and \U$61487 ( \61830 , \61829 , \9513 );
nor \U$61488 ( \61831 , \61828 , \61830 );
xor \U$61489 ( \61832 , \61824 , \61831 );
and \U$61490 ( \61833 , \10424 , RI98702b8_82);
and \U$61491 ( \61834 , RI9870768_92, \10422 );
nor \U$61492 ( \61835 , \61833 , \61834 );
and \U$61493 ( \61836 , \61835 , \9840 );
not \U$61494 ( \61837 , \61835 );
and \U$61495 ( \61838 , \61837 , \10428 );
nor \U$61496 ( \61839 , \61836 , \61838 );
and \U$61497 ( \61840 , \61832 , \61839 );
and \U$61498 ( \61841 , \61824 , \61831 );
or \U$61499 ( \61842 , \61840 , \61841 );
and \U$61500 ( \61843 , \61817 , \61842 );
and \U$61501 ( \61844 , \61797 , \61816 );
or \U$61502 ( \61845 , \61843 , \61844 );
xor \U$61503 ( \61846 , \61551 , \61558 );
xor \U$61504 ( \61847 , \61846 , \61566 );
xor \U$61505 ( \61848 , \61845 , \61847 );
not \U$61506 ( \61849 , \61706 );
not \U$61507 ( \61850 , \61717 );
or \U$61508 ( \61851 , \61849 , \61850 );
or \U$61509 ( \61852 , \61717 , \61706 );
nand \U$61510 ( \61853 , \61851 , \61852 );
not \U$61511 ( \61854 , \61853 );
not \U$61512 ( \61855 , \61698 );
and \U$61513 ( \61856 , \61854 , \61855 );
and \U$61514 ( \61857 , \61853 , \61698 );
nor \U$61515 ( \61858 , \61856 , \61857 );
not \U$61516 ( \61859 , \61734 );
not \U$61517 ( \61860 , \61745 );
or \U$61518 ( \61861 , \61859 , \61860 );
or \U$61519 ( \61862 , \61734 , \61745 );
nand \U$61520 ( \61863 , \61861 , \61862 );
not \U$61521 ( \61864 , \61863 );
not \U$61522 ( \61865 , \61727 );
and \U$61523 ( \61866 , \61864 , \61865 );
and \U$61524 ( \61867 , \61863 , \61727 );
nor \U$61525 ( \61868 , \61866 , \61867 );
or \U$61526 ( \61869 , \61858 , \61868 );
not \U$61527 ( \61870 , \61868 );
not \U$61528 ( \61871 , \61858 );
or \U$61529 ( \61872 , \61870 , \61871 );
xor \U$61530 ( \61873 , \61673 , \61680 );
xor \U$61531 ( \61874 , \61873 , \61688 );
nand \U$61532 ( \61875 , \61872 , \61874 );
nand \U$61533 ( \61876 , \61869 , \61875 );
and \U$61534 ( \61877 , \61848 , \61876 );
and \U$61535 ( \61878 , \61845 , \61847 );
or \U$61536 ( \61879 , \61877 , \61878 );
xor \U$61537 ( \61880 , \61371 , \61378 );
xor \U$61538 ( \61881 , \61880 , \61386 );
xor \U$61539 ( \61882 , \61582 , \61587 );
xor \U$61540 ( \61883 , \61881 , \61882 );
xor \U$61541 ( \61884 , \61879 , \61883 );
xor \U$61542 ( \61885 , \61532 , \8051 );
xor \U$61543 ( \61886 , \61885 , \61540 );
xor \U$61544 ( \61887 , \61652 , \61657 );
xor \U$61545 ( \61888 , \61887 , \61660 );
and \U$61546 ( \61889 , \61886 , \61888 );
xor \U$61547 ( \61890 , \61691 , \61719 );
xor \U$61548 ( \61891 , \61890 , \61747 );
xor \U$61549 ( \61892 , \61652 , \61657 );
xor \U$61550 ( \61893 , \61892 , \61660 );
and \U$61551 ( \61894 , \61891 , \61893 );
and \U$61552 ( \61895 , \61886 , \61891 );
or \U$61553 ( \61896 , \61889 , \61894 , \61895 );
xor \U$61554 ( \61897 , \61884 , \61896 );
xor \U$61555 ( \61898 , \61772 , \61897 );
xor \U$61556 ( \61899 , \61845 , \61847 );
xor \U$61557 ( \61900 , \61899 , \61876 );
not \U$61558 ( \61901 , \61900 );
xor \U$61559 ( \61902 , \61652 , \61657 );
xor \U$61560 ( \61903 , \61902 , \61660 );
xor \U$61561 ( \61904 , \61886 , \61891 );
xor \U$61562 ( \61905 , \61903 , \61904 );
not \U$61563 ( \61906 , \61905 );
or \U$61564 ( \61907 , \61901 , \61906 );
or \U$61565 ( \61908 , \61905 , \61900 );
not \U$61566 ( \61909 , \61874 );
not \U$61567 ( \61910 , \61858 );
or \U$61568 ( \61911 , \61909 , \61910 );
or \U$61569 ( \61912 , \61858 , \61874 );
nand \U$61570 ( \61913 , \61911 , \61912 );
not \U$61571 ( \61914 , \61913 );
not \U$61572 ( \61915 , \61868 );
and \U$61573 ( \61916 , \61914 , \61915 );
and \U$61574 ( \61917 , \61913 , \61868 );
nor \U$61575 ( \61918 , \61916 , \61917 );
nand \U$61576 ( \61919 , RI9870498_86, \9235 );
and \U$61577 ( \61920 , \61919 , \9241 );
not \U$61578 ( \61921 , \61919 );
and \U$61579 ( \61922 , \61921 , \8836 );
nor \U$61580 ( \61923 , \61920 , \61922 );
xor \U$61581 ( \61924 , \61779 , \61786 );
xor \U$61582 ( \61925 , \61924 , \61794 );
and \U$61583 ( \61926 , \61923 , \61925 );
xor \U$61584 ( \61927 , \61824 , \61831 );
xor \U$61585 ( \61928 , \61927 , \61839 );
xor \U$61586 ( \61929 , \61779 , \61786 );
xor \U$61587 ( \61930 , \61929 , \61794 );
and \U$61588 ( \61931 , \61928 , \61930 );
and \U$61589 ( \61932 , \61923 , \61928 );
or \U$61590 ( \61933 , \61926 , \61931 , \61932 );
not \U$61591 ( \61934 , \61933 );
or \U$61592 ( \61935 , \61918 , \61934 );
not \U$61593 ( \61936 , \61934 );
not \U$61594 ( \61937 , \61918 );
or \U$61595 ( \61938 , \61936 , \61937 );
and \U$61596 ( \61939 , \14937 , RI986ffe8_76);
and \U$61597 ( \61940 , RI986fef8_74, \14935 );
nor \U$61598 ( \61941 , \61939 , \61940 );
and \U$61599 ( \61942 , \61941 , \14539 );
not \U$61600 ( \61943 , \61941 );
and \U$61601 ( \61944 , \61943 , \14538 );
nor \U$61602 ( \61945 , \61942 , \61944 );
not \U$61603 ( \61946 , RI9873558_190);
and \U$61604 ( \61947 , \15780 , RI98700d8_78);
and \U$61605 ( \61948 , RI98701c8_80, RI9873648_192);
nor \U$61606 ( \61949 , \61947 , \61948 );
not \U$61607 ( \61950 , \61949 );
or \U$61608 ( \61951 , \61946 , \61950 );
or \U$61609 ( \61952 , \61949 , RI9873558_190);
nand \U$61610 ( \61953 , \61951 , \61952 );
xor \U$61611 ( \61954 , \61945 , \61953 );
and \U$61612 ( \61955 , \13882 , RI986fe08_72);
and \U$61613 ( \61956 , RI986fd18_70, \13880 );
nor \U$61614 ( \61957 , \61955 , \61956 );
and \U$61615 ( \61958 , \61957 , \13358 );
not \U$61616 ( \61959 , \61957 );
and \U$61617 ( \61960 , \61959 , \13359 );
nor \U$61618 ( \61961 , \61958 , \61960 );
and \U$61619 ( \61962 , \61954 , \61961 );
and \U$61620 ( \61963 , \61945 , \61953 );
or \U$61621 ( \61964 , \61962 , \61963 );
and \U$61622 ( \61965 , \10424 , RI98703a8_84);
and \U$61623 ( \61966 , RI98702b8_82, \10422 );
nor \U$61624 ( \61967 , \61965 , \61966 );
and \U$61625 ( \61968 , \61967 , \9840 );
not \U$61626 ( \61969 , \61967 );
and \U$61627 ( \61970 , \61969 , \10428 );
nor \U$61628 ( \61971 , \61968 , \61970 );
and \U$61629 ( \61972 , \9505 , RI9870498_86);
and \U$61630 ( \61973 , RI9870588_88, \9503 );
nor \U$61631 ( \61974 , \61972 , \61973 );
and \U$61632 ( \61975 , \61974 , \9510 );
not \U$61633 ( \61976 , \61974 );
and \U$61634 ( \61977 , \61976 , \9513 );
nor \U$61635 ( \61978 , \61975 , \61977 );
and \U$61636 ( \61979 , \61971 , \61978 );
xor \U$61637 ( \61980 , \61964 , \61979 );
and \U$61638 ( \61981 , \11696 , RI9870768_92);
and \U$61639 ( \61982 , RI9870678_90, \11694 );
nor \U$61640 ( \61983 , \61981 , \61982 );
and \U$61641 ( \61984 , \61983 , \10965 );
not \U$61642 ( \61985 , \61983 );
and \U$61643 ( \61986 , \61985 , \11702 );
nor \U$61644 ( \61987 , \61984 , \61986 );
and \U$61645 ( \61988 , \12293 , RI9870948_96);
and \U$61646 ( \61989 , RI9870858_94, \12291 );
nor \U$61647 ( \61990 , \61988 , \61989 );
and \U$61648 ( \61991 , \61990 , \11687 );
not \U$61649 ( \61992 , \61990 );
and \U$61650 ( \61993 , \61992 , \11686 );
nor \U$61651 ( \61994 , \61991 , \61993 );
xor \U$61652 ( \61995 , \61987 , \61994 );
and \U$61653 ( \61996 , \13045 , RI986fb38_66);
and \U$61654 ( \61997 , RI986fc28_68, \13043 );
nor \U$61655 ( \61998 , \61996 , \61997 );
and \U$61656 ( \61999 , \61998 , \13047 );
not \U$61657 ( \62000 , \61998 );
and \U$61658 ( \62001 , \62000 , \12619 );
nor \U$61659 ( \62002 , \61999 , \62001 );
and \U$61660 ( \62003 , \61995 , \62002 );
and \U$61661 ( \62004 , \61987 , \61994 );
or \U$61662 ( \62005 , \62003 , \62004 );
and \U$61663 ( \62006 , \61980 , \62005 );
and \U$61664 ( \62007 , \61964 , \61979 );
or \U$61665 ( \62008 , \62006 , \62007 );
nand \U$61666 ( \62009 , \61938 , \62008 );
nand \U$61667 ( \62010 , \61935 , \62009 );
nand \U$61668 ( \62011 , \61908 , \62010 );
nand \U$61669 ( \62012 , \61907 , \62011 );
xor \U$61670 ( \62013 , \61898 , \62012 );
not \U$61671 ( \62014 , RI9873558_190);
and \U$61672 ( \62015 , \15780 , RI986fef8_74);
and \U$61673 ( \62016 , RI98700d8_78, RI9873648_192);
nor \U$61674 ( \62017 , \62015 , \62016 );
not \U$61675 ( \62018 , \62017 );
or \U$61676 ( \62019 , \62014 , \62018 );
or \U$61677 ( \62020 , \62017 , RI9873558_190);
nand \U$61678 ( \62021 , \62019 , \62020 );
and \U$61679 ( \62022 , \62021 , \9513 );
not \U$61680 ( \62023 , \62021 );
not \U$61681 ( \62024 , \9513 );
and \U$61682 ( \62025 , \62023 , \62024 );
and \U$61683 ( \62026 , \14937 , RI986fd18_70);
and \U$61684 ( \62027 , RI986ffe8_76, \14935 );
nor \U$61685 ( \62028 , \62026 , \62027 );
and \U$61686 ( \62029 , \62028 , \14538 );
not \U$61687 ( \62030 , \62028 );
and \U$61688 ( \62031 , \62030 , \14539 );
nor \U$61689 ( \62032 , \62029 , \62031 );
nor \U$61690 ( \62033 , \62025 , \62032 );
nor \U$61691 ( \62034 , \62022 , \62033 );
and \U$61692 ( \62035 , \10424 , RI9870588_88);
and \U$61693 ( \62036 , RI98703a8_84, \10422 );
nor \U$61694 ( \62037 , \62035 , \62036 );
and \U$61695 ( \62038 , \62037 , \10428 );
not \U$61696 ( \62039 , \62037 );
and \U$61697 ( \62040 , \62039 , \9840 );
nor \U$61698 ( \62041 , \62038 , \62040 );
nand \U$61699 ( \62042 , RI9870498_86, \9503 );
and \U$61700 ( \62043 , \62042 , \9513 );
not \U$61701 ( \62044 , \62042 );
and \U$61702 ( \62045 , \62044 , \9510 );
nor \U$61703 ( \62046 , \62043 , \62045 );
xor \U$61704 ( \62047 , \62041 , \62046 );
and \U$61705 ( \62048 , \11696 , RI98702b8_82);
and \U$61706 ( \62049 , RI9870768_92, \11694 );
nor \U$61707 ( \62050 , \62048 , \62049 );
and \U$61708 ( \62051 , \62050 , \11702 );
not \U$61709 ( \62052 , \62050 );
and \U$61710 ( \62053 , \62052 , \10965 );
nor \U$61711 ( \62054 , \62051 , \62053 );
and \U$61712 ( \62055 , \62047 , \62054 );
and \U$61713 ( \62056 , \62041 , \62046 );
or \U$61714 ( \62057 , \62055 , \62056 );
xor \U$61715 ( \62058 , \62034 , \62057 );
and \U$61716 ( \62059 , \13045 , RI9870858_94);
and \U$61717 ( \62060 , RI986fb38_66, \13043 );
nor \U$61718 ( \62061 , \62059 , \62060 );
and \U$61719 ( \62062 , \62061 , \13047 );
not \U$61720 ( \62063 , \62061 );
and \U$61721 ( \62064 , \62063 , \12619 );
nor \U$61722 ( \62065 , \62062 , \62064 );
and \U$61723 ( \62066 , \13882 , RI986fc28_68);
and \U$61724 ( \62067 , RI986fe08_72, \13880 );
nor \U$61725 ( \62068 , \62066 , \62067 );
and \U$61726 ( \62069 , \62068 , \13358 );
not \U$61727 ( \62070 , \62068 );
and \U$61728 ( \62071 , \62070 , \13359 );
nor \U$61729 ( \62072 , \62069 , \62071 );
xor \U$61730 ( \62073 , \62065 , \62072 );
and \U$61731 ( \62074 , \12293 , RI9870678_90);
and \U$61732 ( \62075 , RI9870948_96, \12291 );
nor \U$61733 ( \62076 , \62074 , \62075 );
and \U$61734 ( \62077 , \62076 , \11687 );
not \U$61735 ( \62078 , \62076 );
and \U$61736 ( \62079 , \62078 , \11686 );
nor \U$61737 ( \62080 , \62077 , \62079 );
and \U$61738 ( \62081 , \62073 , \62080 );
and \U$61739 ( \62082 , \62065 , \62072 );
nor \U$61740 ( \62083 , \62081 , \62082 );
and \U$61741 ( \62084 , \62058 , \62083 );
and \U$61742 ( \62085 , \62034 , \62057 );
nor \U$61743 ( \62086 , \62084 , \62085 );
xor \U$61744 ( \62087 , \61805 , \8836 );
xor \U$61745 ( \62088 , \62087 , \61813 );
xor \U$61746 ( \62089 , \62086 , \62088 );
xor \U$61747 ( \62090 , \61971 , \61978 );
xor \U$61748 ( \62091 , \61945 , \61953 );
xor \U$61749 ( \62092 , \62091 , \61961 );
and \U$61750 ( \62093 , \62090 , \62092 );
xor \U$61751 ( \62094 , \61987 , \61994 );
xor \U$61752 ( \62095 , \62094 , \62002 );
xor \U$61753 ( \62096 , \61945 , \61953 );
xor \U$61754 ( \62097 , \62096 , \61961 );
and \U$61755 ( \62098 , \62095 , \62097 );
and \U$61756 ( \62099 , \62090 , \62095 );
or \U$61757 ( \62100 , \62093 , \62098 , \62099 );
and \U$61758 ( \62101 , \62089 , \62100 );
and \U$61759 ( \62102 , \62086 , \62088 );
or \U$61760 ( \62103 , \62101 , \62102 );
xor \U$61761 ( \62104 , \61797 , \61816 );
xor \U$61762 ( \62105 , \62104 , \61842 );
xor \U$61763 ( \62106 , \62103 , \62105 );
xor \U$61764 ( \62107 , \61964 , \61979 );
xor \U$61765 ( \62108 , \62107 , \62005 );
xor \U$61766 ( \62109 , \61779 , \61786 );
xor \U$61767 ( \62110 , \62109 , \61794 );
xor \U$61768 ( \62111 , \61923 , \61928 );
xor \U$61769 ( \62112 , \62110 , \62111 );
and \U$61770 ( \62113 , \62108 , \62112 );
and \U$61771 ( \62114 , \62106 , \62113 );
and \U$61772 ( \62115 , \62103 , \62105 );
or \U$61773 ( \62116 , \62114 , \62115 );
not \U$61774 ( \62117 , \62116 );
xnor \U$61775 ( \62118 , \62010 , \61900 );
not \U$61776 ( \62119 , \62118 );
not \U$61777 ( \62120 , \61905 );
and \U$61778 ( \62121 , \62119 , \62120 );
and \U$61779 ( \62122 , \62118 , \61905 );
nor \U$61780 ( \62123 , \62121 , \62122 );
nor \U$61781 ( \62124 , \62117 , \62123 );
and \U$61782 ( \62125 , \62013 , \62124 );
xor \U$61783 ( \62126 , \62124 , \62013 );
not \U$61784 ( \62127 , \62123 );
not \U$61785 ( \62128 , \62116 );
and \U$61786 ( \62129 , \62127 , \62128 );
and \U$61787 ( \62130 , \62123 , \62116 );
nor \U$61788 ( \62131 , \62129 , \62130 );
not \U$61789 ( \62132 , \62008 );
not \U$61790 ( \62133 , \61934 );
or \U$61791 ( \62134 , \62132 , \62133 );
or \U$61792 ( \62135 , \61934 , \62008 );
nand \U$61793 ( \62136 , \62134 , \62135 );
not \U$61794 ( \62137 , \62136 );
not \U$61795 ( \62138 , \61918 );
and \U$61796 ( \62139 , \62137 , \62138 );
and \U$61797 ( \62140 , \62136 , \61918 );
nor \U$61798 ( \62141 , \62139 , \62140 );
not \U$61799 ( \62142 , \62141 );
xor \U$61800 ( \62143 , \62103 , \62105 );
xor \U$61801 ( \62144 , \62143 , \62113 );
nand \U$61802 ( \62145 , \62142 , \62144 );
or \U$61803 ( \62146 , \62131 , \62145 );
xnor \U$61804 ( \62147 , \62145 , \62131 );
not \U$61805 ( \62148 , \62141 );
not \U$61806 ( \62149 , \62144 );
or \U$61807 ( \62150 , \62148 , \62149 );
or \U$61808 ( \62151 , \62144 , \62141 );
nand \U$61809 ( \62152 , \62150 , \62151 );
xor \U$61810 ( \62153 , \62108 , \62112 );
not \U$61811 ( \62154 , \62153 );
xor \U$61812 ( \62155 , \62086 , \62088 );
xor \U$61813 ( \62156 , \62155 , \62100 );
not \U$61814 ( \62157 , \62156 );
or \U$61815 ( \62158 , \62154 , \62157 );
or \U$61816 ( \62159 , \62156 , \62153 );
xor \U$61817 ( \62160 , \62065 , \62072 );
xor \U$61818 ( \62161 , \62160 , \62080 );
not \U$61819 ( \62162 , \9510 );
not \U$61820 ( \62163 , \62021 );
not \U$61821 ( \62164 , \62032 );
or \U$61822 ( \62165 , \62163 , \62164 );
or \U$61823 ( \62166 , \62032 , \62021 );
nand \U$61824 ( \62167 , \62165 , \62166 );
not \U$61825 ( \62168 , \62167 );
or \U$61826 ( \62169 , \62162 , \62168 );
or \U$61827 ( \62170 , \62167 , \9510 );
nand \U$61828 ( \62171 , \62169 , \62170 );
and \U$61829 ( \62172 , \62161 , \62171 );
not \U$61830 ( \62173 , \62172 );
xor \U$61831 ( \62174 , \61945 , \61953 );
xor \U$61832 ( \62175 , \62174 , \61961 );
xor \U$61833 ( \62176 , \62090 , \62095 );
xor \U$61834 ( \62177 , \62175 , \62176 );
not \U$61835 ( \62178 , \62177 );
or \U$61836 ( \62179 , \62173 , \62178 );
or \U$61837 ( \62180 , \62177 , \62172 );
xor \U$61838 ( \62181 , \62041 , \62046 );
xor \U$61839 ( \62182 , \62181 , \62054 );
and \U$61840 ( \62183 , \13045 , RI9870948_96);
and \U$61841 ( \62184 , RI9870858_94, \13043 );
nor \U$61842 ( \62185 , \62183 , \62184 );
and \U$61843 ( \62186 , \62185 , \13047 );
not \U$61844 ( \62187 , \62185 );
and \U$61845 ( \62188 , \62187 , \12619 );
nor \U$61846 ( \62189 , \62186 , \62188 );
and \U$61847 ( \62190 , \11696 , RI98703a8_84);
and \U$61848 ( \62191 , RI98702b8_82, \11694 );
nor \U$61849 ( \62192 , \62190 , \62191 );
and \U$61850 ( \62193 , \62192 , \10965 );
not \U$61851 ( \62194 , \62192 );
and \U$61852 ( \62195 , \62194 , \11702 );
nor \U$61853 ( \62196 , \62193 , \62195 );
xor \U$61854 ( \62197 , \62189 , \62196 );
and \U$61855 ( \62198 , \12293 , RI9870768_92);
and \U$61856 ( \62199 , RI9870678_90, \12291 );
nor \U$61857 ( \62200 , \62198 , \62199 );
and \U$61858 ( \62201 , \62200 , \11687 );
not \U$61859 ( \62202 , \62200 );
and \U$61860 ( \62203 , \62202 , \11686 );
nor \U$61861 ( \62204 , \62201 , \62203 );
and \U$61862 ( \62205 , \62197 , \62204 );
and \U$61863 ( \62206 , \62189 , \62196 );
or \U$61864 ( \62207 , \62205 , \62206 );
not \U$61865 ( \62208 , \62207 );
or \U$61866 ( \62209 , \62182 , \62208 );
and \U$61867 ( \62210 , \62182 , \62208 );
and \U$61868 ( \62211 , \14937 , RI986fe08_72);
and \U$61869 ( \62212 , RI986fd18_70, \14935 );
nor \U$61870 ( \62213 , \62211 , \62212 );
and \U$61871 ( \62214 , \62213 , \14539 );
not \U$61872 ( \62215 , \62213 );
and \U$61873 ( \62216 , \62215 , \14538 );
nor \U$61874 ( \62217 , \62214 , \62216 );
not \U$61875 ( \62218 , RI9873558_190);
and \U$61876 ( \62219 , \15780 , RI986ffe8_76);
and \U$61877 ( \62220 , RI986fef8_74, RI9873648_192);
nor \U$61878 ( \62221 , \62219 , \62220 );
not \U$61879 ( \62222 , \62221 );
or \U$61880 ( \62223 , \62218 , \62222 );
or \U$61881 ( \62224 , \62221 , RI9873558_190);
nand \U$61882 ( \62225 , \62223 , \62224 );
xor \U$61883 ( \62226 , \62217 , \62225 );
and \U$61884 ( \62227 , \13882 , RI986fb38_66);
and \U$61885 ( \62228 , RI986fc28_68, \13880 );
nor \U$61886 ( \62229 , \62227 , \62228 );
and \U$61887 ( \62230 , \62229 , \13358 );
not \U$61888 ( \62231 , \62229 );
and \U$61889 ( \62232 , \62231 , \13359 );
nor \U$61890 ( \62233 , \62230 , \62232 );
and \U$61891 ( \62234 , \62226 , \62233 );
and \U$61892 ( \62235 , \62217 , \62225 );
nor \U$61893 ( \62236 , \62234 , \62235 );
nor \U$61894 ( \62237 , \62210 , \62236 );
not \U$61895 ( \62238 , \62237 );
nand \U$61896 ( \62239 , \62209 , \62238 );
nand \U$61897 ( \62240 , \62180 , \62239 );
nand \U$61898 ( \62241 , \62179 , \62240 );
nand \U$61899 ( \62242 , \62159 , \62241 );
nand \U$61900 ( \62243 , \62158 , \62242 );
and \U$61901 ( \62244 , \62152 , \62243 );
xor \U$61902 ( \62245 , \62243 , \62152 );
xor \U$61903 ( \62246 , \62217 , \62225 );
xor \U$61904 ( \62247 , \62246 , \62233 );
not \U$61905 ( \62248 , RI9873558_190);
and \U$61906 ( \62249 , \15780 , RI986fd18_70);
and \U$61907 ( \62250 , RI986ffe8_76, RI9873648_192);
nor \U$61908 ( \62251 , \62249 , \62250 );
not \U$61909 ( \62252 , \62251 );
or \U$61910 ( \62253 , \62248 , \62252 );
or \U$61911 ( \62254 , \62251 , RI9873558_190);
nand \U$61912 ( \62255 , \62253 , \62254 );
xor \U$61913 ( \62256 , \62255 , \10428 );
and \U$61914 ( \62257 , \14937 , RI986fc28_68);
and \U$61915 ( \62258 , RI986fe08_72, \14935 );
nor \U$61916 ( \62259 , \62257 , \62258 );
and \U$61917 ( \62260 , \62259 , \14539 );
not \U$61918 ( \62261 , \62259 );
and \U$61919 ( \62262 , \62261 , \14538 );
nor \U$61920 ( \62263 , \62260 , \62262 );
and \U$61921 ( \62264 , \62256 , \62263 );
and \U$61922 ( \62265 , \62255 , \10428 );
or \U$61923 ( \62266 , \62264 , \62265 );
and \U$61924 ( \62267 , \10424 , RI9870498_86);
and \U$61925 ( \62268 , RI9870588_88, \10422 );
nor \U$61926 ( \62269 , \62267 , \62268 );
and \U$61927 ( \62270 , \62269 , \9840 );
not \U$61928 ( \62271 , \62269 );
and \U$61929 ( \62272 , \62271 , \10428 );
nor \U$61930 ( \62273 , \62270 , \62272 );
xor \U$61931 ( \62274 , \62266 , \62273 );
and \U$61932 ( \62275 , \13882 , RI9870858_94);
and \U$61933 ( \62276 , RI986fb38_66, \13880 );
nor \U$61934 ( \62277 , \62275 , \62276 );
and \U$61935 ( \62278 , \62277 , \13358 );
not \U$61936 ( \62279 , \62277 );
and \U$61937 ( \62280 , \62279 , \13359 );
nor \U$61938 ( \62281 , \62278 , \62280 );
and \U$61939 ( \62282 , \12293 , RI98702b8_82);
and \U$61940 ( \62283 , RI9870768_92, \12291 );
nor \U$61941 ( \62284 , \62282 , \62283 );
and \U$61942 ( \62285 , \62284 , \11687 );
not \U$61943 ( \62286 , \62284 );
and \U$61944 ( \62287 , \62286 , \11686 );
nor \U$61945 ( \62288 , \62285 , \62287 );
xor \U$61946 ( \62289 , \62281 , \62288 );
and \U$61947 ( \62290 , \13045 , RI9870678_90);
and \U$61948 ( \62291 , RI9870948_96, \13043 );
nor \U$61949 ( \62292 , \62290 , \62291 );
and \U$61950 ( \62293 , \62292 , \13047 );
not \U$61951 ( \62294 , \62292 );
and \U$61952 ( \62295 , \62294 , \12619 );
nor \U$61953 ( \62296 , \62293 , \62295 );
and \U$61954 ( \62297 , \62289 , \62296 );
and \U$61955 ( \62298 , \62281 , \62288 );
or \U$61956 ( \62299 , \62297 , \62298 );
xor \U$61957 ( \62300 , \62274 , \62299 );
and \U$61958 ( \62301 , \62247 , \62300 );
and \U$61959 ( \62302 , \13882 , RI9870948_96);
and \U$61960 ( \62303 , RI9870858_94, \13880 );
nor \U$61961 ( \62304 , \62302 , \62303 );
and \U$61962 ( \62305 , \62304 , \13359 );
not \U$61963 ( \62306 , \62304 );
and \U$61964 ( \62307 , \62306 , \13358 );
nor \U$61965 ( \62308 , \62305 , \62307 );
and \U$61966 ( \62309 , \15780 , RI986fe08_72);
and \U$61967 ( \62310 , RI986fd18_70, RI9873648_192);
nor \U$61968 ( \62311 , \62309 , \62310 );
not \U$61969 ( \62312 , \62311 );
not \U$61970 ( \62313 , RI9873558_190);
and \U$61971 ( \62314 , \62312 , \62313 );
and \U$61972 ( \62315 , \62311 , RI9873558_190);
nor \U$61973 ( \62316 , \62314 , \62315 );
or \U$61974 ( \62317 , \62308 , \62316 );
not \U$61975 ( \62318 , \62316 );
not \U$61976 ( \62319 , \62308 );
or \U$61977 ( \62320 , \62318 , \62319 );
and \U$61978 ( \62321 , \14937 , RI986fb38_66);
and \U$61979 ( \62322 , RI986fc28_68, \14935 );
nor \U$61980 ( \62323 , \62321 , \62322 );
and \U$61981 ( \62324 , \62323 , \14539 );
not \U$61982 ( \62325 , \62323 );
and \U$61983 ( \62326 , \62325 , \14538 );
nor \U$61984 ( \62327 , \62324 , \62326 );
nand \U$61985 ( \62328 , \62320 , \62327 );
nand \U$61986 ( \62329 , \62317 , \62328 );
and \U$61987 ( \62330 , \11696 , RI9870588_88);
and \U$61988 ( \62331 , RI98703a8_84, \11694 );
nor \U$61989 ( \62332 , \62330 , \62331 );
and \U$61990 ( \62333 , \62332 , \10965 );
not \U$61991 ( \62334 , \62332 );
and \U$61992 ( \62335 , \62334 , \11702 );
nor \U$61993 ( \62336 , \62333 , \62335 );
xor \U$61994 ( \62337 , \62329 , \62336 );
and \U$61995 ( \62338 , \11696 , RI9870498_86);
and \U$61996 ( \62339 , RI9870588_88, \11694 );
nor \U$61997 ( \62340 , \62338 , \62339 );
and \U$61998 ( \62341 , \62340 , \11702 );
not \U$61999 ( \62342 , \62340 );
and \U$62000 ( \62343 , \62342 , \10965 );
nor \U$62001 ( \62344 , \62341 , \62343 );
and \U$62002 ( \62345 , \12293 , RI98703a8_84);
and \U$62003 ( \62346 , RI98702b8_82, \12291 );
nor \U$62004 ( \62347 , \62345 , \62346 );
and \U$62005 ( \62348 , \62347 , \11686 );
not \U$62006 ( \62349 , \62347 );
and \U$62007 ( \62350 , \62349 , \11687 );
nor \U$62008 ( \62351 , \62348 , \62350 );
or \U$62009 ( \62352 , \62344 , \62351 );
not \U$62010 ( \62353 , \62351 );
not \U$62011 ( \62354 , \62344 );
or \U$62012 ( \62355 , \62353 , \62354 );
and \U$62013 ( \62356 , \13045 , RI9870768_92);
and \U$62014 ( \62357 , RI9870678_90, \13043 );
nor \U$62015 ( \62358 , \62356 , \62357 );
and \U$62016 ( \62359 , \62358 , \13047 );
not \U$62017 ( \62360 , \62358 );
and \U$62018 ( \62361 , \62360 , \12619 );
nor \U$62019 ( \62362 , \62359 , \62361 );
nand \U$62020 ( \62363 , \62355 , \62362 );
nand \U$62021 ( \62364 , \62352 , \62363 );
and \U$62022 ( \62365 , \62337 , \62364 );
and \U$62023 ( \62366 , \62329 , \62336 );
or \U$62024 ( \62367 , \62365 , \62366 );
xor \U$62025 ( \62368 , \62189 , \62196 );
xor \U$62026 ( \62369 , \62368 , \62204 );
xor \U$62027 ( \62370 , \62367 , \62369 );
nand \U$62028 ( \62371 , RI9870498_86, \10422 );
and \U$62029 ( \62372 , \62371 , \9840 );
not \U$62030 ( \62373 , \62371 );
and \U$62031 ( \62374 , \62373 , \10428 );
nor \U$62032 ( \62375 , \62372 , \62374 );
xor \U$62033 ( \62376 , \62281 , \62288 );
xor \U$62034 ( \62377 , \62376 , \62296 );
and \U$62035 ( \62378 , \62375 , \62377 );
xor \U$62036 ( \62379 , \62255 , \10428 );
xor \U$62037 ( \62380 , \62379 , \62263 );
xor \U$62038 ( \62381 , \62281 , \62288 );
xor \U$62039 ( \62382 , \62381 , \62296 );
and \U$62040 ( \62383 , \62380 , \62382 );
and \U$62041 ( \62384 , \62375 , \62380 );
or \U$62042 ( \62385 , \62378 , \62383 , \62384 );
and \U$62043 ( \62386 , \62370 , \62385 );
and \U$62044 ( \62387 , \62367 , \62369 );
or \U$62045 ( \62388 , \62386 , \62387 );
xnor \U$62046 ( \62389 , \62301 , \62388 );
not \U$62047 ( \62390 , \62389 );
xor \U$62048 ( \62391 , \62161 , \62171 );
xor \U$62049 ( \62392 , \62266 , \62273 );
and \U$62050 ( \62393 , \62392 , \62299 );
and \U$62051 ( \62394 , \62266 , \62273 );
or \U$62052 ( \62395 , \62393 , \62394 );
not \U$62053 ( \62396 , \62395 );
not \U$62054 ( \62397 , \62207 );
not \U$62055 ( \62398 , \62236 );
or \U$62056 ( \62399 , \62397 , \62398 );
or \U$62057 ( \62400 , \62236 , \62207 );
nand \U$62058 ( \62401 , \62399 , \62400 );
not \U$62059 ( \62402 , \62401 );
not \U$62060 ( \62403 , \62182 );
and \U$62061 ( \62404 , \62402 , \62403 );
and \U$62062 ( \62405 , \62401 , \62182 );
nor \U$62063 ( \62406 , \62404 , \62405 );
not \U$62064 ( \62407 , \62406 );
or \U$62065 ( \62408 , \62396 , \62407 );
or \U$62066 ( \62409 , \62406 , \62395 );
nand \U$62067 ( \62410 , \62408 , \62409 );
xor \U$62068 ( \62411 , \62391 , \62410 );
not \U$62069 ( \62412 , \62411 );
and \U$62070 ( \62413 , \62390 , \62412 );
and \U$62071 ( \62414 , \62389 , \62411 );
nor \U$62072 ( \62415 , \62413 , \62414 );
xor \U$62073 ( \62416 , \62247 , \62300 );
not \U$62074 ( \62417 , \62351 );
not \U$62075 ( \62418 , \62362 );
or \U$62076 ( \62419 , \62417 , \62418 );
or \U$62077 ( \62420 , \62351 , \62362 );
nand \U$62078 ( \62421 , \62419 , \62420 );
not \U$62079 ( \62422 , \62421 );
not \U$62080 ( \62423 , \62344 );
and \U$62081 ( \62424 , \62422 , \62423 );
and \U$62082 ( \62425 , \62421 , \62344 );
nor \U$62083 ( \62426 , \62424 , \62425 );
not \U$62084 ( \62427 , RI9873558_190);
and \U$62085 ( \62428 , \15780 , RI986fc28_68);
and \U$62086 ( \62429 , RI986fe08_72, RI9873648_192);
nor \U$62087 ( \62430 , \62428 , \62429 );
not \U$62088 ( \62431 , \62430 );
or \U$62089 ( \62432 , \62427 , \62431 );
or \U$62090 ( \62433 , \62430 , RI9873558_190);
nand \U$62091 ( \62434 , \62432 , \62433 );
and \U$62092 ( \62435 , \62434 , \11702 );
not \U$62093 ( \62436 , \62434 );
not \U$62094 ( \62437 , \11702 );
and \U$62095 ( \62438 , \62436 , \62437 );
and \U$62096 ( \62439 , \14937 , RI9870858_94);
and \U$62097 ( \62440 , RI986fb38_66, \14935 );
nor \U$62098 ( \62441 , \62439 , \62440 );
and \U$62099 ( \62442 , \62441 , \14538 );
not \U$62100 ( \62443 , \62441 );
and \U$62101 ( \62444 , \62443 , \14539 );
nor \U$62102 ( \62445 , \62442 , \62444 );
nor \U$62103 ( \62446 , \62438 , \62445 );
nor \U$62104 ( \62447 , \62435 , \62446 );
or \U$62105 ( \62448 , \62426 , \62447 );
not \U$62106 ( \62449 , \62447 );
not \U$62107 ( \62450 , \62426 );
or \U$62108 ( \62451 , \62449 , \62450 );
and \U$62109 ( \62452 , \12293 , RI9870588_88);
and \U$62110 ( \62453 , RI98703a8_84, \12291 );
nor \U$62111 ( \62454 , \62452 , \62453 );
and \U$62112 ( \62455 , \62454 , \11686 );
not \U$62113 ( \62456 , \62454 );
and \U$62114 ( \62457 , \62456 , \11687 );
nor \U$62115 ( \62458 , \62455 , \62457 );
and \U$62116 ( \62459 , \13045 , RI98702b8_82);
and \U$62117 ( \62460 , RI9870768_92, \13043 );
nor \U$62118 ( \62461 , \62459 , \62460 );
and \U$62119 ( \62462 , \62461 , \12619 );
not \U$62120 ( \62463 , \62461 );
and \U$62121 ( \62464 , \62463 , \13047 );
nor \U$62122 ( \62465 , \62462 , \62464 );
or \U$62123 ( \62466 , \62458 , \62465 );
not \U$62124 ( \62467 , \62465 );
not \U$62125 ( \62468 , \62458 );
or \U$62126 ( \62469 , \62467 , \62468 );
and \U$62127 ( \62470 , \13882 , RI9870678_90);
and \U$62128 ( \62471 , RI9870948_96, \13880 );
nor \U$62129 ( \62472 , \62470 , \62471 );
and \U$62130 ( \62473 , \62472 , \13358 );
not \U$62131 ( \62474 , \62472 );
and \U$62132 ( \62475 , \62474 , \13359 );
nor \U$62133 ( \62476 , \62473 , \62475 );
nand \U$62134 ( \62477 , \62469 , \62476 );
nand \U$62135 ( \62478 , \62466 , \62477 );
nand \U$62136 ( \62479 , \62451 , \62478 );
nand \U$62137 ( \62480 , \62448 , \62479 );
xor \U$62138 ( \62481 , \62329 , \62336 );
xor \U$62139 ( \62482 , \62481 , \62364 );
and \U$62140 ( \62483 , \62480 , \62482 );
xor \U$62141 ( \62484 , \62281 , \62288 );
xor \U$62142 ( \62485 , \62484 , \62296 );
xor \U$62143 ( \62486 , \62375 , \62380 );
xor \U$62144 ( \62487 , \62485 , \62486 );
xor \U$62145 ( \62488 , \62329 , \62336 );
xor \U$62146 ( \62489 , \62488 , \62364 );
and \U$62147 ( \62490 , \62487 , \62489 );
and \U$62148 ( \62491 , \62480 , \62487 );
or \U$62149 ( \62492 , \62483 , \62490 , \62491 );
xor \U$62150 ( \62493 , \62416 , \62492 );
xor \U$62151 ( \62494 , \62367 , \62369 );
xor \U$62152 ( \62495 , \62494 , \62385 );
and \U$62153 ( \62496 , \62493 , \62495 );
and \U$62154 ( \62497 , \62416 , \62492 );
nor \U$62155 ( \62498 , \62496 , \62497 );
or \U$62156 ( \62499 , \62415 , \62498 );
xnor \U$62157 ( \62500 , \62415 , \62498 );
not \U$62158 ( \62501 , RI9873558_190);
and \U$62159 ( \62502 , \15780 , RI9870858_94);
and \U$62160 ( \62503 , RI986fb38_66, RI9873648_192);
nor \U$62161 ( \62504 , \62502 , \62503 );
not \U$62162 ( \62505 , \62504 );
or \U$62163 ( \62506 , \62501 , \62505 );
or \U$62164 ( \62507 , \62504 , RI9873558_190);
nand \U$62165 ( \62508 , \62506 , \62507 );
xor \U$62166 ( \62509 , \62508 , \11686 );
and \U$62167 ( \62510 , \14937 , RI9870678_90);
and \U$62168 ( \62511 , RI9870948_96, \14935 );
nor \U$62169 ( \62512 , \62510 , \62511 );
and \U$62170 ( \62513 , \62512 , \14539 );
not \U$62171 ( \62514 , \62512 );
and \U$62172 ( \62515 , \62514 , \14538 );
nor \U$62173 ( \62516 , \62513 , \62515 );
and \U$62174 ( \62517 , \62509 , \62516 );
and \U$62175 ( \62518 , \62508 , \11686 );
or \U$62176 ( \62519 , \62517 , \62518 );
and \U$62177 ( \62520 , \13045 , RI98703a8_84);
and \U$62178 ( \62521 , RI98702b8_82, \13043 );
nor \U$62179 ( \62522 , \62520 , \62521 );
and \U$62180 ( \62523 , \62522 , \13047 );
not \U$62181 ( \62524 , \62522 );
and \U$62182 ( \62525 , \62524 , \12619 );
nor \U$62183 ( \62526 , \62523 , \62525 );
xor \U$62184 ( \62527 , \62519 , \62526 );
and \U$62185 ( \62528 , \13045 , RI9870588_88);
and \U$62186 ( \62529 , RI98703a8_84, \13043 );
nor \U$62187 ( \62530 , \62528 , \62529 );
and \U$62188 ( \62531 , \62530 , \13047 );
not \U$62189 ( \62532 , \62530 );
and \U$62190 ( \62533 , \62532 , \12619 );
nor \U$62191 ( \62534 , \62531 , \62533 );
nand \U$62192 ( \62535 , RI9870498_86, \12291 );
and \U$62193 ( \62536 , \62535 , \11687 );
not \U$62194 ( \62537 , \62535 );
and \U$62195 ( \62538 , \62537 , \11686 );
nor \U$62196 ( \62539 , \62536 , \62538 );
xor \U$62197 ( \62540 , \62534 , \62539 );
and \U$62198 ( \62541 , \13882 , RI98702b8_82);
and \U$62199 ( \62542 , RI9870768_92, \13880 );
nor \U$62200 ( \62543 , \62541 , \62542 );
and \U$62201 ( \62544 , \62543 , \13358 );
not \U$62202 ( \62545 , \62543 );
and \U$62203 ( \62546 , \62545 , \13359 );
nor \U$62204 ( \62547 , \62544 , \62546 );
and \U$62205 ( \62548 , \62540 , \62547 );
and \U$62206 ( \62549 , \62534 , \62539 );
or \U$62207 ( \62550 , \62548 , \62549 );
and \U$62208 ( \62551 , \62527 , \62550 );
and \U$62209 ( \62552 , \62519 , \62526 );
or \U$62210 ( \62553 , \62551 , \62552 );
not \U$62211 ( \62554 , \10965 );
not \U$62212 ( \62555 , \62434 );
not \U$62213 ( \62556 , \62445 );
or \U$62214 ( \62557 , \62555 , \62556 );
or \U$62215 ( \62558 , \62445 , \62434 );
nand \U$62216 ( \62559 , \62557 , \62558 );
not \U$62217 ( \62560 , \62559 );
or \U$62218 ( \62561 , \62554 , \62560 );
or \U$62219 ( \62562 , \62559 , \10965 );
nand \U$62220 ( \62563 , \62561 , \62562 );
xor \U$62221 ( \62564 , \62553 , \62563 );
and \U$62222 ( \62565 , \12293 , RI9870498_86);
and \U$62223 ( \62566 , RI9870588_88, \12291 );
nor \U$62224 ( \62567 , \62565 , \62566 );
and \U$62225 ( \62568 , \62567 , \11687 );
not \U$62226 ( \62569 , \62567 );
and \U$62227 ( \62570 , \62569 , \11686 );
nor \U$62228 ( \62571 , \62568 , \62570 );
and \U$62229 ( \62572 , \13882 , RI9870768_92);
and \U$62230 ( \62573 , RI9870678_90, \13880 );
nor \U$62231 ( \62574 , \62572 , \62573 );
and \U$62232 ( \62575 , \62574 , \13359 );
not \U$62233 ( \62576 , \62574 );
and \U$62234 ( \62577 , \62576 , \13358 );
nor \U$62235 ( \62578 , \62575 , \62577 );
not \U$62236 ( \62579 , \62578 );
and \U$62237 ( \62580 , \15780 , RI986fb38_66);
and \U$62238 ( \62581 , RI986fc28_68, RI9873648_192);
nor \U$62239 ( \62582 , \62580 , \62581 );
not \U$62240 ( \62583 , \62582 );
not \U$62241 ( \62584 , RI9873558_190);
and \U$62242 ( \62585 , \62583 , \62584 );
and \U$62243 ( \62586 , \62582 , RI9873558_190);
nor \U$62244 ( \62587 , \62585 , \62586 );
and \U$62245 ( \62588 , \14937 , RI9870948_96);
and \U$62246 ( \62589 , RI9870858_94, \14935 );
nor \U$62247 ( \62590 , \62588 , \62589 );
and \U$62248 ( \62591 , \62590 , \14538 );
not \U$62249 ( \62592 , \62590 );
and \U$62250 ( \62593 , \62592 , \14539 );
nor \U$62251 ( \62594 , \62591 , \62593 );
xor \U$62252 ( \62595 , \62587 , \62594 );
not \U$62253 ( \62596 , \62595 );
or \U$62254 ( \62597 , \62579 , \62596 );
or \U$62255 ( \62598 , \62595 , \62578 );
nand \U$62256 ( \62599 , \62597 , \62598 );
and \U$62257 ( \62600 , \62571 , \62599 );
and \U$62258 ( \62601 , \62564 , \62600 );
and \U$62259 ( \62602 , \62553 , \62563 );
or \U$62260 ( \62603 , \62601 , \62602 );
not \U$62261 ( \62604 , \62603 );
not \U$62262 ( \62605 , \62578 );
not \U$62263 ( \62606 , \62587 );
and \U$62264 ( \62607 , \62605 , \62606 );
and \U$62265 ( \62608 , \62578 , \62587 );
nor \U$62266 ( \62609 , \62608 , \62594 );
nor \U$62267 ( \62610 , \62607 , \62609 );
nand \U$62268 ( \62611 , RI9870498_86, \11694 );
and \U$62269 ( \62612 , \62611 , \11702 );
not \U$62270 ( \62613 , \62611 );
and \U$62271 ( \62614 , \62613 , \10965 );
nor \U$62272 ( \62615 , \62612 , \62614 );
xor \U$62273 ( \62616 , \62610 , \62615 );
not \U$62274 ( \62617 , \62465 );
not \U$62275 ( \62618 , \62476 );
or \U$62276 ( \62619 , \62617 , \62618 );
or \U$62277 ( \62620 , \62465 , \62476 );
nand \U$62278 ( \62621 , \62619 , \62620 );
not \U$62279 ( \62622 , \62621 );
not \U$62280 ( \62623 , \62458 );
and \U$62281 ( \62624 , \62622 , \62623 );
and \U$62282 ( \62625 , \62621 , \62458 );
nor \U$62283 ( \62626 , \62624 , \62625 );
and \U$62284 ( \62627 , \62616 , \62626 );
and \U$62285 ( \62628 , \62610 , \62615 );
or \U$62286 ( \62629 , \62627 , \62628 );
not \U$62287 ( \62630 , \62316 );
not \U$62288 ( \62631 , \62327 );
or \U$62289 ( \62632 , \62630 , \62631 );
or \U$62290 ( \62633 , \62327 , \62316 );
nand \U$62291 ( \62634 , \62632 , \62633 );
not \U$62292 ( \62635 , \62634 );
not \U$62293 ( \62636 , \62308 );
and \U$62294 ( \62637 , \62635 , \62636 );
and \U$62295 ( \62638 , \62634 , \62308 );
nor \U$62296 ( \62639 , \62637 , \62638 );
xor \U$62297 ( \62640 , \62629 , \62639 );
not \U$62298 ( \62641 , \62447 );
not \U$62299 ( \62642 , \62478 );
or \U$62300 ( \62643 , \62641 , \62642 );
or \U$62301 ( \62644 , \62478 , \62447 );
nand \U$62302 ( \62645 , \62643 , \62644 );
not \U$62303 ( \62646 , \62645 );
not \U$62304 ( \62647 , \62426 );
and \U$62305 ( \62648 , \62646 , \62647 );
and \U$62306 ( \62649 , \62645 , \62426 );
nor \U$62307 ( \62650 , \62648 , \62649 );
xor \U$62308 ( \62651 , \62640 , \62650 );
not \U$62309 ( \62652 , \62651 );
or \U$62310 ( \62653 , \62604 , \62652 );
or \U$62311 ( \62654 , \62651 , \62603 );
nand \U$62312 ( \62655 , \62653 , \62654 );
xor \U$62313 ( \62656 , \62553 , \62563 );
xor \U$62314 ( \62657 , \62656 , \62600 );
not \U$62315 ( \62658 , \62657 );
xor \U$62316 ( \62659 , \62610 , \62615 );
xor \U$62317 ( \62660 , \62659 , \62626 );
nor \U$62318 ( \62661 , \62658 , \62660 );
and \U$62319 ( \62662 , \62655 , \62661 );
xor \U$62320 ( \62663 , \62661 , \62655 );
and \U$62321 ( \62664 , \15780 , RI9870948_96);
and \U$62322 ( \62665 , RI9870858_94, RI9873648_192);
nor \U$62323 ( \62666 , \62664 , \62665 );
not \U$62324 ( \62667 , \62666 );
not \U$62325 ( \62668 , RI9873558_190);
and \U$62326 ( \62669 , \62667 , \62668 );
and \U$62327 ( \62670 , \62666 , RI9873558_190);
nor \U$62328 ( \62671 , \62669 , \62670 );
not \U$62329 ( \62672 , \62671 );
and \U$62330 ( \62673 , \14937 , RI9870768_92);
and \U$62331 ( \62674 , RI9870678_90, \14935 );
nor \U$62332 ( \62675 , \62673 , \62674 );
and \U$62333 ( \62676 , \62675 , \14539 );
not \U$62334 ( \62677 , \62675 );
and \U$62335 ( \62678 , \62677 , \14538 );
nor \U$62336 ( \62679 , \62676 , \62678 );
not \U$62337 ( \62680 , \62679 );
or \U$62338 ( \62681 , \62672 , \62680 );
or \U$62339 ( \62682 , \62679 , \62671 );
nand \U$62340 ( \62683 , \62681 , \62682 );
not \U$62341 ( \62684 , \62683 );
and \U$62342 ( \62685 , \13882 , RI98703a8_84);
and \U$62343 ( \62686 , RI98702b8_82, \13880 );
nor \U$62344 ( \62687 , \62685 , \62686 );
and \U$62345 ( \62688 , \62687 , \13359 );
not \U$62346 ( \62689 , \62687 );
and \U$62347 ( \62690 , \62689 , \13358 );
nor \U$62348 ( \62691 , \62688 , \62690 );
not \U$62349 ( \62692 , \62691 );
and \U$62350 ( \62693 , \62684 , \62692 );
and \U$62351 ( \62694 , \62683 , \62691 );
nor \U$62352 ( \62695 , \62693 , \62694 );
not \U$62353 ( \62696 , \62695 );
and \U$62354 ( \62697 , \13045 , RI9870498_86);
and \U$62355 ( \62698 , RI9870588_88, \13043 );
nor \U$62356 ( \62699 , \62697 , \62698 );
and \U$62357 ( \62700 , \62699 , \12619 );
not \U$62358 ( \62701 , \62699 );
and \U$62359 ( \62702 , \62701 , \13047 );
nor \U$62360 ( \62703 , \62700 , \62702 );
not \U$62361 ( \62704 , \62703 );
and \U$62362 ( \62705 , \13882 , RI9870588_88);
and \U$62363 ( \62706 , RI98703a8_84, \13880 );
nor \U$62364 ( \62707 , \62705 , \62706 );
and \U$62365 ( \62708 , \62707 , \13359 );
not \U$62366 ( \62709 , \62707 );
and \U$62367 ( \62710 , \62709 , \13358 );
nor \U$62368 ( \62711 , \62708 , \62710 );
not \U$62369 ( \62712 , \62711 );
nand \U$62370 ( \62713 , RI9870498_86, \13043 );
and \U$62371 ( \62714 , \62713 , \13047 );
not \U$62372 ( \62715 , \62713 );
and \U$62373 ( \62716 , \62715 , \12619 );
nor \U$62374 ( \62717 , \62714 , \62716 );
nand \U$62375 ( \62718 , \62712 , \62717 );
not \U$62376 ( \62719 , \62718 );
not \U$62377 ( \62720 , RI9873558_190);
and \U$62378 ( \62721 , \15780 , RI9870678_90);
and \U$62379 ( \62722 , RI9870948_96, RI9873648_192);
nor \U$62380 ( \62723 , \62721 , \62722 );
not \U$62381 ( \62724 , \62723 );
or \U$62382 ( \62725 , \62720 , \62724 );
or \U$62383 ( \62726 , \62723 , RI9873558_190);
nand \U$62384 ( \62727 , \62725 , \62726 );
xor \U$62385 ( \62728 , \62727 , \12619 );
and \U$62386 ( \62729 , \14937 , RI98702b8_82);
and \U$62387 ( \62730 , RI9870768_92, \14935 );
nor \U$62388 ( \62731 , \62729 , \62730 );
and \U$62389 ( \62732 , \62731 , \14539 );
not \U$62390 ( \62733 , \62731 );
and \U$62391 ( \62734 , \62733 , \14538 );
nor \U$62392 ( \62735 , \62732 , \62734 );
and \U$62393 ( \62736 , \62728 , \62735 );
and \U$62394 ( \62737 , \62727 , \12619 );
or \U$62395 ( \62738 , \62736 , \62737 );
not \U$62396 ( \62739 , \62738 );
or \U$62397 ( \62740 , \62719 , \62739 );
or \U$62398 ( \62741 , \62738 , \62718 );
nand \U$62399 ( \62742 , \62740 , \62741 );
not \U$62400 ( \62743 , \62742 );
or \U$62401 ( \62744 , \62704 , \62743 );
or \U$62402 ( \62745 , \62742 , \62703 );
nand \U$62403 ( \62746 , \62744 , \62745 );
nand \U$62404 ( \62747 , \62696 , \62746 );
xor \U$62405 ( \62748 , \62508 , \11686 );
xor \U$62406 ( \62749 , \62748 , \62516 );
or \U$62407 ( \62750 , \62691 , \62671 );
not \U$62408 ( \62751 , \62671 );
not \U$62409 ( \62752 , \62691 );
or \U$62410 ( \62753 , \62751 , \62752 );
nand \U$62411 ( \62754 , \62753 , \62679 );
nand \U$62412 ( \62755 , \62750 , \62754 );
xor \U$62413 ( \62756 , \62534 , \62539 );
xor \U$62414 ( \62757 , \62756 , \62547 );
xor \U$62415 ( \62758 , \62755 , \62757 );
xor \U$62416 ( \62759 , \62749 , \62758 );
not \U$62417 ( \62760 , \62759 );
not \U$62418 ( \62761 , \62718 );
not \U$62419 ( \62762 , \62703 );
and \U$62420 ( \62763 , \62761 , \62762 );
and \U$62421 ( \62764 , \62718 , \62703 );
not \U$62422 ( \62765 , \62738 );
nor \U$62423 ( \62766 , \62764 , \62765 );
nor \U$62424 ( \62767 , \62763 , \62766 );
not \U$62425 ( \62768 , \62767 );
and \U$62426 ( \62769 , \62760 , \62768 );
and \U$62427 ( \62770 , \62759 , \62767 );
nor \U$62428 ( \62771 , \62769 , \62770 );
xor \U$62429 ( \62772 , \62747 , \62771 );
not \U$62430 ( \62773 , \62695 );
not \U$62431 ( \62774 , \62746 );
or \U$62432 ( \62775 , \62773 , \62774 );
or \U$62433 ( \62776 , \62746 , \62695 );
nand \U$62434 ( \62777 , \62775 , \62776 );
and \U$62435 ( \62778 , \13882 , RI9870498_86);
and \U$62436 ( \62779 , RI9870588_88, \13880 );
nor \U$62437 ( \62780 , \62778 , \62779 );
and \U$62438 ( \62781 , \62780 , \13359 );
not \U$62439 ( \62782 , \62780 );
and \U$62440 ( \62783 , \62782 , \13358 );
nor \U$62441 ( \62784 , \62781 , \62783 );
and \U$62442 ( \62785 , \15780 , RI9870768_92);
and \U$62443 ( \62786 , RI9870678_90, RI9873648_192);
nor \U$62444 ( \62787 , \62785 , \62786 );
not \U$62445 ( \62788 , \62787 );
not \U$62446 ( \62789 , RI9873558_190);
and \U$62447 ( \62790 , \62788 , \62789 );
and \U$62448 ( \62791 , \62787 , RI9873558_190);
nor \U$62449 ( \62792 , \62790 , \62791 );
or \U$62450 ( \62793 , \62784 , \62792 );
not \U$62451 ( \62794 , \62792 );
not \U$62452 ( \62795 , \62784 );
or \U$62453 ( \62796 , \62794 , \62795 );
and \U$62454 ( \62797 , \14937 , RI98703a8_84);
and \U$62455 ( \62798 , RI98702b8_82, \14935 );
nor \U$62456 ( \62799 , \62797 , \62798 );
and \U$62457 ( \62800 , \62799 , \14539 );
not \U$62458 ( \62801 , \62799 );
and \U$62459 ( \62802 , \62801 , \14538 );
nor \U$62460 ( \62803 , \62800 , \62802 );
nand \U$62461 ( \62804 , \62796 , \62803 );
nand \U$62462 ( \62805 , \62793 , \62804 );
not \U$62463 ( \62806 , \62717 );
not \U$62464 ( \62807 , \62711 );
or \U$62465 ( \62808 , \62806 , \62807 );
or \U$62466 ( \62809 , \62711 , \62717 );
nand \U$62467 ( \62810 , \62808 , \62809 );
xor \U$62468 ( \62811 , \62805 , \62810 );
xor \U$62469 ( \62812 , \62727 , \12619 );
xor \U$62470 ( \62813 , \62812 , \62735 );
and \U$62471 ( \62814 , \62811 , \62813 );
and \U$62472 ( \62815 , \62805 , \62810 );
or \U$62473 ( \62816 , \62814 , \62815 );
and \U$62474 ( \62817 , \62777 , \62816 );
nand \U$62475 ( \62818 , RI9870498_86, \13880 );
and \U$62476 ( \62819 , \62818 , \13359 );
not \U$62477 ( \62820 , \62818 );
and \U$62478 ( \62821 , \62820 , \13358 );
nor \U$62479 ( \62822 , \62819 , \62821 );
not \U$62480 ( \62823 , \62822 );
not \U$62481 ( \62824 , RI9873558_190);
and \U$62482 ( \62825 , \15780 , RI98702b8_82);
and \U$62483 ( \62826 , RI9870768_92, RI9873648_192);
nor \U$62484 ( \62827 , \62825 , \62826 );
not \U$62485 ( \62828 , \62827 );
or \U$62486 ( \62829 , \62824 , \62828 );
or \U$62487 ( \62830 , \62827 , RI9873558_190);
nand \U$62488 ( \62831 , \62829 , \62830 );
xor \U$62489 ( \62832 , \62831 , \13359 );
and \U$62490 ( \62833 , \14937 , RI9870588_88);
and \U$62491 ( \62834 , RI98703a8_84, \14935 );
nor \U$62492 ( \62835 , \62833 , \62834 );
and \U$62493 ( \62836 , \62835 , \14539 );
not \U$62494 ( \62837 , \62835 );
and \U$62495 ( \62838 , \62837 , \14538 );
nor \U$62496 ( \62839 , \62836 , \62838 );
xor \U$62497 ( \62840 , \62832 , \62839 );
nand \U$62498 ( \62841 , \62823 , \62840 );
not \U$62499 ( \62842 , \62792 );
not \U$62500 ( \62843 , \62803 );
or \U$62501 ( \62844 , \62842 , \62843 );
or \U$62502 ( \62845 , \62803 , \62792 );
nand \U$62503 ( \62846 , \62844 , \62845 );
not \U$62504 ( \62847 , \62846 );
not \U$62505 ( \62848 , \62784 );
and \U$62506 ( \62849 , \62847 , \62848 );
and \U$62507 ( \62850 , \62846 , \62784 );
nor \U$62508 ( \62851 , \62849 , \62850 );
not \U$62509 ( \62852 , \62851 );
xor \U$62510 ( \62853 , \62831 , \13359 );
and \U$62511 ( \62854 , \62853 , \62839 );
and \U$62512 ( \62855 , \62831 , \13359 );
or \U$62513 ( \62856 , \62854 , \62855 );
not \U$62514 ( \62857 , \62856 );
and \U$62515 ( \62858 , \62852 , \62857 );
and \U$62516 ( \62859 , \62851 , \62856 );
nor \U$62517 ( \62860 , \62858 , \62859 );
xor \U$62518 ( \62861 , \62841 , \62860 );
and \U$62519 ( \62862 , \14937 , RI9870498_86);
and \U$62520 ( \62863 , RI9870588_88, \14935 );
nor \U$62521 ( \62864 , \62862 , \62863 );
and \U$62522 ( \62865 , \62864 , \14539 );
not \U$62523 ( \62866 , \62864 );
and \U$62524 ( \62867 , \62866 , \14538 );
nor \U$62525 ( \62868 , \62865 , \62867 );
not \U$62526 ( \62869 , \62868 );
and \U$62527 ( \62870 , \15780 , RI98703a8_84);
and \U$62528 ( \62871 , RI98702b8_82, RI9873648_192);
nor \U$62529 ( \62872 , \62870 , \62871 );
not \U$62530 ( \62873 , \62872 );
not \U$62531 ( \62874 , RI9873558_190);
and \U$62532 ( \62875 , \62873 , \62874 );
and \U$62533 ( \62876 , \62872 , RI9873558_190);
nor \U$62534 ( \62877 , \62875 , \62876 );
nor \U$62535 ( \62878 , \62869 , \62877 );
not \U$62536 ( \62879 , \62822 );
not \U$62537 ( \62880 , \62840 );
or \U$62538 ( \62881 , \62879 , \62880 );
or \U$62539 ( \62882 , \62840 , \62822 );
nand \U$62540 ( \62883 , \62881 , \62882 );
xor \U$62541 ( \62884 , \62878 , \62883 );
not \U$62542 ( \62885 , RI9873558_190);
and \U$62543 ( \62886 , \15780 , RI9870588_88);
and \U$62544 ( \62887 , RI98703a8_84, RI9873648_192);
nor \U$62545 ( \62888 , \62886 , \62887 );
not \U$62546 ( \62889 , \62888 );
or \U$62547 ( \62890 , \62885 , \62889 );
or \U$62548 ( \62891 , \62888 , RI9873558_190);
nand \U$62549 ( \62892 , \62890 , \62891 );
nand \U$62550 ( \62893 , \14538 , \62892 );
not \U$62551 ( \62894 , \62868 );
not \U$62552 ( \62895 , \62877 );
and \U$62553 ( \62896 , \62894 , \62895 );
and \U$62554 ( \62897 , \62868 , \62877 );
nor \U$62555 ( \62898 , \62896 , \62897 );
xnor \U$62556 ( \62899 , \62893 , \62898 );
nand \U$62557 ( \62900 , RI9870498_86, \14935 );
and \U$62558 ( \62901 , \62900 , \14539 );
not \U$62559 ( \62902 , \62900 );
and \U$62560 ( \62903 , \62902 , \14538 );
nor \U$62561 ( \62904 , \62901 , \62903 );
and \U$62562 ( \62905 , \62892 , \14538 );
not \U$62563 ( \62906 , \62892 );
and \U$62564 ( \62907 , \62906 , \14539 );
nor \U$62565 ( \62908 , \62905 , \62907 );
xor \U$62566 ( \62909 , \62904 , \62908 );
nand \U$62567 ( \62910 , RI9870498_86, RI9873648_192);
and \U$62568 ( \62911 , \62910 , RI9873558_190);
not \U$62569 ( \62912 , RI9873558_190);
and \U$62570 ( \62913 , \15780 , RI9870498_86);
and \U$62571 ( \62914 , RI9870588_88, RI9873648_192);
nor \U$62572 ( \62915 , \62913 , \62914 );
not \U$62573 ( \62916 , \62915 );
or \U$62574 ( \62917 , \62912 , \62916 );
or \U$62575 ( \62918 , \62915 , RI9873558_190);
nand \U$62576 ( \62919 , \62917 , \62918 );
and \U$62577 ( \62920 , \62911 , \62919 );
and \U$62578 ( \62921 , \62909 , \62920 );
and \U$62579 ( \62922 , \62904 , \62908 );
nor \U$62580 ( \62923 , \62921 , \62922 );
or \U$62581 ( \62924 , \62899 , \62923 );
or \U$62582 ( \62925 , \62893 , \62898 );
nand \U$62583 ( \62926 , \62924 , \62925 );
and \U$62584 ( \62927 , \62884 , \62926 );
and \U$62585 ( \62928 , \62878 , \62883 );
nor \U$62586 ( \62929 , \62927 , \62928 );
and \U$62587 ( \62930 , \62861 , \62929 );
and \U$62588 ( \62931 , \62841 , \62860 );
nor \U$62589 ( \62932 , \62930 , \62931 );
not \U$62590 ( \62933 , \62856 );
nor \U$62591 ( \62934 , \62933 , \62851 );
xor \U$62592 ( \62935 , \62805 , \62810 );
xor \U$62593 ( \62936 , \62935 , \62813 );
xor \U$62594 ( \62937 , \62934 , \62936 );
and \U$62595 ( \62938 , \62932 , \62937 );
and \U$62596 ( \62939 , \62934 , \62936 );
nor \U$62597 ( \62940 , \62938 , \62939 );
xnor \U$62598 ( \62941 , \62816 , \62777 );
nor \U$62599 ( \62942 , \62940 , \62941 );
nor \U$62600 ( \62943 , \62817 , \62942 );
and \U$62601 ( \62944 , \62772 , \62943 );
and \U$62602 ( \62945 , \62747 , \62771 );
nor \U$62603 ( \62946 , \62944 , \62945 );
not \U$62604 ( \62947 , \62759 );
nor \U$62605 ( \62948 , \62947 , \62767 );
xor \U$62606 ( \62949 , \62571 , \62599 );
xor \U$62607 ( \62950 , \62519 , \62526 );
xor \U$62608 ( \62951 , \62950 , \62550 );
xor \U$62609 ( \62952 , \62949 , \62951 );
xor \U$62610 ( \62953 , \62508 , \11686 );
xor \U$62611 ( \62954 , \62953 , \62516 );
and \U$62612 ( \62955 , \62755 , \62954 );
xor \U$62613 ( \62956 , \62508 , \11686 );
xor \U$62614 ( \62957 , \62956 , \62516 );
and \U$62615 ( \62958 , \62757 , \62957 );
and \U$62616 ( \62959 , \62755 , \62757 );
or \U$62617 ( \62960 , \62955 , \62958 , \62959 );
xor \U$62618 ( \62961 , \62952 , \62960 );
xor \U$62619 ( \62962 , \62948 , \62961 );
and \U$62620 ( \62963 , \62946 , \62962 );
and \U$62621 ( \62964 , \62948 , \62961 );
nor \U$62622 ( \62965 , \62963 , \62964 );
xor \U$62623 ( \62966 , \62949 , \62951 );
and \U$62624 ( \62967 , \62966 , \62960 );
and \U$62625 ( \62968 , \62949 , \62951 );
nor \U$62626 ( \62969 , \62967 , \62968 );
not \U$62627 ( \62970 , \62657 );
not \U$62628 ( \62971 , \62660 );
and \U$62629 ( \62972 , \62970 , \62971 );
and \U$62630 ( \62973 , \62657 , \62660 );
nor \U$62631 ( \62974 , \62972 , \62973 );
xnor \U$62632 ( \62975 , \62969 , \62974 );
or \U$62633 ( \62976 , \62965 , \62975 );
or \U$62634 ( \62977 , \62969 , \62974 );
nand \U$62635 ( \62978 , \62976 , \62977 );
and \U$62636 ( \62979 , \62663 , \62978 );
nor \U$62637 ( \62980 , \62662 , \62979 );
not \U$62638 ( \62981 , \62651 );
nand \U$62639 ( \62982 , \62981 , \62603 );
xor \U$62640 ( \62983 , \62329 , \62336 );
xor \U$62641 ( \62984 , \62983 , \62364 );
xor \U$62642 ( \62985 , \62480 , \62487 );
xor \U$62643 ( \62986 , \62984 , \62985 );
not \U$62644 ( \62987 , \62986 );
xor \U$62645 ( \62988 , \62629 , \62639 );
and \U$62646 ( \62989 , \62988 , \62650 );
and \U$62647 ( \62990 , \62629 , \62639 );
or \U$62648 ( \62991 , \62989 , \62990 );
not \U$62649 ( \62992 , \62991 );
and \U$62650 ( \62993 , \62987 , \62992 );
and \U$62651 ( \62994 , \62986 , \62991 );
nor \U$62652 ( \62995 , \62993 , \62994 );
xnor \U$62653 ( \62996 , \62982 , \62995 );
or \U$62654 ( \62997 , \62980 , \62996 );
or \U$62655 ( \62998 , \62982 , \62995 );
nand \U$62656 ( \62999 , \62997 , \62998 );
not \U$62657 ( \63000 , \62986 );
nor \U$62658 ( \63001 , \63000 , \62991 );
xor \U$62659 ( \63002 , \62416 , \62492 );
xor \U$62660 ( \63003 , \63002 , \62495 );
xor \U$62661 ( \63004 , \63001 , \63003 );
and \U$62662 ( \63005 , \62999 , \63004 );
and \U$62663 ( \63006 , \63001 , \63003 );
nor \U$62664 ( \63007 , \63005 , \63006 );
or \U$62665 ( \63008 , \62500 , \63007 );
nand \U$62666 ( \63009 , \62499 , \63008 );
xnor \U$62667 ( \63010 , \62172 , \62239 );
not \U$62668 ( \63011 , \63010 );
not \U$62669 ( \63012 , \62177 );
and \U$62670 ( \63013 , \63011 , \63012 );
and \U$62671 ( \63014 , \63010 , \62177 );
nor \U$62672 ( \63015 , \63013 , \63014 );
not \U$62673 ( \63016 , \63015 );
xor \U$62674 ( \63017 , \62034 , \62057 );
xor \U$62675 ( \63018 , \63017 , \62083 );
and \U$62676 ( \63019 , \62391 , \62395 );
not \U$62677 ( \63020 , \62391 );
not \U$62678 ( \63021 , \62395 );
and \U$62679 ( \63022 , \63020 , \63021 );
nor \U$62680 ( \63023 , \63022 , \62406 );
nor \U$62681 ( \63024 , \63019 , \63023 );
xor \U$62682 ( \63025 , \63018 , \63024 );
not \U$62683 ( \63026 , \63025 );
or \U$62684 ( \63027 , \63016 , \63026 );
or \U$62685 ( \63028 , \63025 , \63015 );
nand \U$62686 ( \63029 , \63027 , \63028 );
not \U$62687 ( \63030 , \62301 );
not \U$62688 ( \63031 , \62411 );
or \U$62689 ( \63032 , \63030 , \63031 );
or \U$62690 ( \63033 , \62411 , \62301 );
nand \U$62691 ( \63034 , \63033 , \62388 );
nand \U$62692 ( \63035 , \63032 , \63034 );
xor \U$62693 ( \63036 , \63029 , \63035 );
and \U$62694 ( \63037 , \63009 , \63036 );
and \U$62695 ( \63038 , \63029 , \63035 );
nor \U$62696 ( \63039 , \63037 , \63038 );
not \U$62697 ( \63040 , \63015 );
not \U$62698 ( \63041 , \63018 );
and \U$62699 ( \63042 , \63040 , \63041 );
and \U$62700 ( \63043 , \63015 , \63018 );
nor \U$62701 ( \63044 , \63043 , \63024 );
nor \U$62702 ( \63045 , \63042 , \63044 );
xnor \U$62703 ( \63046 , \62241 , \62156 );
not \U$62704 ( \63047 , \63046 );
not \U$62705 ( \63048 , \62153 );
and \U$62706 ( \63049 , \63047 , \63048 );
and \U$62707 ( \63050 , \63046 , \62153 );
nor \U$62708 ( \63051 , \63049 , \63050 );
xnor \U$62709 ( \63052 , \63045 , \63051 );
or \U$62710 ( \63053 , \63039 , \63052 );
or \U$62711 ( \63054 , \63045 , \63051 );
nand \U$62712 ( \63055 , \63053 , \63054 );
and \U$62713 ( \63056 , \62245 , \63055 );
nor \U$62714 ( \63057 , \62244 , \63056 );
or \U$62715 ( \63058 , \62147 , \63057 );
nand \U$62716 ( \63059 , \62146 , \63058 );
and \U$62717 ( \63060 , \62126 , \63059 );
nor \U$62718 ( \63061 , \62125 , \63060 );
and \U$62719 ( \63062 , \61769 , \61771 );
xor \U$62720 ( \63063 , \61879 , \61883 );
and \U$62721 ( \63064 , \63063 , \61896 );
and \U$62722 ( \63065 , \61879 , \61883 );
or \U$62723 ( \63066 , \63064 , \63065 );
xnor \U$62724 ( \63067 , \63062 , \63066 );
not \U$62725 ( \63068 , \63067 );
xor \U$62726 ( \63069 , \61645 , \61753 );
xor \U$62727 ( \63070 , \63069 , \61756 );
not \U$62728 ( \63071 , \63070 );
and \U$62729 ( \63072 , \63068 , \63071 );
and \U$62730 ( \63073 , \63067 , \63070 );
nor \U$62731 ( \63074 , \63072 , \63073 );
xor \U$62732 ( \63075 , \61772 , \61897 );
and \U$62733 ( \63076 , \63075 , \62012 );
and \U$62734 ( \63077 , \61772 , \61897 );
nor \U$62735 ( \63078 , \63076 , \63077 );
xnor \U$62736 ( \63079 , \63074 , \63078 );
or \U$62737 ( \63080 , \63061 , \63079 );
or \U$62738 ( \63081 , \63074 , \63078 );
nand \U$62739 ( \63082 , \63080 , \63081 );
xor \U$62740 ( \63083 , \61644 , \61759 );
xor \U$62741 ( \63084 , \63083 , \61762 );
not \U$62742 ( \63085 , \63062 );
not \U$62743 ( \63086 , \63070 );
or \U$62744 ( \63087 , \63085 , \63086 );
or \U$62745 ( \63088 , \63070 , \63062 );
nand \U$62746 ( \63089 , \63088 , \63066 );
nand \U$62747 ( \63090 , \63087 , \63089 );
xor \U$62748 ( \63091 , \63084 , \63090 );
and \U$62749 ( \63092 , \63082 , \63091 );
and \U$62750 ( \63093 , \63084 , \63090 );
nor \U$62751 ( \63094 , \63092 , \63093 );
or \U$62752 ( \63095 , \61767 , \63094 );
nand \U$62753 ( \63096 , \61766 , \63095 );
or \U$62754 ( \63097 , \61635 , \61480 );
not \U$62755 ( \63098 , \61480 );
not \U$62756 ( \63099 , \61635 );
or \U$62757 ( \63100 , \63098 , \63099 );
nand \U$62758 ( \63101 , \63100 , \61598 );
nand \U$62759 ( \63102 , \63097 , \63101 );
xor \U$62760 ( \63103 , \61217 , \61352 );
xor \U$62761 ( \63104 , \63103 , \61357 );
xor \U$62762 ( \63105 , \61149 , \61155 );
xor \U$62763 ( \63106 , \63105 , \61171 );
xor \U$62764 ( \63107 , \63104 , \63106 );
or \U$62765 ( \63108 , \61631 , \61609 );
not \U$62766 ( \63109 , \61609 );
not \U$62767 ( \63110 , \61631 );
or \U$62768 ( \63111 , \63109 , \63110 );
nand \U$62769 ( \63112 , \63111 , \61616 );
nand \U$62770 ( \63113 , \63108 , \63112 );
xor \U$62771 ( \63114 , \63107 , \63113 );
xor \U$62772 ( \63115 , \63102 , \63114 );
and \U$62773 ( \63116 , \63096 , \63115 );
and \U$62774 ( \63117 , \63102 , \63114 );
nor \U$62775 ( \63118 , \63116 , \63117 );
xor \U$62776 ( \63119 , \63104 , \63106 );
and \U$62777 ( \63120 , \63119 , \63113 );
and \U$62778 ( \63121 , \63104 , \63106 );
nor \U$62779 ( \63122 , \63120 , \63121 );
xnor \U$62780 ( \63123 , \61194 , \61360 );
not \U$62781 ( \63124 , \63123 );
not \U$62782 ( \63125 , \61197 );
and \U$62783 ( \63126 , \63124 , \63125 );
and \U$62784 ( \63127 , \63123 , \61197 );
nor \U$62785 ( \63128 , \63126 , \63127 );
xnor \U$62786 ( \63129 , \63122 , \63128 );
or \U$62787 ( \63130 , \63118 , \63129 );
or \U$62788 ( \63131 , \63122 , \63128 );
nand \U$62789 ( \63132 , \63130 , \63131 );
and \U$62790 ( \63133 , \61364 , \63132 );
nor \U$62791 ( \63134 , \61363 , \63133 );
or \U$62792 ( \63135 , \61186 , \63134 );
nand \U$62793 ( \63136 , \61185 , \63135 );
and \U$62794 ( \63137 , \61040 , \63136 );
nor \U$62795 ( \63138 , \61039 , \63137 );
or \U$62796 ( \63139 , \61015 , \63138 );
nand \U$62797 ( \63140 , \61014 , \63139 );
xor \U$62798 ( \63141 , \60300 , \60453 );
xor \U$62799 ( \63142 , \63141 , \60456 );
and \U$62800 ( \63143 , \60849 , \60851 );
xor \U$62801 ( \63144 , \63142 , \63143 );
not \U$62802 ( \63145 , \60838 );
not \U$62803 ( \63146 , \60832 );
or \U$62804 ( \63147 , \63145 , \63146 );
or \U$62805 ( \63148 , \60832 , \60838 );
nand \U$62806 ( \63149 , \63148 , \60828 );
nand \U$62807 ( \63150 , \63147 , \63149 );
xor \U$62808 ( \63151 , \63144 , \63150 );
not \U$62809 ( \63152 , \60852 );
or \U$62810 ( \63153 , \60842 , \63152 );
not \U$62811 ( \63154 , \63152 );
not \U$62812 ( \63155 , \60842 );
or \U$62813 ( \63156 , \63154 , \63155 );
nand \U$62814 ( \63157 , \63156 , \60819 );
nand \U$62815 ( \63158 , \63153 , \63157 );
xor \U$62816 ( \63159 , \63151 , \63158 );
and \U$62817 ( \63160 , \63140 , \63159 );
and \U$62818 ( \63161 , \63158 , \63151 );
nor \U$62819 ( \63162 , \63160 , \63161 );
xor \U$62820 ( \63163 , \63142 , \63143 );
and \U$62821 ( \63164 , \63163 , \63150 );
and \U$62822 ( \63165 , \63142 , \63143 );
nor \U$62823 ( \63166 , \63164 , \63165 );
xnor \U$62824 ( \63167 , \60296 , \60459 );
not \U$62825 ( \63168 , \63167 );
not \U$62826 ( \63169 , \60293 );
and \U$62827 ( \63170 , \63168 , \63169 );
and \U$62828 ( \63171 , \63167 , \60293 );
nor \U$62829 ( \63172 , \63170 , \63171 );
xnor \U$62830 ( \63173 , \63166 , \63172 );
or \U$62831 ( \63174 , \63162 , \63173 );
or \U$62832 ( \63175 , \63166 , \63172 );
nand \U$62833 ( \63176 , \63174 , \63175 );
and \U$62834 ( \63177 , \60463 , \63176 );
nor \U$62835 ( \63178 , \60462 , \63177 );
or \U$62836 ( \63179 , \60290 , \63178 );
nand \U$62837 ( \63180 , \60289 , \63179 );
not \U$62838 ( \63181 , \60276 );
not \U$62839 ( \63182 , \60284 );
or \U$62840 ( \63183 , \63181 , \63182 );
or \U$62841 ( \63184 , \60284 , \60276 );
nand \U$62842 ( \63185 , \63184 , \60280 );
nand \U$62843 ( \63186 , \63183 , \63185 );
xor \U$62844 ( \63187 , \59730 , \59912 );
xor \U$62845 ( \63188 , \63187 , \59915 );
xor \U$62846 ( \63189 , \63186 , \63188 );
and \U$62847 ( \63190 , \63180 , \63189 );
and \U$62848 ( \63191 , \63186 , \63188 );
nor \U$62849 ( \63192 , \63190 , \63191 );
or \U$62850 ( \63193 , \59920 , \63192 );
nand \U$62851 ( \63194 , \59919 , \63193 );
and \U$62852 ( \63195 , \59722 , \63194 );
nor \U$62853 ( \63196 , \59721 , \63195 );
xor \U$62854 ( \63197 , \59294 , \59299 );
and \U$62855 ( \63198 , \63197 , \59492 );
and \U$62856 ( \63199 , \59294 , \59299 );
nor \U$62857 ( \63200 , \63198 , \63199 );
xnor \U$62858 ( \63201 , \59096 , \59286 );
not \U$62859 ( \63202 , \63201 );
not \U$62860 ( \63203 , \59099 );
and \U$62861 ( \63204 , \63202 , \63203 );
and \U$62862 ( \63205 , \63201 , \59099 );
nor \U$62863 ( \63206 , \63204 , \63205 );
xnor \U$62864 ( \63207 , \63200 , \63206 );
or \U$62865 ( \63208 , \63196 , \63207 );
or \U$62866 ( \63209 , \63200 , \63206 );
nand \U$62867 ( \63210 , \63208 , \63209 );
and \U$62868 ( \63211 , \59290 , \63210 );
nor \U$62869 ( \63212 , \59289 , \63211 );
or \U$62870 ( \63213 , \59088 , \63212 );
nand \U$62871 ( \63214 , \59087 , \63213 );
and \U$62872 ( \63215 , \58837 , \63214 );
nor \U$62873 ( \63216 , \58836 , \63215 );
not \U$62874 ( \63217 , \58822 );
nand \U$62875 ( \63218 , \63217 , \58825 );
not \U$62876 ( \63219 , \58235 );
not \U$62877 ( \63220 , \58520 );
and \U$62878 ( \63221 , \63219 , \63220 );
and \U$62879 ( \63222 , \58235 , \58520 );
nor \U$62880 ( \63223 , \63221 , \63222 );
xnor \U$62881 ( \63224 , \63218 , \63223 );
or \U$62882 ( \63225 , \63216 , \63224 );
or \U$62883 ( \63226 , \63218 , \63223 );
nand \U$62884 ( \63227 , \63225 , \63226 );
and \U$62885 ( \63228 , \58523 , \63227 );
nor \U$62886 ( \63229 , \58522 , \63228 );
or \U$62887 ( \63230 , \58229 , \63229 );
nand \U$62888 ( \63231 , \58228 , \63230 );
not \U$62889 ( \63232 , \58223 );
nor \U$62890 ( \63233 , \63232 , \58218 );
xor \U$62891 ( \63234 , \57415 , \57417 );
xor \U$62892 ( \63235 , \63234 , \57666 );
xor \U$62893 ( \63236 , \63233 , \63235 );
and \U$62894 ( \63237 , \63231 , \63236 );
and \U$62895 ( \63238 , \63233 , \63235 );
nor \U$62896 ( \63239 , \63237 , \63238 );
or \U$62897 ( \63240 , \57671 , \63239 );
nand \U$62898 ( \63241 , \57670 , \63240 );
xor \U$62899 ( \63242 , \56606 , \56859 );
xor \U$62900 ( \63243 , \63242 , \56862 );
and \U$62901 ( \63244 , \57406 , \57408 );
xor \U$62902 ( \63245 , \63243 , \63244 );
xor \U$62903 ( \63246 , \56881 , \56885 );
and \U$62904 ( \63247 , \63246 , \57121 );
and \U$62905 ( \63248 , \56881 , \56885 );
or \U$62906 ( \63249 , \63247 , \63248 );
xor \U$62907 ( \63250 , \63245 , \63249 );
not \U$62908 ( \63251 , \57409 );
not \U$62909 ( \63252 , \57122 );
or \U$62910 ( \63253 , \63251 , \63252 );
or \U$62911 ( \63254 , \57122 , \57409 );
nand \U$62912 ( \63255 , \63254 , \57402 );
nand \U$62913 ( \63256 , \63253 , \63255 );
xor \U$62914 ( \63257 , \63250 , \63256 );
and \U$62915 ( \63258 , \63241 , \63257 );
and \U$62916 ( \63259 , \63256 , \63250 );
nor \U$62917 ( \63260 , \63258 , \63259 );
xor \U$62918 ( \63261 , \63243 , \63244 );
and \U$62919 ( \63262 , \63261 , \63249 );
and \U$62920 ( \63263 , \63243 , \63244 );
nor \U$62921 ( \63264 , \63262 , \63263 );
xnor \U$62922 ( \63265 , \56598 , \56865 );
not \U$62923 ( \63266 , \63265 );
not \U$62924 ( \63267 , \56587 );
and \U$62925 ( \63268 , \63266 , \63267 );
and \U$62926 ( \63269 , \63265 , \56587 );
nor \U$62927 ( \63270 , \63268 , \63269 );
xnor \U$62928 ( \63271 , \63264 , \63270 );
or \U$62929 ( \63272 , \63260 , \63271 );
or \U$62930 ( \63273 , \63264 , \63270 );
nand \U$62931 ( \63274 , \63272 , \63273 );
and \U$62932 ( \63275 , \56869 , \63274 );
nor \U$62933 ( \63276 , \56868 , \63275 );
not \U$62934 ( \63277 , \55973 );
not \U$62935 ( \63278 , \56287 );
or \U$62936 ( \63279 , \63277 , \63278 );
or \U$62937 ( \63280 , \56287 , \55973 );
nand \U$62938 ( \63281 , \63279 , \63280 );
not \U$62939 ( \63282 , \63281 );
not \U$62940 ( \63283 , \55967 );
and \U$62941 ( \63284 , \63282 , \63283 );
and \U$62942 ( \63285 , \63281 , \55967 );
nor \U$62943 ( \63286 , \63284 , \63285 );
and \U$62944 ( \63287 , \56293 , \56299 );
not \U$62945 ( \63288 , \56293 );
not \U$62946 ( \63289 , \56299 );
and \U$62947 ( \63290 , \63288 , \63289 );
nor \U$62948 ( \63291 , \63290 , \56578 );
nor \U$62949 ( \63292 , \63287 , \63291 );
xnor \U$62950 ( \63293 , \63286 , \63292 );
or \U$62951 ( \63294 , \63276 , \63293 );
or \U$62952 ( \63295 , \63286 , \63292 );
nand \U$62953 ( \63296 , \63294 , \63295 );
and \U$62954 ( \63297 , \56291 , \63296 );
nor \U$62955 ( \63298 , \56290 , \63297 );
not \U$62956 ( \63299 , \55597 );
nand \U$62957 ( \63300 , \63299 , \55957 );
and \U$62958 ( \63301 , \63300 , \55936 );
not \U$62959 ( \63302 , \55957 );
and \U$62960 ( \63303 , \63302 , \55597 );
nor \U$62961 ( \63304 , \63301 , \63303 );
not \U$62962 ( \63305 , \54919 );
not \U$62963 ( \63306 , \54631 );
or \U$62964 ( \63307 , \63305 , \63306 );
or \U$62965 ( \63308 , \54631 , \54919 );
nand \U$62966 ( \63309 , \63307 , \63308 );
not \U$62967 ( \63310 , \63309 );
not \U$62968 ( \63311 , \54637 );
and \U$62969 ( \63312 , \63310 , \63311 );
and \U$62970 ( \63313 , \63309 , \54637 );
nor \U$62971 ( \63314 , \63312 , \63313 );
not \U$62972 ( \63315 , \63314 );
xor \U$62973 ( \63316 , \55236 , \55585 );
and \U$62974 ( \63317 , \63316 , \55596 );
and \U$62975 ( \63318 , \55236 , \55585 );
or \U$62976 ( \63319 , \63317 , \63318 );
not \U$62977 ( \63320 , \63319 );
or \U$62978 ( \63321 , \63315 , \63320 );
or \U$62979 ( \63322 , \63319 , \63314 );
nand \U$62980 ( \63323 , \63321 , \63322 );
not \U$62981 ( \63324 , \63323 );
or \U$62982 ( \63325 , \55946 , \55953 );
not \U$62983 ( \63326 , \55953 );
not \U$62984 ( \63327 , \55946 );
or \U$62985 ( \63328 , \63326 , \63327 );
nand \U$62986 ( \63329 , \63328 , \55941 );
nand \U$62987 ( \63330 , \63325 , \63329 );
xor \U$62988 ( \63331 , \54681 , \54901 );
xor \U$62989 ( \63332 , \63331 , \54916 );
and \U$62990 ( \63333 , \55590 , \63332 );
xor \U$62991 ( \63334 , \54681 , \54901 );
xor \U$62992 ( \63335 , \63334 , \54916 );
and \U$62993 ( \63336 , \55594 , \63335 );
and \U$62994 ( \63337 , \55590 , \55594 );
or \U$62995 ( \63338 , \63333 , \63336 , \63337 );
xnor \U$62996 ( \63339 , \63330 , \63338 );
not \U$62997 ( \63340 , \63339 );
xor \U$62998 ( \63341 , \54290 , \54520 );
xor \U$62999 ( \63342 , \63341 , \54534 );
xor \U$63000 ( \63343 , \54923 , \54930 );
xor \U$63001 ( \63344 , \63342 , \63343 );
not \U$63002 ( \63345 , \63344 );
and \U$63003 ( \63346 , \63340 , \63345 );
and \U$63004 ( \63347 , \63339 , \63344 );
nor \U$63005 ( \63348 , \63346 , \63347 );
not \U$63006 ( \63349 , \63348 );
and \U$63007 ( \63350 , \63324 , \63349 );
and \U$63008 ( \63351 , \63323 , \63348 );
nor \U$63009 ( \63352 , \63350 , \63351 );
xnor \U$63010 ( \63353 , \63304 , \63352 );
or \U$63011 ( \63354 , \63298 , \63353 );
or \U$63012 ( \63355 , \63304 , \63352 );
nand \U$63013 ( \63356 , \63354 , \63355 );
or \U$63014 ( \63357 , \63348 , \63314 );
not \U$63015 ( \63358 , \63314 );
not \U$63016 ( \63359 , \63348 );
or \U$63017 ( \63360 , \63358 , \63359 );
nand \U$63018 ( \63361 , \63360 , \63319 );
nand \U$63019 ( \63362 , \63357 , \63361 );
xor \U$63020 ( \63363 , \54921 , \54935 );
xor \U$63021 ( \63364 , \63363 , \54940 );
xor \U$63022 ( \63365 , \54537 , \54539 );
xor \U$63023 ( \63366 , \63365 , \54564 );
xor \U$63024 ( \63367 , \63364 , \63366 );
not \U$63025 ( \63368 , \63338 );
not \U$63026 ( \63369 , \63344 );
or \U$63027 ( \63370 , \63368 , \63369 );
or \U$63028 ( \63371 , \63344 , \63338 );
nand \U$63029 ( \63372 , \63371 , \63330 );
nand \U$63030 ( \63373 , \63370 , \63372 );
xor \U$63031 ( \63374 , \63367 , \63373 );
xor \U$63032 ( \63375 , \63362 , \63374 );
and \U$63033 ( \63376 , \63356 , \63375 );
and \U$63034 ( \63377 , \63362 , \63374 );
nor \U$63035 ( \63378 , \63376 , \63377 );
xor \U$63036 ( \63379 , \63364 , \63366 );
and \U$63037 ( \63380 , \63379 , \63373 );
and \U$63038 ( \63381 , \63364 , \63366 );
nor \U$63039 ( \63382 , \63380 , \63381 );
xnor \U$63040 ( \63383 , \54943 , \54611 );
not \U$63041 ( \63384 , \63383 );
not \U$63042 ( \63385 , \54608 );
and \U$63043 ( \63386 , \63384 , \63385 );
and \U$63044 ( \63387 , \63383 , \54608 );
nor \U$63045 ( \63388 , \63386 , \63387 );
xnor \U$63046 ( \63389 , \63382 , \63388 );
or \U$63047 ( \63390 , \63378 , \63389 );
or \U$63048 ( \63391 , \63382 , \63388 );
nand \U$63049 ( \63392 , \63390 , \63391 );
and \U$63050 ( \63393 , \54947 , \63392 );
nor \U$63051 ( \63394 , \54946 , \63393 );
or \U$63052 ( \63395 , \54593 , \63394 );
nand \U$63053 ( \63396 , \54592 , \63395 );
or \U$63054 ( \63397 , \54224 , \53537 );
not \U$63055 ( \63398 , \53537 );
not \U$63056 ( \63399 , \54224 );
or \U$63057 ( \63400 , \63398 , \63399 );
nand \U$63058 ( \63401 , \63400 , \54193 );
nand \U$63059 ( \63402 , \63397 , \63401 );
not \U$63060 ( \63403 , \53110 );
not \U$63061 ( \63404 , \52738 );
or \U$63062 ( \63405 , \63403 , \63404 );
or \U$63063 ( \63406 , \52738 , \53110 );
nand \U$63064 ( \63407 , \63405 , \63406 );
or \U$63065 ( \63408 , \54220 , \54209 );
not \U$63066 ( \63409 , \54209 );
not \U$63067 ( \63410 , \54220 );
or \U$63068 ( \63411 , \63409 , \63410 );
nand \U$63069 ( \63412 , \63411 , \54202 );
nand \U$63070 ( \63413 , \63408 , \63412 );
xor \U$63071 ( \63414 , \63407 , \63413 );
xor \U$63072 ( \63415 , \53452 , \53454 );
xor \U$63073 ( \63416 , \63415 , \53471 );
xor \U$63074 ( \63417 , \63414 , \63416 );
xor \U$63075 ( \63418 , \63402 , \63417 );
and \U$63076 ( \63419 , \63396 , \63418 );
and \U$63077 ( \63420 , \63402 , \63417 );
nor \U$63078 ( \63421 , \63419 , \63420 );
xor \U$63079 ( \63422 , \63407 , \63413 );
and \U$63080 ( \63423 , \63422 , \63416 );
and \U$63081 ( \63424 , \63407 , \63413 );
nor \U$63082 ( \63425 , \63423 , \63424 );
not \U$63083 ( \63426 , \53517 );
not \U$63084 ( \63427 , \53524 );
and \U$63085 ( \63428 , \63426 , \63427 );
and \U$63086 ( \63429 , \53517 , \53524 );
nor \U$63087 ( \63430 , \63428 , \63429 );
xnor \U$63088 ( \63431 , \63425 , \63430 );
or \U$63089 ( \63432 , \63421 , \63431 );
or \U$63090 ( \63433 , \63425 , \63430 );
nand \U$63091 ( \63434 , \63432 , \63433 );
and \U$63092 ( \63435 , \53527 , \63434 );
nor \U$63093 ( \63436 , \53526 , \63435 );
not \U$63094 ( \63437 , \53478 );
nand \U$63095 ( \63438 , \63437 , \53503 );
xor \U$63096 ( \63439 , \52704 , \52706 );
xor \U$63097 ( \63440 , \63439 , \52709 );
not \U$63098 ( \63441 , \63440 );
xor \U$63099 ( \63442 , \53481 , \53499 );
and \U$63100 ( \63443 , \63442 , \53502 );
and \U$63101 ( \63444 , \53481 , \53499 );
nor \U$63102 ( \63445 , \63443 , \63444 );
not \U$63103 ( \63446 , \63445 );
and \U$63104 ( \63447 , \63441 , \63446 );
and \U$63105 ( \63448 , \63440 , \63445 );
nor \U$63106 ( \63449 , \63447 , \63448 );
xnor \U$63107 ( \63450 , \63438 , \63449 );
or \U$63108 ( \63451 , \63436 , \63450 );
or \U$63109 ( \63452 , \63438 , \63449 );
nand \U$63110 ( \63453 , \63451 , \63452 );
not \U$63111 ( \63454 , \63440 );
nor \U$63112 ( \63455 , \63454 , \63445 );
not \U$63113 ( \63456 , \52712 );
not \U$63114 ( \63457 , \52308 );
or \U$63115 ( \63458 , \63456 , \63457 );
or \U$63116 ( \63459 , \52308 , \52712 );
nand \U$63117 ( \63460 , \63458 , \63459 );
xor \U$63118 ( \63461 , \63455 , \63460 );
and \U$63119 ( \63462 , \63453 , \63461 );
and \U$63120 ( \63463 , \63455 , \63460 );
nor \U$63121 ( \63464 , \63462 , \63463 );
or \U$63122 ( \63465 , \52715 , \63464 );
nand \U$63123 ( \63466 , \52714 , \63465 );
and \U$63124 ( \63467 , \52288 , \63466 );
nor \U$63125 ( \63468 , \52287 , \63467 );
and \U$63126 ( \63469 , \51851 , \63468 );
and \U$63127 ( \63470 , \51837 , \51850 );
nor \U$63128 ( \63471 , \63469 , \63470 );
not \U$63129 ( \63472 , \51841 );
nor \U$63130 ( \63473 , \63472 , \51846 );
xor \U$63131 ( \63474 , \51034 , \51036 );
xor \U$63132 ( \63475 , \63474 , \51039 );
xor \U$63133 ( \63476 , \63473 , \63475 );
and \U$63134 ( \63477 , \63471 , \63476 );
and \U$63135 ( \63478 , \63473 , \63475 );
nor \U$63136 ( \63479 , \63477 , \63478 );
not \U$63137 ( \63480 , \63479 );
and \U$63138 ( \63481 , \51044 , \63480 );
nor \U$63139 ( \63482 , \51043 , \63481 );
not \U$63140 ( \63483 , \50562 );
nand \U$63141 ( \63484 , \63483 , \50565 );
xor \U$63142 ( \63485 , \50140 , \50145 );
xor \U$63143 ( \63486 , \63485 , \50152 );
and \U$63144 ( \63487 , \63484 , \63486 );
not \U$63145 ( \63488 , \63484 );
not \U$63146 ( \63489 , \63486 );
and \U$63147 ( \63490 , \63488 , \63489 );
nor \U$63148 ( \63491 , \63487 , \63490 );
or \U$63149 ( \63492 , \63482 , \63491 );
or \U$63150 ( \63493 , \63484 , \63489 );
nand \U$63151 ( \63494 , \63492 , \63493 );
and \U$63152 ( \63495 , \50157 , \63494 );
nor \U$63153 ( \63496 , \50156 , \63495 );
or \U$63154 ( \63497 , \49735 , \63496 );
nand \U$63155 ( \63498 , \49734 , \63497 );
and \U$63156 ( \63499 , \49281 , \63498 );
nor \U$63157 ( \63500 , \49280 , \63499 );
not \U$63158 ( \63501 , \63500 );
xor \U$63159 ( \63502 , \48817 , \48826 );
and \U$63160 ( \63503 , \63502 , \48837 );
and \U$63161 ( \63504 , \48817 , \48826 );
or \U$63162 ( \63505 , \63503 , \63504 );
not \U$63163 ( \63506 , \47864 );
not \U$63164 ( \63507 , \48363 );
not \U$63165 ( \63508 , \47859 );
and \U$63166 ( \63509 , \63507 , \63508 );
and \U$63167 ( \63510 , \48363 , \47859 );
nor \U$63168 ( \63511 , \63509 , \63510 );
not \U$63169 ( \63512 , \63511 );
or \U$63170 ( \63513 , \63506 , \63512 );
or \U$63171 ( \63514 , \63511 , \47864 );
nand \U$63172 ( \63515 , \63513 , \63514 );
xor \U$63173 ( \63516 , \63505 , \63515 );
and \U$63174 ( \63517 , \63501 , \63516 );
and \U$63175 ( \63518 , \63505 , \63515 );
nor \U$63176 ( \63519 , \63517 , \63518 );
and \U$63177 ( \63520 , \48366 , \63519 );
and \U$63178 ( \63521 , \47849 , \48365 );
nor \U$63179 ( \63522 , \63520 , \63521 );
or \U$63180 ( \63523 , \47844 , \47358 );
not \U$63181 ( \63524 , \47358 );
not \U$63182 ( \63525 , \47844 );
or \U$63183 ( \63526 , \63524 , \63525 );
nand \U$63184 ( \63527 , \63526 , \47343 );
nand \U$63185 ( \63528 , \63523 , \63527 );
xor \U$63186 ( \63529 , \46797 , \46799 );
xor \U$63187 ( \63530 , \63529 , \46840 );
and \U$63188 ( \63531 , \47309 , \63530 );
xor \U$63189 ( \63532 , \46797 , \46799 );
xor \U$63190 ( \63533 , \63532 , \46840 );
and \U$63191 ( \63534 , \47341 , \63533 );
and \U$63192 ( \63535 , \47309 , \47341 );
or \U$63193 ( \63536 , \63531 , \63534 , \63535 );
xor \U$63194 ( \63537 , \47325 , \47329 );
and \U$63195 ( \63538 , \63537 , \47338 );
and \U$63196 ( \63539 , \47325 , \47329 );
or \U$63197 ( \63540 , \63538 , \63539 );
xor \U$63198 ( \63541 , \47311 , \47313 );
and \U$63199 ( \63542 , \63541 , \47318 );
and \U$63200 ( \63543 , \47311 , \47313 );
or \U$63201 ( \63544 , \63542 , \63543 );
xor \U$63202 ( \63545 , \63540 , \63544 );
xor \U$63203 ( \63546 , \45225 , \45227 );
xor \U$63204 ( \63547 , \63546 , \45230 );
xor \U$63205 ( \63548 , \46027 , \46034 );
xor \U$63206 ( \63549 , \63547 , \63548 );
xor \U$63207 ( \63550 , \63545 , \63549 );
xor \U$63208 ( \63551 , \63536 , \63550 );
xor \U$63209 ( \63552 , \46797 , \46799 );
and \U$63210 ( \63553 , \63552 , \46840 );
and \U$63211 ( \63554 , \46797 , \46799 );
or \U$63212 ( \63555 , \63553 , \63554 );
xor \U$63213 ( \63556 , \45678 , \46004 );
xor \U$63214 ( \63557 , \63556 , \46019 );
xor \U$63215 ( \63558 , \63555 , \63557 );
xor \U$63216 ( \63559 , \47311 , \47313 );
xor \U$63217 ( \63560 , \63559 , \47318 );
and \U$63218 ( \63561 , \47321 , \63560 );
xor \U$63219 ( \63562 , \47311 , \47313 );
xor \U$63220 ( \63563 , \63562 , \47318 );
and \U$63221 ( \63564 , \47339 , \63563 );
and \U$63222 ( \63565 , \47321 , \47339 );
or \U$63223 ( \63566 , \63561 , \63564 , \63565 );
xor \U$63224 ( \63567 , \63558 , \63566 );
xor \U$63225 ( \63568 , \63551 , \63567 );
xor \U$63226 ( \63569 , \63528 , \63568 );
and \U$63227 ( \63570 , \63522 , \63569 );
and \U$63228 ( \63571 , \63528 , \63568 );
nor \U$63229 ( \63572 , \63570 , \63571 );
not \U$63230 ( \63573 , \63572 );
xor \U$63231 ( \63574 , \63555 , \63557 );
and \U$63232 ( \63575 , \63574 , \63566 );
and \U$63233 ( \63576 , \63555 , \63557 );
or \U$63234 ( \63577 , \63575 , \63576 );
not \U$63235 ( \63578 , \63577 );
xor \U$63236 ( \63579 , \63540 , \63544 );
and \U$63237 ( \63580 , \63579 , \63549 );
and \U$63238 ( \63581 , \63540 , \63544 );
or \U$63239 ( \63582 , \63580 , \63581 );
xor \U$63240 ( \63583 , \46022 , \46024 );
xor \U$63241 ( \63584 , \63583 , \46039 );
xnor \U$63242 ( \63585 , \63582 , \63584 );
not \U$63243 ( \63586 , \63585 );
xor \U$63244 ( \63587 , \45598 , \45600 );
xor \U$63245 ( \63588 , \63587 , \45605 );
xor \U$63246 ( \63589 , \45635 , \45640 );
xor \U$63247 ( \63590 , \63588 , \63589 );
not \U$63248 ( \63591 , \63590 );
and \U$63249 ( \63592 , \63586 , \63591 );
and \U$63250 ( \63593 , \63585 , \63590 );
nor \U$63251 ( \63594 , \63592 , \63593 );
not \U$63252 ( \63595 , \63594 );
or \U$63253 ( \63596 , \63578 , \63595 );
or \U$63254 ( \63597 , \63594 , \63577 );
nand \U$63255 ( \63598 , \63596 , \63597 );
xor \U$63256 ( \63599 , \63536 , \63550 );
and \U$63257 ( \63600 , \63599 , \63567 );
and \U$63258 ( \63601 , \63536 , \63550 );
or \U$63259 ( \63602 , \63600 , \63601 );
xor \U$63260 ( \63603 , \63598 , \63602 );
and \U$63261 ( \63604 , \63573 , \63603 );
and \U$63262 ( \63605 , \63598 , \63602 );
nor \U$63263 ( \63606 , \63604 , \63605 );
not \U$63264 ( \63607 , \63594 );
nand \U$63265 ( \63608 , \63607 , \63577 );
not \U$63266 ( \63609 , \63590 );
not \U$63267 ( \63610 , \63584 );
or \U$63268 ( \63611 , \63609 , \63610 );
or \U$63269 ( \63612 , \63584 , \63590 );
nand \U$63270 ( \63613 , \63612 , \63582 );
nand \U$63271 ( \63614 , \63611 , \63613 );
xor \U$63272 ( \63615 , \45596 , \45608 );
xor \U$63273 ( \63616 , \63615 , \45613 );
xor \U$63274 ( \63617 , \63614 , \63616 );
xor \U$63275 ( \63618 , \45633 , \45645 );
xor \U$63276 ( \63619 , \63618 , \46042 );
xor \U$63277 ( \63620 , \63617 , \63619 );
and \U$63278 ( \63621 , \63608 , \63620 );
not \U$63279 ( \63622 , \63608 );
not \U$63280 ( \63623 , \63620 );
and \U$63281 ( \63624 , \63622 , \63623 );
nor \U$63282 ( \63625 , \63621 , \63624 );
or \U$63283 ( \63626 , \63606 , \63625 );
or \U$63284 ( \63627 , \63608 , \63623 );
nand \U$63285 ( \63628 , \63626 , \63627 );
not \U$63286 ( \63629 , \46045 );
not \U$63287 ( \63630 , \46048 );
or \U$63288 ( \63631 , \63629 , \63630 );
or \U$63289 ( \63632 , \46048 , \46045 );
nand \U$63290 ( \63633 , \63631 , \63632 );
xor \U$63291 ( \63634 , \63614 , \63616 );
and \U$63292 ( \63635 , \63634 , \63619 );
and \U$63293 ( \63636 , \63614 , \63616 );
or \U$63294 ( \63637 , \63635 , \63636 );
xor \U$63295 ( \63638 , \63633 , \63637 );
and \U$63296 ( \63639 , \63628 , \63638 );
and \U$63297 ( \63640 , \63633 , \63637 );
nor \U$63298 ( \63641 , \63639 , \63640 );
or \U$63299 ( \63642 , \46055 , \63641 );
nand \U$63300 ( \63643 , \46050 , \63642 );
and \U$63301 ( \63644 , \45629 , \63643 );
nor \U$63302 ( \63645 , \45628 , \63644 );
xnor \U$63303 ( \63646 , \45205 , \45215 );
or \U$63304 ( \63647 , \63645 , \63646 );
nand \U$63305 ( \63648 , \45217 , \63647 );
xor \U$63306 ( \63649 , \44388 , \44390 );
and \U$63307 ( \63650 , \45210 , \45214 );
xor \U$63308 ( \63651 , \63649 , \63650 );
and \U$63309 ( \63652 , \63648 , \63651 );
and \U$63310 ( \63653 , \63649 , \63650 );
nor \U$63311 ( \63654 , \63652 , \63653 );
xnor \U$63312 ( \63655 , \44391 , \44393 );
or \U$63313 ( \63656 , \63654 , \63655 );
nand \U$63314 ( \63657 , \44395 , \63656 );
and \U$63315 ( \63658 , \43999 , \63657 );
nor \U$63316 ( \63659 , \43998 , \63658 );
xnor \U$63317 ( \63660 , \43579 , \43587 );
or \U$63318 ( \63661 , \63659 , \63660 );
nand \U$63319 ( \63662 , \43589 , \63661 );
and \U$63320 ( \63663 , \43584 , \43586 );
xor \U$63321 ( \63664 , \42819 , \42829 );
xor \U$63322 ( \63665 , \63663 , \63664 );
and \U$63323 ( \63666 , \63662 , \63665 );
and \U$63324 ( \63667 , \63663 , \63664 );
nor \U$63325 ( \63668 , \63666 , \63667 );
xnor \U$63326 ( \63669 , \42830 , \42838 );
or \U$63327 ( \63670 , \63668 , \63669 );
nand \U$63328 ( \63671 , \42840 , \63670 );
not \U$63329 ( \63672 , \42094 );
not \U$63330 ( \63673 , \41733 );
or \U$63331 ( \63674 , \63672 , \63673 );
or \U$63332 ( \63675 , \41733 , \42094 );
nand \U$63333 ( \63676 , \63674 , \63675 );
and \U$63334 ( \63677 , \42835 , \42837 );
xor \U$63335 ( \63678 , \63676 , \63677 );
and \U$63336 ( \63679 , \63671 , \63678 );
and \U$63337 ( \63680 , \63676 , \63677 );
nor \U$63338 ( \63681 , \63679 , \63680 );
or \U$63339 ( \63682 , \42097 , \63681 );
nand \U$63340 ( \63683 , \42096 , \63682 );
and \U$63341 ( \63684 , \41718 , \63683 );
nor \U$63342 ( \63685 , \41717 , \63684 );
not \U$63343 ( \63686 , \41321 );
nand \U$63344 ( \63687 , \63686 , \41340 );
xor \U$63345 ( \63688 , \40571 , \40573 );
xor \U$63346 ( \63689 , \63688 , \40576 );
not \U$63347 ( \63690 , \63689 );
and \U$63348 ( \63691 , \41324 , \41332 );
not \U$63349 ( \63692 , \41324 );
not \U$63350 ( \63693 , \41332 );
and \U$63351 ( \63694 , \63692 , \63693 );
nor \U$63352 ( \63695 , \63694 , \41329 );
nor \U$63353 ( \63696 , \63691 , \63695 );
not \U$63354 ( \63697 , \63696 );
and \U$63355 ( \63698 , \63690 , \63697 );
and \U$63356 ( \63699 , \63689 , \63696 );
nor \U$63357 ( \63700 , \63698 , \63699 );
xnor \U$63358 ( \63701 , \63687 , \63700 );
or \U$63359 ( \63702 , \63685 , \63701 );
or \U$63360 ( \63703 , \63687 , \63700 );
nand \U$63361 ( \63704 , \63702 , \63703 );
not \U$63362 ( \63705 , \63689 );
nor \U$63363 ( \63706 , \63705 , \63696 );
xor \U$63364 ( \63707 , \40579 , \40581 );
xor \U$63365 ( \63708 , \63706 , \63707 );
and \U$63366 ( \63709 , \63704 , \63708 );
and \U$63367 ( \63710 , \63706 , \63707 );
nor \U$63368 ( \63711 , \63709 , \63710 );
xnor \U$63369 ( \63712 , \40204 , \40582 );
or \U$63370 ( \63713 , \63711 , \63712 );
nand \U$63371 ( \63714 , \40584 , \63713 );
and \U$63372 ( \63715 , \40203 , \63714 );
nor \U$63373 ( \63716 , \40202 , \63715 );
xnor \U$63374 ( \63717 , \39848 , \39853 );
or \U$63375 ( \63718 , \63716 , \63717 );
nand \U$63376 ( \63719 , \39855 , \63718 );
and \U$63377 ( \63720 , \39514 , \63719 );
nor \U$63378 ( \63721 , \39513 , \63720 );
not \U$63379 ( \63722 , \63721 );
xor \U$63380 ( \63723 , \39506 , \39508 );
and \U$63381 ( \63724 , \63723 , \39511 );
and \U$63382 ( \63725 , \39506 , \39508 );
or \U$63383 ( \63726 , \63724 , \63725 );
xor \U$63384 ( \63727 , \38625 , \38627 );
xor \U$63385 ( \63728 , \63727 , \38630 );
xor \U$63386 ( \63729 , \63726 , \63728 );
and \U$63387 ( \63730 , \63722 , \63729 );
and \U$63388 ( \63731 , \63726 , \63728 );
nor \U$63389 ( \63732 , \63730 , \63731 );
not \U$63390 ( \63733 , \63732 );
and \U$63391 ( \63734 , \38640 , \63733 );
nor \U$63392 ( \63735 , \38639 , \63734 );
or \U$63393 ( \63736 , \38344 , \63735 );
nand \U$63394 ( \63737 , \38339 , \63736 );
and \U$63395 ( \63738 , \38016 , \38061 );
xor \U$63396 ( \63739 , \38020 , \38038 );
and \U$63397 ( \63740 , \63739 , \38060 );
and \U$63398 ( \63741 , \38020 , \38038 );
or \U$63399 ( \63742 , \63740 , \63741 );
xor \U$63400 ( \63743 , \38047 , \38051 );
and \U$63401 ( \63744 , \63743 , \38059 );
and \U$63402 ( \63745 , \38047 , \38051 );
or \U$63403 ( \63746 , \63744 , \63745 );
xor \U$63404 ( \63747 , \37015 , \37020 );
xor \U$63405 ( \63748 , \63747 , \37053 );
xor \U$63406 ( \63749 , \63746 , \63748 );
xor \U$63407 ( \63750 , \38028 , \38032 );
and \U$63408 ( \63751 , \63750 , \38037 );
and \U$63409 ( \63752 , \38028 , \38032 );
or \U$63410 ( \63753 , \63751 , \63752 );
xor \U$63411 ( \63754 , \36914 , \36935 );
xor \U$63412 ( \63755 , \63754 , \37012 );
and \U$63413 ( \63756 , \38055 , \63755 );
xor \U$63414 ( \63757 , \36914 , \36935 );
xor \U$63415 ( \63758 , \63757 , \37012 );
and \U$63416 ( \63759 , \38057 , \63758 );
and \U$63417 ( \63760 , \38055 , \38057 );
or \U$63418 ( \63761 , \63756 , \63759 , \63760 );
xor \U$63419 ( \63762 , \63753 , \63761 );
xor \U$63420 ( \63763 , \37063 , \37068 );
xor \U$63421 ( \63764 , \63763 , \37079 );
xor \U$63422 ( \63765 , \63762 , \63764 );
xor \U$63423 ( \63766 , \63749 , \63765 );
xor \U$63424 ( \63767 , \63742 , \63766 );
xor \U$63425 ( \63768 , \63738 , \63767 );
and \U$63426 ( \63769 , \63737 , \63768 );
and \U$63427 ( \63770 , \63738 , \63767 );
nor \U$63428 ( \63771 , \63769 , \63770 );
nand \U$63429 ( \63772 , \63742 , \63766 );
xor \U$63430 ( \63773 , \63753 , \63761 );
and \U$63431 ( \63774 , \63773 , \63764 );
and \U$63432 ( \63775 , \63753 , \63761 );
or \U$63433 ( \63776 , \63774 , \63775 );
not \U$63434 ( \63777 , \63776 );
xor \U$63435 ( \63778 , \36717 , \36723 );
xor \U$63436 ( \63779 , \63778 , \36772 );
not \U$63437 ( \63780 , \63779 );
and \U$63438 ( \63781 , \63777 , \63780 );
and \U$63439 ( \63782 , \63776 , \63779 );
nor \U$63440 ( \63783 , \63781 , \63782 );
not \U$63441 ( \63784 , \63783 );
xor \U$63442 ( \63785 , \36830 , \37056 );
xor \U$63443 ( \63786 , \63785 , \37082 );
not \U$63444 ( \63787 , \63786 );
and \U$63445 ( \63788 , \63784 , \63787 );
and \U$63446 ( \63789 , \63783 , \63786 );
nor \U$63447 ( \63790 , \63788 , \63789 );
not \U$63448 ( \63791 , \63790 );
xor \U$63449 ( \63792 , \63746 , \63748 );
and \U$63450 ( \63793 , \63792 , \63765 );
and \U$63451 ( \63794 , \63746 , \63748 );
or \U$63452 ( \63795 , \63793 , \63794 );
not \U$63453 ( \63796 , \63795 );
and \U$63454 ( \63797 , \63791 , \63796 );
and \U$63455 ( \63798 , \63790 , \63795 );
nor \U$63456 ( \63799 , \63797 , \63798 );
xnor \U$63457 ( \63800 , \63772 , \63799 );
or \U$63458 ( \63801 , \63771 , \63800 );
or \U$63459 ( \63802 , \63772 , \63799 );
nand \U$63460 ( \63803 , \63801 , \63802 );
not \U$63461 ( \63804 , \63795 );
nor \U$63462 ( \63805 , \63804 , \63790 );
not \U$63463 ( \63806 , \63786 );
or \U$63464 ( \63807 , \63806 , \63779 );
not \U$63465 ( \63808 , \63779 );
not \U$63466 ( \63809 , \63806 );
or \U$63467 ( \63810 , \63808 , \63809 );
nand \U$63468 ( \63811 , \63810 , \63776 );
nand \U$63469 ( \63812 , \63807 , \63811 );
not \U$63470 ( \63813 , \63812 );
xor \U$63471 ( \63814 , \36809 , \36819 );
xor \U$63472 ( \63815 , \63814 , \37085 );
not \U$63473 ( \63816 , \63815 );
or \U$63474 ( \63817 , \63813 , \63816 );
or \U$63475 ( \63818 , \63815 , \63812 );
nand \U$63476 ( \63819 , \63817 , \63818 );
xor \U$63477 ( \63820 , \63805 , \63819 );
and \U$63478 ( \63821 , \63803 , \63820 );
and \U$63479 ( \63822 , \63805 , \63819 );
nor \U$63480 ( \63823 , \63821 , \63822 );
not \U$63481 ( \63824 , \63815 );
nand \U$63482 ( \63825 , \63824 , \63812 );
not \U$63483 ( \63826 , \36802 );
not \U$63484 ( \63827 , \37088 );
and \U$63485 ( \63828 , \63826 , \63827 );
and \U$63486 ( \63829 , \36802 , \37088 );
nor \U$63487 ( \63830 , \63828 , \63829 );
xnor \U$63488 ( \63831 , \63825 , \63830 );
or \U$63489 ( \63832 , \63823 , \63831 );
or \U$63490 ( \63833 , \63825 , \63830 );
nand \U$63491 ( \63834 , \63832 , \63833 );
and \U$63492 ( \63835 , \37091 , \63834 );
nor \U$63493 ( \63836 , \37090 , \63835 );
and \U$63494 ( \63837 , \36799 , \63836 );
and \U$63495 ( \63838 , \36509 , \36798 );
nor \U$63496 ( \63839 , \63837 , \63838 );
and \U$63497 ( \63840 , \36504 , \63839 );
nor \U$63498 ( \63841 , \36503 , \63840 );
not \U$63499 ( \63842 , \63841 );
and \U$63500 ( \63843 , \36206 , \36225 );
xor \U$63501 ( \63844 , \36207 , \36217 );
and \U$63502 ( \63845 , \63844 , \36224 );
and \U$63503 ( \63846 , \36207 , \36217 );
nor \U$63504 ( \63847 , \63845 , \63846 );
not \U$63505 ( \63848 , \63847 );
not \U$63506 ( \63849 , \35487 );
not \U$63507 ( \63850 , \35497 );
not \U$63508 ( \63851 , \35729 );
or \U$63509 ( \63852 , \63850 , \63851 );
or \U$63510 ( \63853 , \35729 , \35497 );
nand \U$63511 ( \63854 , \63852 , \63853 );
not \U$63512 ( \63855 , \63854 );
or \U$63513 ( \63856 , \63849 , \63855 );
or \U$63514 ( \63857 , \63854 , \35487 );
nand \U$63515 ( \63858 , \63856 , \63857 );
not \U$63516 ( \63859 , \63858 );
or \U$63517 ( \63860 , \63848 , \63859 );
or \U$63518 ( \63861 , \63858 , \63847 );
nand \U$63519 ( \63862 , \63860 , \63861 );
xor \U$63520 ( \63863 , \63843 , \63862 );
and \U$63521 ( \63864 , \63842 , \63863 );
and \U$63522 ( \63865 , \63862 , \63843 );
nor \U$63523 ( \63866 , \63864 , \63865 );
not \U$63524 ( \63867 , \63847 );
nand \U$63525 ( \63868 , \63867 , \63858 );
not \U$63526 ( \63869 , \35484 );
not \U$63527 ( \63870 , \35731 );
and \U$63528 ( \63871 , \63869 , \63870 );
and \U$63529 ( \63872 , \35484 , \35731 );
nor \U$63530 ( \63873 , \63871 , \63872 );
xnor \U$63531 ( \63874 , \63868 , \63873 );
or \U$63532 ( \63875 , \63866 , \63874 );
or \U$63533 ( \63876 , \63868 , \63873 );
nand \U$63534 ( \63877 , \63875 , \63876 );
and \U$63535 ( \63878 , \35734 , \63877 );
nor \U$63536 ( \63879 , \35733 , \63878 );
xnor \U$63537 ( \63880 , \35463 , \35445 );
or \U$63538 ( \63881 , \63879 , \63880 );
nand \U$63539 ( \63882 , \35464 , \63881 );
not \U$63540 ( \63883 , \34778 );
not \U$63541 ( \63884 , \34781 );
or \U$63542 ( \63885 , \63883 , \63884 );
or \U$63543 ( \63886 , \34781 , \34778 );
nand \U$63544 ( \63887 , \63885 , \63886 );
not \U$63545 ( \63888 , \35459 );
or \U$63546 ( \63889 , \35447 , \63888 );
not \U$63547 ( \63890 , \63888 );
not \U$63548 ( \63891 , \35447 );
or \U$63549 ( \63892 , \63890 , \63891 );
nand \U$63550 ( \63893 , \63892 , \35452 );
nand \U$63551 ( \63894 , \63889 , \63893 );
xor \U$63552 ( \63895 , \63887 , \63894 );
and \U$63553 ( \63896 , \63882 , \63895 );
and \U$63554 ( \63897 , \63887 , \63894 );
nor \U$63555 ( \63898 , \63896 , \63897 );
and \U$63556 ( \63899 , \34788 , \63898 );
and \U$63557 ( \63900 , \34782 , \34787 );
nor \U$63558 ( \63901 , \63899 , \63900 );
and \U$63559 ( \63902 , \34593 , \63901 );
nor \U$63560 ( \63903 , \34592 , \63902 );
or \U$63561 ( \63904 , \34409 , \63903 );
nand \U$63562 ( \63905 , \34408 , \63904 );
not \U$63563 ( \63906 , \34046 );
nor \U$63564 ( \63907 , \63906 , \34215 );
not \U$63565 ( \63908 , \34008 );
not \U$63566 ( \63909 , \34019 );
or \U$63567 ( \63910 , \63908 , \63909 );
or \U$63568 ( \63911 , \34019 , \34008 );
nand \U$63569 ( \63912 , \63910 , \63911 );
xor \U$63570 ( \63913 , \63907 , \63912 );
and \U$63571 ( \63914 , \63905 , \63913 );
and \U$63572 ( \63915 , \63907 , \63912 );
nor \U$63573 ( \63916 , \63914 , \63915 );
and \U$63574 ( \63917 , \34036 , \63916 );
and \U$63575 ( \63918 , \34020 , \34035 );
nor \U$63576 ( \63919 , \63917 , \63918 );
not \U$63577 ( \63920 , \33657 );
not \U$63578 ( \63921 , \33497 );
or \U$63579 ( \63922 , \63920 , \63921 );
or \U$63580 ( \63923 , \33497 , \33657 );
nand \U$63581 ( \63924 , \63922 , \63923 );
not \U$63582 ( \63925 , \34031 );
nor \U$63583 ( \63926 , \63925 , \34026 );
xor \U$63584 ( \63927 , \63924 , \63926 );
and \U$63585 ( \63928 , \63919 , \63927 );
and \U$63586 ( \63929 , \63924 , \63926 );
nor \U$63587 ( \63930 , \63928 , \63929 );
and \U$63588 ( \63931 , \33689 , \63930 );
and \U$63589 ( \63932 , \33658 , \33688 );
nor \U$63590 ( \63933 , \63931 , \63932 );
xor \U$63591 ( \63934 , \33678 , \33680 );
and \U$63592 ( \63935 , \63934 , \33683 );
and \U$63593 ( \63936 , \33678 , \33680 );
or \U$63594 ( \63937 , \63935 , \63936 );
not \U$63595 ( \63938 , \63937 );
not \U$63596 ( \63939 , \33054 );
not \U$63597 ( \63940 , \33158 );
not \U$63598 ( \63941 , \33056 );
and \U$63599 ( \63942 , \63940 , \63941 );
and \U$63600 ( \63943 , \33158 , \33056 );
nor \U$63601 ( \63944 , \63942 , \63943 );
not \U$63602 ( \63945 , \63944 );
or \U$63603 ( \63946 , \63939 , \63945 );
or \U$63604 ( \63947 , \63944 , \33054 );
nand \U$63605 ( \63948 , \63946 , \63947 );
not \U$63606 ( \63949 , \63948 );
or \U$63607 ( \63950 , \63938 , \63949 );
or \U$63608 ( \63951 , \63937 , \63948 );
nand \U$63609 ( \63952 , \63950 , \63951 );
or \U$63610 ( \63953 , \33684 , \33662 );
not \U$63611 ( \63954 , \33662 );
not \U$63612 ( \63955 , \33684 );
or \U$63613 ( \63956 , \63954 , \63955 );
nand \U$63614 ( \63957 , \63956 , \33669 );
nand \U$63615 ( \63958 , \63953 , \63957 );
xor \U$63616 ( \63959 , \63952 , \63958 );
and \U$63617 ( \63960 , \63933 , \63959 );
and \U$63618 ( \63961 , \63952 , \63958 );
nor \U$63619 ( \63962 , \63960 , \63961 );
not \U$63620 ( \63963 , \63937 );
nand \U$63621 ( \63964 , \63963 , \63948 );
not \U$63622 ( \63965 , \33051 );
not \U$63623 ( \63966 , \33160 );
and \U$63624 ( \63967 , \63965 , \63966 );
and \U$63625 ( \63968 , \33051 , \33160 );
nor \U$63626 ( \63969 , \63967 , \63968 );
xnor \U$63627 ( \63970 , \63964 , \63969 );
or \U$63628 ( \63971 , \63962 , \63970 );
or \U$63629 ( \63972 , \63964 , \63969 );
nand \U$63630 ( \63973 , \63971 , \63972 );
and \U$63631 ( \63974 , \33163 , \63973 );
nor \U$63632 ( \63975 , \33162 , \63974 );
not \U$63633 ( \63976 , \33045 );
nand \U$63634 ( \63977 , \63976 , \33034 );
xor \U$63635 ( \63978 , \33039 , \33041 );
and \U$63636 ( \63979 , \63978 , \33044 );
and \U$63637 ( \63980 , \33039 , \33041 );
or \U$63638 ( \63981 , \63979 , \63980 );
xor \U$63639 ( \63982 , \970 , \1010 );
xor \U$63640 ( \63983 , \63982 , \1059 );
xnor \U$63641 ( \63984 , \63981 , \63983 );
xnor \U$63642 ( \63985 , \63977 , \63984 );
or \U$63643 ( \63986 , \63975 , \63985 );
or \U$63644 ( \63987 , \63977 , \63984 );
or \U$63645 ( \63988 , \63981 , \63983 );
nand \U$63646 ( \63989 , \63986 , \63987 , \63988 );
not \U$63647 ( \63990 , \63989 );
or \U$63648 ( \63991 , \32834 , \63990 );
or \U$63649 ( \63992 , \63989 , \32833 );
nand \U$63650 ( \63993 , \63991 , \63992 );
not \U$63651 ( \63994 , \63993 );
xor \U$63652 ( \63995 , \1196 , \32716 );
xor \U$63653 ( \63996 , \63985 , \63975 );
xor \U$63654 ( \63997 , \63995 , \63996 );
xor \U$63655 ( \63998 , \63970 , \63962 );
xor \U$63656 ( \63999 , \32702 , \32686 );
or \U$63657 ( \64000 , \63998 , \63999 );
xnor \U$63658 ( \64001 , \32683 , \32649 );
xnor \U$63659 ( \64002 , \63959 , \63933 );
or \U$63660 ( \64003 , \64001 , \64002 );
not \U$63661 ( \64004 , \64001 );
not \U$63662 ( \64005 , \64002 );
or \U$63663 ( \64006 , \64004 , \64005 );
xor \U$63664 ( \64007 , \63927 , \63919 );
xor \U$63665 ( \64008 , \2026 , \32593 );
and \U$63666 ( \64009 , \64007 , \64008 );
or \U$63667 ( \64010 , \64007 , \64008 );
xor \U$63668 ( \64011 , \63913 , \63905 );
xor \U$63669 ( \64012 , \32579 , \32563 );
and \U$63670 ( \64013 , \64011 , \64012 );
not \U$63671 ( \64014 , \64011 );
not \U$63672 ( \64015 , \64012 );
and \U$63673 ( \64016 , \64014 , \64015 );
xor \U$63674 ( \64017 , \34409 , \63903 );
not \U$63675 ( \64018 , \64017 );
xor \U$63676 ( \64019 , \32560 , \32528 );
not \U$63677 ( \64020 , \64019 );
and \U$63678 ( \64021 , \64018 , \64020 );
xnor \U$63679 ( \64022 , \34593 , \63901 );
xnor \U$63680 ( \64023 , \32525 , \32485 );
and \U$63681 ( \64024 , \64022 , \64023 );
nor \U$63682 ( \64025 , \64021 , \64024 );
xor \U$63683 ( \64026 , \34782 , \34787 );
xor \U$63684 ( \64027 , \64026 , \63898 );
xor \U$63685 ( \64028 , \2848 , \2911 );
xor \U$63686 ( \64029 , \64028 , \32482 );
or \U$63687 ( \64030 , \64027 , \64029 );
not \U$63688 ( \64031 , \64029 );
not \U$63689 ( \64032 , \64027 );
or \U$63690 ( \64033 , \64031 , \64032 );
xor \U$63691 ( \64034 , \63895 , \63882 );
xor \U$63692 ( \64035 , \3125 , \32480 );
or \U$63693 ( \64036 , \64034 , \64035 );
nand \U$63694 ( \64037 , \64033 , \64036 );
and \U$63695 ( \64038 , \64034 , \64035 );
xnor \U$63696 ( \64039 , \35734 , \63877 );
xnor \U$63697 ( \64040 , \3862 , \32458 );
or \U$63698 ( \64041 , \64039 , \64040 );
not \U$63699 ( \64042 , \64040 );
not \U$63700 ( \64043 , \64039 );
or \U$63701 ( \64044 , \64042 , \64043 );
xnor \U$63702 ( \64045 , \36504 , \63839 );
xnor \U$63703 ( \64046 , \32449 , \32445 );
or \U$63704 ( \64047 , \64045 , \64046 );
not \U$63705 ( \64048 , \64046 );
not \U$63706 ( \64049 , \64045 );
or \U$63707 ( \64050 , \64048 , \64049 );
xor \U$63708 ( \64051 , \37091 , \63834 );
xor \U$63709 ( \64052 , \5249 , \32419 );
and \U$63710 ( \64053 , \64051 , \64052 );
or \U$63711 ( \64054 , \64051 , \64052 );
xor \U$63712 ( \64055 , \63831 , \63823 );
xor \U$63713 ( \64056 , \5517 , \32417 );
xor \U$63714 ( \64057 , \64055 , \64056 );
xor \U$63715 ( \64058 , \63800 , \63771 );
xor \U$63716 ( \64059 , \6067 , \32404 );
and \U$63717 ( \64060 , \64058 , \64059 );
or \U$63718 ( \64061 , \64058 , \64059 );
xnor \U$63719 ( \64062 , \63768 , \63737 );
xnor \U$63720 ( \64063 , \6362 , \32402 );
or \U$63721 ( \64064 , \64062 , \64063 );
not \U$63722 ( \64065 , \64063 );
not \U$63723 ( \64066 , \64062 );
or \U$63724 ( \64067 , \64065 , \64066 );
and \U$63725 ( \64068 , \63729 , \63722 );
not \U$63726 ( \64069 , \63729 );
and \U$63727 ( \64070 , \64069 , \63721 );
nor \U$63728 ( \64071 , \64068 , \64070 );
xor \U$63729 ( \64072 , \32369 , \32368 );
xor \U$63730 ( \64073 , \64071 , \64072 );
xor \U$63731 ( \64074 , \39514 , \63719 );
xor \U$63732 ( \64075 , \32365 , \32356 );
xor \U$63733 ( \64076 , \64074 , \64075 );
xor \U$63734 ( \64077 , \63717 , \63716 );
xor \U$63735 ( \64078 , \8333 , \32354 );
xor \U$63736 ( \64079 , \64077 , \64078 );
xor \U$63737 ( \64080 , \63708 , \63704 );
xor \U$63738 ( \64081 , \9490 , \32339 );
xor \U$63739 ( \64082 , \64080 , \64081 );
xor \U$63740 ( \64083 , \63701 , \63685 );
xor \U$63741 ( \64084 , \32336 , \32328 );
xor \U$63742 ( \64085 , \64083 , \64084 );
xor \U$63743 ( \64086 , \63678 , \63671 );
xor \U$63744 ( \64087 , \32261 , \32222 );
xor \U$63745 ( \64088 , \64086 , \64087 );
xor \U$63746 ( \64089 , \63660 , \63659 );
xor \U$63747 ( \64090 , \32211 , \32210 );
xor \U$63748 ( \64091 , \64089 , \64090 );
xor \U$63749 ( \64092 , \43999 , \63657 );
xor \U$63750 ( \64093 , \32207 , \32204 );
xor \U$63751 ( \64094 , \64092 , \64093 );
xor \U$63752 ( \64095 , \63655 , \63654 );
xor \U$63753 ( \64096 , \32202 , \32201 );
xor \U$63754 ( \64097 , \64095 , \64096 );
xor \U$63755 ( \64098 , \63638 , \63628 );
xor \U$63756 ( \64099 , \15144 , \32181 );
xor \U$63757 ( \64100 , \64098 , \64099 );
xor \U$63758 ( \64101 , \63625 , \63606 );
xor \U$63759 ( \64102 , \15620 , \32179 );
xor \U$63760 ( \64103 , \64101 , \64102 );
not \U$63761 ( \64104 , \63603 );
not \U$63762 ( \64105 , \63572 );
or \U$63763 ( \64106 , \64104 , \64105 );
or \U$63764 ( \64107 , \63572 , \63603 );
nand \U$63765 ( \64108 , \64106 , \64107 );
xor \U$63766 ( \64109 , \32176 , \32166 );
xor \U$63767 ( \64110 , \64108 , \64109 );
xor \U$63768 ( \64111 , \63569 , \63522 );
xor \U$63769 ( \64112 , \32164 , \32163 );
xor \U$63770 ( \64113 , \64111 , \64112 );
not \U$63771 ( \64114 , \63516 );
not \U$63772 ( \64115 , \63500 );
or \U$63773 ( \64116 , \64114 , \64115 );
or \U$63774 ( \64117 , \63500 , \63516 );
nand \U$63775 ( \64118 , \64116 , \64117 );
xor \U$63776 ( \64119 , \32148 , \32126 );
and \U$63777 ( \64120 , \64118 , \64119 );
or \U$63778 ( \64121 , \64118 , \64119 );
xor \U$63779 ( \64122 , \50157 , \63494 );
xor \U$63780 ( \64123 , \32104 , \32073 );
xor \U$63781 ( \64124 , \64122 , \64123 );
xor \U$63782 ( \64125 , \63491 , \63482 );
xor \U$63783 ( \64126 , \32069 , \32031 );
xor \U$63784 ( \64127 , \64125 , \64126 );
and \U$63785 ( \64128 , \51044 , \63480 );
not \U$63786 ( \64129 , \51044 );
and \U$63787 ( \64130 , \64129 , \63479 );
nor \U$63788 ( \64131 , \64128 , \64130 );
xor \U$63789 ( \64132 , \19704 , \32029 );
xor \U$63790 ( \64133 , \64131 , \64132 );
xor \U$63791 ( \64134 , \63476 , \63471 );
xor \U$63792 ( \64135 , \20113 , \32027 );
xor \U$63793 ( \64136 , \64134 , \64135 );
xor \U$63794 ( \64137 , \52288 , \63466 );
xor \U$63795 ( \64138 , \32013 , \31997 );
and \U$63796 ( \64139 , \64137 , \64138 );
xor \U$63797 ( \64140 , \52715 , \63464 );
xor \U$63798 ( \64141 , \31994 , \31962 );
xor \U$63799 ( \64142 , \64140 , \64141 );
xor \U$63800 ( \64143 , \63461 , \63453 );
xor \U$63801 ( \64144 , \31959 , \31891 );
xor \U$63802 ( \64145 , \64143 , \64144 );
xor \U$63803 ( \64146 , \63450 , \63436 );
xor \U$63804 ( \64147 , \31888 , \31827 );
xor \U$63805 ( \64148 , \64146 , \64147 );
xor \U$63806 ( \64149 , \53527 , \63434 );
xor \U$63807 ( \64150 , \21969 , \31825 );
xor \U$63808 ( \64151 , \64149 , \64150 );
xor \U$63809 ( \64152 , \63431 , \63421 );
xor \U$63810 ( \64153 , \22343 , \31823 );
xor \U$63811 ( \64154 , \64152 , \64153 );
xor \U$63812 ( \64155 , \63418 , \63396 );
xor \U$63813 ( \64156 , \22677 , \31821 );
xor \U$63814 ( \64157 , \64155 , \64156 );
xor \U$63815 ( \64158 , \54593 , \63394 );
xor \U$63816 ( \64159 , \31818 , \31809 );
xor \U$63817 ( \64160 , \64158 , \64159 );
xor \U$63818 ( \64161 , \54947 , \63392 );
xor \U$63819 ( \64162 , \23358 , \31807 );
xor \U$63820 ( \64163 , \64161 , \64162 );
xor \U$63821 ( \64164 , \63389 , \63378 );
xor \U$63822 ( \64165 , \23684 , \31805 );
xor \U$63823 ( \64166 , \64164 , \64165 );
xor \U$63824 ( \64167 , \63375 , \63356 );
xor \U$63825 ( \64168 , \31802 , \31791 );
xor \U$63826 ( \64169 , \64167 , \64168 );
xor \U$63827 ( \64170 , \63353 , \63298 );
xor \U$63828 ( \64171 , \24349 , \31789 );
xor \U$63829 ( \64172 , \64170 , \64171 );
xor \U$63830 ( \64173 , \56291 , \63296 );
xor \U$63831 ( \64174 , \31786 , \31775 );
xor \U$63832 ( \64175 , \64173 , \64174 );
xor \U$63833 ( \64176 , \24941 , \31773 );
xor \U$63834 ( \64177 , \63293 , \63276 );
xor \U$63835 ( \64178 , \64176 , \64177 );
xor \U$63836 ( \64179 , \56869 , \63274 );
xor \U$63837 ( \64180 , \31770 , \31759 );
xor \U$63838 ( \64181 , \64179 , \64180 );
xor \U$63839 ( \64182 , \63271 , \63260 );
xor \U$63840 ( \64183 , \25480 , \31757 );
xor \U$63841 ( \64184 , \64182 , \64183 );
xor \U$63842 ( \64185 , \63257 , \63241 );
xor \U$63843 ( \64186 , \31754 , \31743 );
xor \U$63844 ( \64187 , \64185 , \64186 );
xor \U$63845 ( \64188 , \26101 , \31741 );
xor \U$63846 ( \64189 , \57671 , \63239 );
xor \U$63847 ( \64190 , \64188 , \64189 );
xor \U$63848 ( \64191 , \31738 , \31729 );
xor \U$63849 ( \64192 , \63236 , \63231 );
xor \U$63850 ( \64193 , \64191 , \64192 );
xor \U$63851 ( \64194 , \58229 , \63229 );
xor \U$63852 ( \64195 , \31726 , \31704 );
xor \U$63853 ( \64196 , \64194 , \64195 );
xor \U$63854 ( \64197 , \31701 , \31670 );
xor \U$63855 ( \64198 , \58523 , \63227 );
xor \U$63856 ( \64199 , \64197 , \64198 );
xor \U$63857 ( \64200 , \63224 , \63216 );
xor \U$63858 ( \64201 , \31667 , \31605 );
xor \U$63859 ( \64202 , \64200 , \64201 );
xor \U$63860 ( \64203 , \31602 , \31528 );
xor \U$63861 ( \64204 , \58837 , \63214 );
xor \U$63862 ( \64205 , \64203 , \64204 );
xor \U$63863 ( \64206 , \31525 , \31437 );
xor \U$63864 ( \64207 , \59088 , \63212 );
xor \U$63865 ( \64208 , \64206 , \64207 );
xor \U$63866 ( \64209 , \59290 , \63210 );
xor \U$63867 ( \64210 , \31434 , \31242 );
xor \U$63868 ( \64211 , \64209 , \64210 );
xor \U$63869 ( \64212 , \31239 , \30957 );
xor \U$63870 ( \64213 , \63207 , \63196 );
xor \U$63871 ( \64214 , \64212 , \64213 );
xor \U$63872 ( \64215 , \30954 , \30697 );
xor \U$63873 ( \64216 , \59722 , \63194 );
xor \U$63874 ( \64217 , \64215 , \64216 );
xor \U$63875 ( \64218 , \30694 , \30431 );
xor \U$63876 ( \64219 , \59920 , \63192 );
xor \U$63877 ( \64220 , \64218 , \64219 );
xor \U$63878 ( \64221 , \63189 , \63180 );
xor \U$63879 ( \64222 , \27360 , \30429 );
xor \U$63880 ( \64223 , \64221 , \64222 );
xor \U$63881 ( \64224 , \27584 , \30427 );
xor \U$63882 ( \64225 , \60290 , \63178 );
xor \U$63883 ( \64226 , \64224 , \64225 );
xor \U$63884 ( \64227 , \30424 , \30409 );
xor \U$63885 ( \64228 , \60463 , \63176 );
xor \U$63886 ( \64229 , \64227 , \64228 );
xor \U$63887 ( \64230 , \63173 , \63162 );
xor \U$63888 ( \64231 , \27962 , \30407 );
xor \U$63889 ( \64232 , \64230 , \64231 );
xor \U$63890 ( \64233 , \63159 , \63140 );
xor \U$63891 ( \64234 , \30404 , \30393 );
xor \U$63892 ( \64235 , \64233 , \64234 );
xor \U$63893 ( \64236 , \61015 , \63138 );
xor \U$63894 ( \64237 , \30390 , \30374 );
xor \U$63895 ( \64238 , \64236 , \64237 );
xor \U$63896 ( \64239 , \28317 , \30372 );
xor \U$63897 ( \64240 , \61040 , \63136 );
xor \U$63898 ( \64241 , \64239 , \64240 );
xor \U$63899 ( \64242 , \61186 , \63134 );
xor \U$63900 ( \64243 , \30369 , \30357 );
xor \U$63901 ( \64244 , \64242 , \64243 );
xor \U$63902 ( \64245 , \30354 , \30328 );
xor \U$63903 ( \64246 , \61364 , \63132 );
xor \U$63904 ( \64247 , \64245 , \64246 );
xor \U$63905 ( \64248 , \63129 , \63118 );
xor \U$63906 ( \64249 , \30325 , \30289 );
xor \U$63907 ( \64250 , \64248 , \64249 );
xor \U$63908 ( \64251 , \63115 , \63096 );
xor \U$63909 ( \64252 , \28843 , \30287 );
xor \U$63910 ( \64253 , \64251 , \64252 );
xor \U$63911 ( \64254 , \30284 , \30275 );
xor \U$63912 ( \64255 , \61767 , \63094 );
xor \U$63913 ( \64256 , \64254 , \64255 );
xor \U$63914 ( \64257 , \30272 , \30242 );
xor \U$63915 ( \64258 , \63091 , \63082 );
xor \U$63916 ( \64259 , \64257 , \64258 );
xor \U$63917 ( \64260 , \63079 , \63061 );
xor \U$63918 ( \64261 , \30239 , \30216 );
xor \U$63919 ( \64262 , \64260 , \64261 );
xor \U$63920 ( \64263 , \30213 , \30165 );
xor \U$63921 ( \64264 , \62126 , \63059 );
xor \U$63922 ( \64265 , \64263 , \64264 );
xor \U$63923 ( \64266 , \29260 , \30163 );
xor \U$63924 ( \64267 , \62147 , \63057 );
xor \U$63925 ( \64268 , \64266 , \64267 );
xor \U$63926 ( \64269 , \30160 , \30148 );
xor \U$63927 ( \64270 , \62245 , \63055 );
xor \U$63928 ( \64271 , \64269 , \64270 );
xor \U$63929 ( \64272 , \30145 , \30121 );
xor \U$63930 ( \64273 , \63052 , \63039 );
xor \U$63931 ( \64274 , \64272 , \64273 );
xor \U$63932 ( \64275 , \30118 , \30083 );
xor \U$63933 ( \64276 , \63036 , \63009 );
xor \U$63934 ( \64277 , \64275 , \64276 );
xor \U$63935 ( \64278 , \29562 , \30081 );
xor \U$63936 ( \64279 , \62500 , \63007 );
xor \U$63937 ( \64280 , \64278 , \64279 );
xor \U$63938 ( \64281 , \30078 , \30069 );
xor \U$63939 ( \64282 , \63004 , \62999 );
xor \U$63940 ( \64283 , \64281 , \64282 );
xor \U$63941 ( \64284 , \30066 , \30050 );
xor \U$63942 ( \64285 , \62996 , \62980 );
xor \U$63943 ( \64286 , \64284 , \64285 );
xor \U$63944 ( \64287 , \29721 , \30048 );
xor \U$63945 ( \64288 , \62663 , \62978 );
xor \U$63946 ( \64289 , \64287 , \64288 );
xor \U$63947 ( \64290 , \30045 , \30032 );
xor \U$63948 ( \64291 , \62975 , \62965 );
xor \U$63949 ( \64292 , \64290 , \64291 );
xor \U$63950 ( \64293 , \29809 , \29834 );
xor \U$63951 ( \64294 , \64293 , \30029 );
xnor \U$63952 ( \64295 , \62962 , \62946 );
or \U$63953 ( \64296 , \64294 , \64295 );
xnor \U$63954 ( \64297 , \30026 , \30018 );
xor \U$63955 ( \64298 , \62747 , \62771 );
xor \U$63956 ( \64299 , \64298 , \62943 );
or \U$63957 ( \64300 , \64297 , \64299 );
xor \U$63958 ( \64301 , \29874 , \29891 );
xor \U$63959 ( \64302 , \64301 , \30015 );
xor \U$63960 ( \64303 , \62937 , \62932 );
xor \U$63961 ( \64304 , \30012 , \29999 );
and \U$63962 ( \64305 , \64303 , \64304 );
xor \U$63963 ( \64306 , \29916 , \29927 );
xor \U$63964 ( \64307 , \64306 , \29996 );
xor \U$63965 ( \64308 , \62841 , \62860 );
xor \U$63966 ( \64309 , \64308 , \62929 );
or \U$63967 ( \64310 , \64307 , \64309 );
not \U$63968 ( \64311 , \64309 );
not \U$63969 ( \64312 , \64307 );
or \U$63970 ( \64313 , \64311 , \64312 );
xnor \U$63971 ( \64314 , \29993 , \29951 );
xor \U$63972 ( \64315 , \29990 , \29966 );
xnor \U$63973 ( \64316 , \62920 , \62909 );
xor \U$63974 ( \64317 , \62911 , \62919 );
nor \U$63975 ( \64318 , \29985 , \62910 );
and \U$63976 ( \64319 , \64317 , \64318 );
and \U$63977 ( \64320 , \29984 , \29986 );
nor \U$63978 ( \64321 , \64317 , \64318 );
nor \U$63979 ( \64322 , \64320 , \64321 , \29987 );
nor \U$63980 ( \64323 , \64319 , \64322 );
or \U$63981 ( \64324 , \64316 , \64323 );
not \U$63982 ( \64325 , \64323 );
not \U$63983 ( \64326 , \64316 );
or \U$63984 ( \64327 , \64325 , \64326 );
xor \U$63985 ( \64328 , \29987 , \29976 );
nand \U$63986 ( \64329 , \64327 , \64328 );
nand \U$63987 ( \64330 , \64324 , \64329 );
or \U$63988 ( \64331 , \64315 , \64330 );
xor \U$63989 ( \64332 , \62923 , \62899 );
and \U$63990 ( \64333 , \64331 , \64332 );
and \U$63991 ( \64334 , \64330 , \64315 );
nor \U$63992 ( \64335 , \64333 , \64334 );
or \U$63993 ( \64336 , \64314 , \64335 );
not \U$63994 ( \64337 , \64335 );
not \U$63995 ( \64338 , \64314 );
or \U$63996 ( \64339 , \64337 , \64338 );
xor \U$63997 ( \64340 , \62926 , \62884 );
nand \U$63998 ( \64341 , \64339 , \64340 );
nand \U$63999 ( \64342 , \64336 , \64341 );
nand \U$64000 ( \64343 , \64313 , \64342 );
nand \U$64001 ( \64344 , \64310 , \64343 );
or \U$64002 ( \64345 , \64304 , \64303 );
and \U$64003 ( \64346 , \64344 , \64345 );
nor \U$64004 ( \64347 , \64305 , \64346 );
or \U$64005 ( \64348 , \64302 , \64347 );
nand \U$64006 ( \64349 , \64300 , \64348 );
and \U$64007 ( \64350 , \62941 , \62940 );
and \U$64008 ( \64351 , \64302 , \64347 );
nor \U$64009 ( \64352 , \64350 , \64351 , \62942 );
or \U$64010 ( \64353 , \64349 , \64352 );
and \U$64011 ( \64354 , \64297 , \64299 );
and \U$64012 ( \64355 , \64295 , \64294 );
nor \U$64013 ( \64356 , \64354 , \64355 );
nand \U$64014 ( \64357 , \64353 , \64356 );
nand \U$64015 ( \64358 , \64296 , \64357 );
and \U$64016 ( \64359 , \64292 , \64358 );
and \U$64017 ( \64360 , \64290 , \64291 );
or \U$64018 ( \64361 , \64359 , \64360 );
and \U$64019 ( \64362 , \64289 , \64361 );
and \U$64020 ( \64363 , \64287 , \64288 );
or \U$64021 ( \64364 , \64362 , \64363 );
and \U$64022 ( \64365 , \64286 , \64364 );
and \U$64023 ( \64366 , \64284 , \64285 );
or \U$64024 ( \64367 , \64365 , \64366 );
and \U$64025 ( \64368 , \64283 , \64367 );
and \U$64026 ( \64369 , \64281 , \64282 );
or \U$64027 ( \64370 , \64368 , \64369 );
and \U$64028 ( \64371 , \64280 , \64370 );
and \U$64029 ( \64372 , \64278 , \64279 );
or \U$64030 ( \64373 , \64371 , \64372 );
and \U$64031 ( \64374 , \64277 , \64373 );
and \U$64032 ( \64375 , \64275 , \64276 );
or \U$64033 ( \64376 , \64374 , \64375 );
and \U$64034 ( \64377 , \64274 , \64376 );
and \U$64035 ( \64378 , \64272 , \64273 );
or \U$64036 ( \64379 , \64377 , \64378 );
and \U$64037 ( \64380 , \64271 , \64379 );
and \U$64038 ( \64381 , \64269 , \64270 );
or \U$64039 ( \64382 , \64380 , \64381 );
and \U$64040 ( \64383 , \64268 , \64382 );
and \U$64041 ( \64384 , \64266 , \64267 );
or \U$64042 ( \64385 , \64383 , \64384 );
and \U$64043 ( \64386 , \64265 , \64385 );
and \U$64044 ( \64387 , \64263 , \64264 );
or \U$64045 ( \64388 , \64386 , \64387 );
and \U$64046 ( \64389 , \64262 , \64388 );
and \U$64047 ( \64390 , \64260 , \64261 );
or \U$64048 ( \64391 , \64389 , \64390 );
and \U$64049 ( \64392 , \64259 , \64391 );
and \U$64050 ( \64393 , \64257 , \64258 );
or \U$64051 ( \64394 , \64392 , \64393 );
and \U$64052 ( \64395 , \64256 , \64394 );
and \U$64053 ( \64396 , \64254 , \64255 );
or \U$64054 ( \64397 , \64395 , \64396 );
and \U$64055 ( \64398 , \64253 , \64397 );
and \U$64056 ( \64399 , \64251 , \64252 );
or \U$64057 ( \64400 , \64398 , \64399 );
and \U$64058 ( \64401 , \64250 , \64400 );
and \U$64059 ( \64402 , \64248 , \64249 );
or \U$64060 ( \64403 , \64401 , \64402 );
and \U$64061 ( \64404 , \64247 , \64403 );
and \U$64062 ( \64405 , \64245 , \64246 );
or \U$64063 ( \64406 , \64404 , \64405 );
and \U$64064 ( \64407 , \64244 , \64406 );
and \U$64065 ( \64408 , \64242 , \64243 );
or \U$64066 ( \64409 , \64407 , \64408 );
and \U$64067 ( \64410 , \64241 , \64409 );
and \U$64068 ( \64411 , \64239 , \64240 );
or \U$64069 ( \64412 , \64410 , \64411 );
and \U$64070 ( \64413 , \64238 , \64412 );
and \U$64071 ( \64414 , \64236 , \64237 );
or \U$64072 ( \64415 , \64413 , \64414 );
and \U$64073 ( \64416 , \64235 , \64415 );
and \U$64074 ( \64417 , \64233 , \64234 );
or \U$64075 ( \64418 , \64416 , \64417 );
and \U$64076 ( \64419 , \64232 , \64418 );
and \U$64077 ( \64420 , \64230 , \64231 );
or \U$64078 ( \64421 , \64419 , \64420 );
and \U$64079 ( \64422 , \64229 , \64421 );
and \U$64080 ( \64423 , \64227 , \64228 );
or \U$64081 ( \64424 , \64422 , \64423 );
and \U$64082 ( \64425 , \64226 , \64424 );
and \U$64083 ( \64426 , \64224 , \64225 );
or \U$64084 ( \64427 , \64425 , \64426 );
and \U$64085 ( \64428 , \64223 , \64427 );
and \U$64086 ( \64429 , \64221 , \64222 );
or \U$64087 ( \64430 , \64428 , \64429 );
and \U$64088 ( \64431 , \64220 , \64430 );
and \U$64089 ( \64432 , \64218 , \64219 );
or \U$64090 ( \64433 , \64431 , \64432 );
and \U$64091 ( \64434 , \64217 , \64433 );
and \U$64092 ( \64435 , \64215 , \64216 );
or \U$64093 ( \64436 , \64434 , \64435 );
and \U$64094 ( \64437 , \64214 , \64436 );
and \U$64095 ( \64438 , \64212 , \64213 );
or \U$64096 ( \64439 , \64437 , \64438 );
and \U$64097 ( \64440 , \64211 , \64439 );
and \U$64098 ( \64441 , \64209 , \64210 );
or \U$64099 ( \64442 , \64440 , \64441 );
and \U$64100 ( \64443 , \64208 , \64442 );
and \U$64101 ( \64444 , \64206 , \64207 );
or \U$64102 ( \64445 , \64443 , \64444 );
and \U$64103 ( \64446 , \64205 , \64445 );
and \U$64104 ( \64447 , \64203 , \64204 );
or \U$64105 ( \64448 , \64446 , \64447 );
and \U$64106 ( \64449 , \64202 , \64448 );
and \U$64107 ( \64450 , \64200 , \64201 );
or \U$64108 ( \64451 , \64449 , \64450 );
and \U$64109 ( \64452 , \64199 , \64451 );
and \U$64110 ( \64453 , \64197 , \64198 );
or \U$64111 ( \64454 , \64452 , \64453 );
and \U$64112 ( \64455 , \64196 , \64454 );
and \U$64113 ( \64456 , \64194 , \64195 );
or \U$64114 ( \64457 , \64455 , \64456 );
and \U$64115 ( \64458 , \64193 , \64457 );
and \U$64116 ( \64459 , \64191 , \64192 );
or \U$64117 ( \64460 , \64458 , \64459 );
and \U$64118 ( \64461 , \64190 , \64460 );
and \U$64119 ( \64462 , \64188 , \64189 );
or \U$64120 ( \64463 , \64461 , \64462 );
and \U$64121 ( \64464 , \64187 , \64463 );
and \U$64122 ( \64465 , \64185 , \64186 );
or \U$64123 ( \64466 , \64464 , \64465 );
and \U$64124 ( \64467 , \64184 , \64466 );
and \U$64125 ( \64468 , \64182 , \64183 );
or \U$64126 ( \64469 , \64467 , \64468 );
and \U$64127 ( \64470 , \64181 , \64469 );
and \U$64128 ( \64471 , \64179 , \64180 );
or \U$64129 ( \64472 , \64470 , \64471 );
and \U$64130 ( \64473 , \64178 , \64472 );
and \U$64131 ( \64474 , \64176 , \64177 );
or \U$64132 ( \64475 , \64473 , \64474 );
and \U$64133 ( \64476 , \64175 , \64475 );
and \U$64134 ( \64477 , \64173 , \64174 );
or \U$64135 ( \64478 , \64476 , \64477 );
and \U$64136 ( \64479 , \64172 , \64478 );
and \U$64137 ( \64480 , \64170 , \64171 );
or \U$64138 ( \64481 , \64479 , \64480 );
and \U$64139 ( \64482 , \64169 , \64481 );
and \U$64140 ( \64483 , \64167 , \64168 );
or \U$64141 ( \64484 , \64482 , \64483 );
and \U$64142 ( \64485 , \64166 , \64484 );
and \U$64143 ( \64486 , \64164 , \64165 );
or \U$64144 ( \64487 , \64485 , \64486 );
and \U$64145 ( \64488 , \64163 , \64487 );
and \U$64146 ( \64489 , \64161 , \64162 );
or \U$64147 ( \64490 , \64488 , \64489 );
and \U$64148 ( \64491 , \64160 , \64490 );
and \U$64149 ( \64492 , \64158 , \64159 );
or \U$64150 ( \64493 , \64491 , \64492 );
and \U$64151 ( \64494 , \64157 , \64493 );
and \U$64152 ( \64495 , \64155 , \64156 );
or \U$64153 ( \64496 , \64494 , \64495 );
and \U$64154 ( \64497 , \64154 , \64496 );
and \U$64155 ( \64498 , \64152 , \64153 );
or \U$64156 ( \64499 , \64497 , \64498 );
and \U$64157 ( \64500 , \64151 , \64499 );
and \U$64158 ( \64501 , \64149 , \64150 );
or \U$64159 ( \64502 , \64500 , \64501 );
and \U$64160 ( \64503 , \64148 , \64502 );
and \U$64161 ( \64504 , \64146 , \64147 );
or \U$64162 ( \64505 , \64503 , \64504 );
and \U$64163 ( \64506 , \64145 , \64505 );
and \U$64164 ( \64507 , \64143 , \64144 );
or \U$64165 ( \64508 , \64506 , \64507 );
and \U$64166 ( \64509 , \64142 , \64508 );
and \U$64167 ( \64510 , \64140 , \64141 );
or \U$64168 ( \64511 , \64509 , \64510 );
or \U$64169 ( \64512 , \64137 , \64138 );
and \U$64170 ( \64513 , \64511 , \64512 );
nor \U$64171 ( \64514 , \64139 , \64513 );
xor \U$64172 ( \64515 , \51837 , \51850 );
xor \U$64173 ( \64516 , \64515 , \63468 );
or \U$64174 ( \64517 , \64514 , \64516 );
not \U$64175 ( \64518 , \64516 );
not \U$64176 ( \64519 , \64514 );
or \U$64177 ( \64520 , \64518 , \64519 );
xor \U$64178 ( \64521 , \32024 , \32016 );
nand \U$64179 ( \64522 , \64520 , \64521 );
nand \U$64180 ( \64523 , \64517 , \64522 );
and \U$64181 ( \64524 , \64136 , \64523 );
and \U$64182 ( \64525 , \64134 , \64135 );
or \U$64183 ( \64526 , \64524 , \64525 );
and \U$64184 ( \64527 , \64133 , \64526 );
and \U$64185 ( \64528 , \64131 , \64132 );
or \U$64186 ( \64529 , \64527 , \64528 );
and \U$64187 ( \64530 , \64127 , \64529 );
and \U$64188 ( \64531 , \64125 , \64126 );
or \U$64189 ( \64532 , \64530 , \64531 );
and \U$64190 ( \64533 , \64124 , \64532 );
and \U$64191 ( \64534 , \64122 , \64123 );
or \U$64192 ( \64535 , \64533 , \64534 );
xor \U$64193 ( \64536 , \49735 , \63496 );
xor \U$64194 ( \64537 , \32121 , \32107 );
or \U$64195 ( \64538 , \64536 , \64537 );
and \U$64196 ( \64539 , \64535 , \64538 );
and \U$64197 ( \64540 , \64537 , \64536 );
nor \U$64198 ( \64541 , \64539 , \64540 );
xnor \U$64199 ( \64542 , \18057 , \32124 );
or \U$64200 ( \64543 , \64541 , \64542 );
not \U$64201 ( \64544 , \64542 );
not \U$64202 ( \64545 , \64541 );
or \U$64203 ( \64546 , \64544 , \64545 );
xor \U$64204 ( \64547 , \49281 , \63498 );
nand \U$64205 ( \64548 , \64546 , \64547 );
nand \U$64206 ( \64549 , \64543 , \64548 );
and \U$64207 ( \64550 , \64121 , \64549 );
nor \U$64208 ( \64551 , \64120 , \64550 );
xor \U$64209 ( \64552 , \47849 , \48365 );
xor \U$64210 ( \64553 , \64552 , \63519 );
or \U$64211 ( \64554 , \64551 , \64553 );
not \U$64212 ( \64555 , \64553 );
not \U$64213 ( \64556 , \64551 );
or \U$64214 ( \64557 , \64555 , \64556 );
xor \U$64215 ( \64558 , \32160 , \32151 );
nand \U$64216 ( \64559 , \64557 , \64558 );
nand \U$64217 ( \64560 , \64554 , \64559 );
and \U$64218 ( \64561 , \64113 , \64560 );
and \U$64219 ( \64562 , \64111 , \64112 );
or \U$64220 ( \64563 , \64561 , \64562 );
and \U$64221 ( \64564 , \64110 , \64563 );
and \U$64222 ( \64565 , \64108 , \64109 );
or \U$64223 ( \64566 , \64564 , \64565 );
and \U$64224 ( \64567 , \64103 , \64566 );
and \U$64225 ( \64568 , \64101 , \64102 );
or \U$64226 ( \64569 , \64567 , \64568 );
and \U$64227 ( \64570 , \64100 , \64569 );
and \U$64228 ( \64571 , \64098 , \64099 );
or \U$64229 ( \64572 , \64570 , \64571 );
xor \U$64230 ( \64573 , \46055 , \63641 );
xor \U$64231 ( \64574 , \14676 , \32183 );
or \U$64232 ( \64575 , \64573 , \64574 );
and \U$64233 ( \64576 , \64572 , \64575 );
and \U$64234 ( \64577 , \64574 , \64573 );
nor \U$64235 ( \64578 , \64576 , \64577 );
xnor \U$64236 ( \64579 , \45629 , \63643 );
or \U$64237 ( \64580 , \64578 , \64579 );
not \U$64238 ( \64581 , \64579 );
not \U$64239 ( \64582 , \64578 );
or \U$64240 ( \64583 , \64581 , \64582 );
xor \U$64241 ( \64584 , \32189 , \32185 );
nand \U$64242 ( \64585 , \64583 , \64584 );
nand \U$64243 ( \64586 , \64580 , \64585 );
xor \U$64244 ( \64587 , \32193 , \32192 );
or \U$64245 ( \64588 , \64586 , \64587 );
xor \U$64246 ( \64589 , \63646 , \63645 );
and \U$64247 ( \64590 , \64588 , \64589 );
and \U$64248 ( \64591 , \64587 , \64586 );
nor \U$64249 ( \64592 , \64590 , \64591 );
xnor \U$64250 ( \64593 , \32198 , \32195 );
or \U$64251 ( \64594 , \64592 , \64593 );
not \U$64252 ( \64595 , \64593 );
not \U$64253 ( \64596 , \64592 );
or \U$64254 ( \64597 , \64595 , \64596 );
xor \U$64255 ( \64598 , \63651 , \63648 );
nand \U$64256 ( \64599 , \64597 , \64598 );
nand \U$64257 ( \64600 , \64594 , \64599 );
and \U$64258 ( \64601 , \64097 , \64600 );
and \U$64259 ( \64602 , \64095 , \64096 );
or \U$64260 ( \64603 , \64601 , \64602 );
and \U$64261 ( \64604 , \64094 , \64603 );
and \U$64262 ( \64605 , \64092 , \64093 );
or \U$64263 ( \64606 , \64604 , \64605 );
and \U$64264 ( \64607 , \64091 , \64606 );
and \U$64265 ( \64608 , \64089 , \64090 );
or \U$64266 ( \64609 , \64607 , \64608 );
xor \U$64267 ( \64610 , \32216 , \32213 );
or \U$64268 ( \64611 , \64609 , \64610 );
xor \U$64269 ( \64612 , \63665 , \63662 );
and \U$64270 ( \64613 , \64611 , \64612 );
and \U$64271 ( \64614 , \64610 , \64609 );
nor \U$64272 ( \64615 , \64613 , \64614 );
xnor \U$64273 ( \64616 , \63669 , \63668 );
or \U$64274 ( \64617 , \64615 , \64616 );
not \U$64275 ( \64618 , \64616 );
not \U$64276 ( \64619 , \64615 );
or \U$64277 ( \64620 , \64618 , \64619 );
xor \U$64278 ( \64621 , \32220 , \32219 );
nand \U$64279 ( \64622 , \64620 , \64621 );
nand \U$64280 ( \64623 , \64617 , \64622 );
and \U$64281 ( \64624 , \64088 , \64623 );
and \U$64282 ( \64625 , \64086 , \64087 );
or \U$64283 ( \64626 , \64624 , \64625 );
xor \U$64284 ( \64627 , \42097 , \63681 );
xor \U$64285 ( \64628 , \32298 , \32264 );
or \U$64286 ( \64629 , \64627 , \64628 );
and \U$64287 ( \64630 , \64626 , \64629 );
and \U$64288 ( \64631 , \64628 , \64627 );
nor \U$64289 ( \64632 , \64630 , \64631 );
xnor \U$64290 ( \64633 , \41718 , \63683 );
or \U$64291 ( \64634 , \64632 , \64633 );
not \U$64292 ( \64635 , \64633 );
not \U$64293 ( \64636 , \64632 );
or \U$64294 ( \64637 , \64635 , \64636 );
xor \U$64295 ( \64638 , \32325 , \32301 );
nand \U$64296 ( \64639 , \64637 , \64638 );
nand \U$64297 ( \64640 , \64634 , \64639 );
and \U$64298 ( \64641 , \64085 , \64640 );
and \U$64299 ( \64642 , \64083 , \64084 );
or \U$64300 ( \64643 , \64641 , \64642 );
and \U$64301 ( \64644 , \64082 , \64643 );
and \U$64302 ( \64645 , \64080 , \64081 );
or \U$64303 ( \64646 , \64644 , \64645 );
xor \U$64304 ( \64647 , \63712 , \63711 );
or \U$64305 ( \64648 , \64646 , \64647 );
xor \U$64306 ( \64649 , \32342 , \32341 );
and \U$64307 ( \64650 , \64648 , \64649 );
and \U$64308 ( \64651 , \64647 , \64646 );
nor \U$64309 ( \64652 , \64650 , \64651 );
xnor \U$64310 ( \64653 , \40203 , \63714 );
or \U$64311 ( \64654 , \64652 , \64653 );
not \U$64312 ( \64655 , \64653 );
not \U$64313 ( \64656 , \64652 );
or \U$64314 ( \64657 , \64655 , \64656 );
xor \U$64315 ( \64658 , \32351 , \32344 );
nand \U$64316 ( \64659 , \64657 , \64658 );
nand \U$64317 ( \64660 , \64654 , \64659 );
and \U$64318 ( \64661 , \64079 , \64660 );
and \U$64319 ( \64662 , \64077 , \64078 );
or \U$64320 ( \64663 , \64661 , \64662 );
and \U$64321 ( \64664 , \64076 , \64663 );
and \U$64322 ( \64665 , \64074 , \64075 );
or \U$64323 ( \64666 , \64664 , \64665 );
and \U$64324 ( \64667 , \64073 , \64666 );
and \U$64325 ( \64668 , \64071 , \64072 );
or \U$64326 ( \64669 , \64667 , \64668 );
not \U$64327 ( \64670 , \38640 );
not \U$64328 ( \64671 , \63732 );
or \U$64329 ( \64672 , \64670 , \64671 );
or \U$64330 ( \64673 , \63732 , \38640 );
nand \U$64331 ( \64674 , \64672 , \64673 );
xor \U$64332 ( \64675 , \32387 , \32371 );
or \U$64333 ( \64676 , \64674 , \64675 );
and \U$64334 ( \64677 , \64669 , \64676 );
and \U$64335 ( \64678 , \64675 , \64674 );
nor \U$64336 ( \64679 , \64677 , \64678 );
xnor \U$64337 ( \64680 , \38344 , \63735 );
or \U$64338 ( \64681 , \64679 , \64680 );
not \U$64339 ( \64682 , \64680 );
not \U$64340 ( \64683 , \64679 );
or \U$64341 ( \64684 , \64682 , \64683 );
xor \U$64342 ( \64685 , \32398 , \32390 );
nand \U$64343 ( \64686 , \64684 , \64685 );
nand \U$64344 ( \64687 , \64681 , \64686 );
nand \U$64345 ( \64688 , \64067 , \64687 );
nand \U$64346 ( \64689 , \64064 , \64688 );
and \U$64347 ( \64690 , \64061 , \64689 );
nor \U$64348 ( \64691 , \64060 , \64690 );
xnor \U$64349 ( \64692 , \32414 , \32406 );
or \U$64350 ( \64693 , \64691 , \64692 );
not \U$64351 ( \64694 , \64692 );
not \U$64352 ( \64695 , \64691 );
or \U$64353 ( \64696 , \64694 , \64695 );
xor \U$64354 ( \64697 , \63820 , \63803 );
nand \U$64355 ( \64698 , \64696 , \64697 );
nand \U$64356 ( \64699 , \64693 , \64698 );
and \U$64357 ( \64700 , \64057 , \64699 );
and \U$64358 ( \64701 , \64055 , \64056 );
or \U$64359 ( \64702 , \64700 , \64701 );
and \U$64360 ( \64703 , \64054 , \64702 );
nor \U$64361 ( \64704 , \64053 , \64703 );
xor \U$64362 ( \64705 , \36509 , \36798 );
xor \U$64363 ( \64706 , \64705 , \63836 );
or \U$64364 ( \64707 , \64704 , \64706 );
not \U$64365 ( \64708 , \64706 );
not \U$64366 ( \64709 , \64704 );
or \U$64367 ( \64710 , \64708 , \64709 );
xor \U$64368 ( \64711 , \32442 , \32421 );
nand \U$64369 ( \64712 , \64710 , \64711 );
nand \U$64370 ( \64713 , \64707 , \64712 );
nand \U$64371 ( \64714 , \64050 , \64713 );
nand \U$64372 ( \64715 , \64047 , \64714 );
not \U$64373 ( \64716 , \63863 );
not \U$64374 ( \64717 , \63841 );
or \U$64375 ( \64718 , \64716 , \64717 );
or \U$64376 ( \64719 , \63841 , \63863 );
nand \U$64377 ( \64720 , \64718 , \64719 );
and \U$64378 ( \64721 , \4437 , \32453 );
not \U$64379 ( \64722 , \4437 );
and \U$64380 ( \64723 , \64722 , \32452 );
nor \U$64381 ( \64724 , \64721 , \64723 );
or \U$64382 ( \64725 , \64720 , \64724 );
and \U$64383 ( \64726 , \64715 , \64725 );
and \U$64384 ( \64727 , \64724 , \64720 );
nor \U$64385 ( \64728 , \64726 , \64727 );
xor \U$64386 ( \64729 , \4139 , \4144 );
xor \U$64387 ( \64730 , \64729 , \32455 );
or \U$64388 ( \64731 , \64728 , \64730 );
not \U$64389 ( \64732 , \64730 );
not \U$64390 ( \64733 , \64728 );
or \U$64391 ( \64734 , \64732 , \64733 );
xor \U$64392 ( \64735 , \63874 , \63866 );
nand \U$64393 ( \64736 , \64734 , \64735 );
nand \U$64394 ( \64737 , \64731 , \64736 );
nand \U$64395 ( \64738 , \64044 , \64737 );
nand \U$64396 ( \64739 , \64041 , \64738 );
xor \U$64397 ( \64740 , \32477 , \32460 );
and \U$64398 ( \64741 , \64739 , \64740 );
not \U$64399 ( \64742 , \64739 );
not \U$64400 ( \64743 , \64740 );
and \U$64401 ( \64744 , \64742 , \64743 );
and \U$64402 ( \64745 , \63879 , \63880 );
nor \U$64403 ( \64746 , \64744 , \64745 );
and \U$64404 ( \64747 , \63881 , \64746 );
nor \U$64405 ( \64748 , \64038 , \64741 , \64747 );
or \U$64406 ( \64749 , \64037 , \64748 );
or \U$64407 ( \64750 , \64023 , \64022 );
nand \U$64408 ( \64751 , \64030 , \64749 , \64750 );
and \U$64409 ( \64752 , \64025 , \64751 );
and \U$64410 ( \64753 , \64017 , \64019 );
nor \U$64411 ( \64754 , \64752 , \64753 );
nor \U$64412 ( \64755 , \64016 , \64754 );
nor \U$64413 ( \64756 , \64013 , \64755 );
xor \U$64414 ( \64757 , \34020 , \34035 );
xor \U$64415 ( \64758 , \64757 , \63916 );
or \U$64416 ( \64759 , \64756 , \64758 );
not \U$64417 ( \64760 , \64758 );
not \U$64418 ( \64761 , \64756 );
or \U$64419 ( \64762 , \64760 , \64761 );
xor \U$64420 ( \64763 , \32590 , \32582 );
nand \U$64421 ( \64764 , \64762 , \64763 );
nand \U$64422 ( \64765 , \64759 , \64764 );
and \U$64423 ( \64766 , \64010 , \64765 );
nor \U$64424 ( \64767 , \64009 , \64766 );
xor \U$64425 ( \64768 , \33658 , \33688 );
xor \U$64426 ( \64769 , \64768 , \63930 );
or \U$64427 ( \64770 , \64767 , \64769 );
not \U$64428 ( \64771 , \64769 );
not \U$64429 ( \64772 , \64767 );
or \U$64430 ( \64773 , \64771 , \64772 );
xor \U$64431 ( \64774 , \32646 , \32595 );
nand \U$64432 ( \64775 , \64773 , \64774 );
nand \U$64433 ( \64776 , \64770 , \64775 );
nand \U$64434 ( \64777 , \64006 , \64776 );
nand \U$64435 ( \64778 , \64003 , \64777 );
and \U$64436 ( \64779 , \64000 , \64778 );
and \U$64437 ( \64780 , \63999 , \63998 );
nor \U$64438 ( \64781 , \64779 , \64780 );
xnor \U$64439 ( \64782 , \32713 , \32705 );
or \U$64440 ( \64783 , \64781 , \64782 );
not \U$64441 ( \64784 , \64782 );
not \U$64442 ( \64785 , \64781 );
or \U$64443 ( \64786 , \64784 , \64785 );
xor \U$64444 ( \64787 , \33163 , \63973 );
nand \U$64445 ( \64788 , \64786 , \64787 );
nand \U$64446 ( \64789 , \64783 , \64788 );
and \U$64447 ( \64790 , \63997 , \64789 );
and \U$64448 ( \64791 , \63995 , \63996 );
or \U$64449 ( \64792 , \64790 , \64791 );
not \U$64450 ( \64793 , \64792 );
and \U$64451 ( \64794 , \376 , RI986e260_13);
and \U$64452 ( \64795 , RI986e350_15, \374 );
nor \U$64453 ( \64796 , \64794 , \64795 );
and \U$64454 ( \64797 , \395 , RI986e170_11);
and \U$64455 ( \64798 , RI986e080_9, \393 );
nor \U$64456 ( \64799 , \64797 , \64798 );
xnor \U$64457 ( \64800 , \64796 , \64799 );
not \U$64458 ( \64801 , \64800 );
and \U$64459 ( \64802 , \64793 , \64801 );
and \U$64460 ( \64803 , \64792 , \64800 );
nor \U$64461 ( \64804 , \64802 , \64803 );
not \U$64462 ( \64805 , \64804 );
and \U$64463 ( \64806 , \354 , RI986ddb0_3);
and \U$64464 ( \64807 , RI986dcc0_1, \352 );
nor \U$64465 ( \64808 , \64806 , \64807 );
and \U$64466 ( \64809 , \416 , RI986df90_7);
and \U$64467 ( \64810 , RI986dea0_5, \414 );
nor \U$64468 ( \64811 , \64809 , \64810 );
xnor \U$64469 ( \64812 , \64808 , \64811 );
not \U$64470 ( \64813 , \64812 );
and \U$64471 ( \64814 , \376 , RI986e2d8_14);
and \U$64472 ( \64815 , RI986e3c8_16, \374 );
nor \U$64473 ( \64816 , \64814 , \64815 );
and \U$64474 ( \64817 , \395 , RI986e1e8_12);
and \U$64475 ( \64818 , RI986e0f8_10, \393 );
nor \U$64476 ( \64819 , \64817 , \64818 );
xor \U$64477 ( \64820 , \64816 , \64819 );
not \U$64478 ( \64821 , \64820 );
or \U$64479 ( \64822 , \64813 , \64821 );
or \U$64480 ( \64823 , \64812 , \64820 );
nand \U$64481 ( \64824 , \64822 , \64823 );
not \U$64482 ( \64825 , \64824 );
and \U$64483 ( \64826 , \64805 , \64825 );
and \U$64484 ( \64827 , \64804 , \64824 );
nor \U$64485 ( \64828 , \64826 , \64827 );
not \U$64486 ( \64829 , \64828 );
or \U$64487 ( \64830 , \63994 , \64829 );
or \U$64488 ( \64831 , \64828 , \63993 );
nand \U$64489 ( \64832 , \64830 , \64831 );
not \U$64490 ( \64833 , \64832 );
or \U$64491 ( \64834 , \32821 , \64833 );
or \U$64492 ( \64835 , \64832 , \32820 );
nand \U$64493 ( \64836 , \64834 , \64835 );
xnor \U$64494 ( \64837 , RI9874ae8_236, RI9874f20_245);
not \U$64495 ( \64838 , \64837 );
xor \U$64496 ( \64839 , RI98745c0_225, RI9874a70_235);
not \U$64497 ( \64840 , \64839 );
and \U$64498 ( \64841 , \64838 , \64840 );
and \U$64499 ( \64842 , \64837 , \64839 );
nor \U$64500 ( \64843 , \64841 , \64842 );
not \U$64501 ( \64844 , \64843 );
xor \U$64502 ( \64845 , RI9874548_224, RI98736c0_193);
not \U$64503 ( \64846 , \64845 );
xnor \U$64504 ( \64847 , RI9873e40_209, RI9874c50_239);
not \U$64505 ( \64848 , \64847 );
or \U$64506 ( \64849 , \64846 , \64848 );
or \U$64507 ( \64850 , \64847 , \64845 );
nand \U$64508 ( \64851 , \64849 , \64850 );
not \U$64509 ( \64852 , \64851 );
and \U$64510 ( \64853 , \64844 , \64852 );
and \U$64511 ( \64854 , \64843 , \64851 );
nor \U$64512 ( \64855 , \64853 , \64854 );
not \U$64513 ( \64856 , \64855 );
xor \U$64514 ( \64857 , RI9874188_216, RI9874278_218);
not \U$64515 ( \64858 , \64857 );
xnor \U$64516 ( \64859 , RI9873f30_211, RI9874ea8_244);
not \U$64517 ( \64860 , \64859 );
or \U$64518 ( \64861 , \64858 , \64860 );
or \U$64519 ( \64862 , \64859 , \64857 );
nand \U$64520 ( \64863 , \64861 , \64862 );
not \U$64521 ( \64864 , \64863 );
xnor \U$64522 ( \64865 , RI98743e0_221, RI98744d0_223);
not \U$64523 ( \64866 , \64865 );
xor \U$64524 ( \64867 , RI9875358_254, RI9873b70_203);
not \U$64525 ( \64868 , \64867 );
and \U$64526 ( \64869 , \64866 , \64868 );
and \U$64527 ( \64870 , \64865 , \64867 );
nor \U$64528 ( \64871 , \64869 , \64870 );
not \U$64529 ( \64872 , \64871 );
or \U$64530 ( \64873 , \64864 , \64872 );
or \U$64531 ( \64874 , \64871 , \64863 );
nand \U$64532 ( \64875 , \64873 , \64874 );
not \U$64533 ( \64876 , \64875 );
and \U$64534 ( \64877 , \64856 , \64876 );
and \U$64535 ( \64878 , \64855 , \64875 );
nor \U$64536 ( \64879 , \64877 , \64878 );
not \U$64537 ( \64880 , \64879 );
xor \U$64538 ( \64881 , RI98749f8_234, RI9875178_250);
not \U$64539 ( \64882 , \64881 );
xnor \U$64540 ( \64883 , RI9874458_222, RI9874098_214);
not \U$64541 ( \64884 , \64883 );
or \U$64542 ( \64885 , \64882 , \64884 );
or \U$64543 ( \64886 , \64883 , \64881 );
nand \U$64544 ( \64887 , \64885 , \64886 );
not \U$64545 ( \64888 , \64887 );
xnor \U$64546 ( \64889 , RI9873eb8_210, RI9874818_230);
not \U$64547 ( \64890 , \64889 );
xor \U$64548 ( \64891 , RI9874db8_242, RI9875088_248);
not \U$64549 ( \64892 , \64891 );
and \U$64550 ( \64893 , \64890 , \64892 );
and \U$64551 ( \64894 , \64889 , \64891 );
nor \U$64552 ( \64895 , \64893 , \64894 );
not \U$64553 ( \64896 , \64895 );
or \U$64554 ( \64897 , \64888 , \64896 );
or \U$64555 ( \64898 , \64895 , \64887 );
nand \U$64556 ( \64899 , \64897 , \64898 );
not \U$64557 ( \64900 , \64899 );
xnor \U$64558 ( \64901 , RI9874638_226, RI9874b60_237);
not \U$64559 ( \64902 , \64901 );
xor \U$64560 ( \64903 , RI9873738_194, RI9874cc8_240);
not \U$64561 ( \64904 , \64903 );
and \U$64562 ( \64905 , \64902 , \64904 );
and \U$64563 ( \64906 , \64901 , \64903 );
nor \U$64564 ( \64907 , \64905 , \64906 );
not \U$64565 ( \64908 , \64907 );
xor \U$64566 ( \64909 , RI9873918_198, RI9873cd8_206);
not \U$64567 ( \64910 , \64909 );
xnor \U$64568 ( \64911 , RI9873be8_204, RI9875010_247);
not \U$64569 ( \64912 , \64911 );
or \U$64570 ( \64913 , \64910 , \64912 );
or \U$64571 ( \64914 , \64911 , \64909 );
nand \U$64572 ( \64915 , \64913 , \64914 );
not \U$64573 ( \64916 , \64915 );
and \U$64574 ( \64917 , \64908 , \64916 );
and \U$64575 ( \64918 , \64907 , \64915 );
nor \U$64576 ( \64919 , \64917 , \64918 );
not \U$64577 ( \64920 , \64919 );
or \U$64578 ( \64921 , \64900 , \64920 );
or \U$64579 ( \64922 , \64919 , \64899 );
nand \U$64580 ( \64923 , \64921 , \64922 );
not \U$64581 ( \64924 , \64923 );
or \U$64582 ( \64925 , \64880 , \64924 );
or \U$64583 ( \64926 , \64879 , \64923 );
nand \U$64584 ( \64927 , \64925 , \64926 );
xnor \U$64585 ( \64928 , RI9875100_249, RI9874980_233);
not \U$64586 ( \64929 , \64928 );
xor \U$64587 ( \64930 , RI98747a0_229, RI9874020_213);
not \U$64588 ( \64931 , \64930 );
and \U$64589 ( \64932 , \64929 , \64931 );
and \U$64590 ( \64933 , \64928 , \64930 );
nor \U$64591 ( \64934 , \64932 , \64933 );
not \U$64592 ( \64935 , \64934 );
xor \U$64593 ( \64936 , RI9874110_215, RI98737b0_195);
not \U$64594 ( \64937 , \64936 );
xnor \U$64595 ( \64938 , RI9874f98_246, RI9874bd8_238);
not \U$64596 ( \64939 , \64938 );
or \U$64597 ( \64940 , \64937 , \64939 );
or \U$64598 ( \64941 , \64938 , \64936 );
nand \U$64599 ( \64942 , \64940 , \64941 );
not \U$64600 ( \64943 , \64942 );
and \U$64601 ( \64944 , \64935 , \64943 );
and \U$64602 ( \64945 , \64934 , \64942 );
nor \U$64603 ( \64946 , \64944 , \64945 );
not \U$64604 ( \64947 , \64946 );
xor \U$64605 ( \64948 , RI9874890_231, RI9873fa8_212);
not \U$64606 ( \64949 , \64948 );
xnor \U$64607 ( \64950 , RI9873a08_200, RI9873af8_202);
not \U$64608 ( \64951 , \64950 );
or \U$64609 ( \64952 , \64949 , \64951 );
or \U$64610 ( \64953 , \64950 , \64948 );
nand \U$64611 ( \64954 , \64952 , \64953 );
not \U$64612 ( \64955 , \64954 );
xnor \U$64613 ( \64956 , RI98742f0_219, RI98751f0_251);
not \U$64614 ( \64957 , \64956 );
xor \U$64615 ( \64958 , RI9874200_217, RI98738a0_197);
not \U$64616 ( \64959 , \64958 );
and \U$64617 ( \64960 , \64957 , \64959 );
and \U$64618 ( \64961 , \64956 , \64958 );
nor \U$64619 ( \64962 , \64960 , \64961 );
not \U$64620 ( \64963 , \64962 );
or \U$64621 ( \64964 , \64955 , \64963 );
or \U$64622 ( \64965 , \64962 , \64954 );
nand \U$64623 ( \64966 , \64964 , \64965 );
not \U$64624 ( \64967 , \64966 );
and \U$64625 ( \64968 , \64947 , \64967 );
and \U$64626 ( \64969 , \64946 , \64966 );
nor \U$64627 ( \64970 , \64968 , \64969 );
not \U$64628 ( \64971 , \64970 );
xor \U$64629 ( \64972 , RI9873828_196, RI9875268_252);
not \U$64630 ( \64973 , \64972 );
xnor \U$64631 ( \64974 , RI9874368_220, RI9873a80_201);
not \U$64632 ( \64975 , \64974 );
or \U$64633 ( \64976 , \64973 , \64975 );
or \U$64634 ( \64977 , \64974 , \64972 );
nand \U$64635 ( \64978 , \64976 , \64977 );
not \U$64636 ( \64979 , \64978 );
xnor \U$64637 ( \64980 , RI9874728_228, RI9873d50_207);
not \U$64638 ( \64981 , \64980 );
xor \U$64639 ( \64982 , RI9873990_199, RI9874908_232);
not \U$64640 ( \64983 , \64982 );
and \U$64641 ( \64984 , \64981 , \64983 );
and \U$64642 ( \64985 , \64980 , \64982 );
nor \U$64643 ( \64986 , \64984 , \64985 );
not \U$64644 ( \64987 , \64986 );
or \U$64645 ( \64988 , \64979 , \64987 );
or \U$64646 ( \64989 , \64986 , \64978 );
nand \U$64647 ( \64990 , \64988 , \64989 );
not \U$64648 ( \64991 , \64990 );
xnor \U$64649 ( \64992 , RI9874d40_241, RI98746b0_227);
not \U$64650 ( \64993 , \64992 );
xor \U$64651 ( \64994 , RI9874e30_243, RI9873c60_205);
not \U$64652 ( \64995 , \64994 );
and \U$64653 ( \64996 , \64993 , \64995 );
and \U$64654 ( \64997 , \64992 , \64994 );
nor \U$64655 ( \64998 , \64996 , \64997 );
not \U$64656 ( \64999 , \64998 );
xor \U$64657 ( \65000 , RI98752e0_253, RI9875448_256);
not \U$64658 ( \65001 , \65000 );
xnor \U$64659 ( \65002 , RI98753d0_255, RI9873dc8_208);
not \U$64660 ( \65003 , \65002 );
or \U$64661 ( \65004 , \65001 , \65003 );
or \U$64662 ( \65005 , \65002 , \65000 );
nand \U$64663 ( \65006 , \65004 , \65005 );
not \U$64664 ( \65007 , \65006 );
and \U$64665 ( \65008 , \64999 , \65007 );
and \U$64666 ( \65009 , \64998 , \65006 );
nor \U$64667 ( \65010 , \65008 , \65009 );
not \U$64668 ( \65011 , \65010 );
or \U$64669 ( \65012 , \64991 , \65011 );
or \U$64670 ( \65013 , \65010 , \64990 );
nand \U$64671 ( \65014 , \65012 , \65013 );
not \U$64672 ( \65015 , \65014 );
and \U$64673 ( \65016 , \64971 , \65015 );
and \U$64674 ( \65017 , \64970 , \65014 );
nor \U$64675 ( \65018 , \65016 , \65017 );
xor \U$64676 ( \65019 , \64927 , \65018 );
_DC gff1e ( \65020_nGff1e , \64836 , \65019 );
buf \U$64677 ( \65021 , \65020_nGff1e );
xor \U$64678 ( \65022 , \63995 , \63996 );
xor \U$64679 ( \65023 , \65022 , \64789 );
_DC gfe5e ( \65024_nGfe5e , \65023 , \65019 );
buf \U$64680 ( \65025 , \65024_nGfe5e );
not \U$64681 ( \65026 , \64778 );
xnor \U$64682 ( \65027 , \63999 , \63998 );
not \U$64683 ( \65028 , \65027 );
or \U$64684 ( \65029 , \65026 , \65028 );
or \U$64685 ( \65030 , \65027 , \64778 );
nand \U$64686 ( \65031 , \65029 , \65030 );
_DC gfcc0 ( \65032_nGfcc0 , \65031 , \65019 );
buf \U$64687 ( \65033 , \65032_nGfcc0 );
not \U$64688 ( \65034 , \64765 );
xnor \U$64689 ( \65035 , \64008 , \64007 );
not \U$64690 ( \65036 , \65035 );
or \U$64691 ( \65037 , \65034 , \65036 );
or \U$64692 ( \65038 , \65035 , \64765 );
nand \U$64693 ( \65039 , \65037 , \65038 );
_DC gf9d4 ( \65040_nGf9d4 , \65039 , \65019 );
buf \U$64694 ( \65041 , \65040_nGf9d4 );
not \U$64695 ( \65042 , \64754 );
xor \U$64696 ( \65043 , \64012 , \64011 );
not \U$64697 ( \65044 , \65043 );
or \U$64698 ( \65045 , \65042 , \65044 );
or \U$64699 ( \65046 , \65043 , \64754 );
nand \U$64700 ( \65047 , \65045 , \65046 );
_DC gf7a2 ( \65048_nGf7a2 , \65047 , \65019 );
buf \U$64701 ( \65049 , \65048_nGf7a2 );
xnor \U$64702 ( \65050 , \64724 , \64720 );
not \U$64703 ( \65051 , \65050 );
not \U$64704 ( \65052 , \64715 );
or \U$64705 ( \65053 , \65051 , \65052 );
or \U$64706 ( \65054 , \64715 , \65050 );
nand \U$64707 ( \65055 , \65053 , \65054 );
_DC gec11 ( \65056_nGec11 , \65055 , \65019 );
buf \U$64708 ( \65057 , \65056_nGec11 );
xnor \U$64709 ( \65058 , \64052 , \64051 );
not \U$64710 ( \65059 , \65058 );
not \U$64711 ( \65060 , \64702 );
or \U$64712 ( \65061 , \65059 , \65060 );
or \U$64713 ( \65062 , \64702 , \65058 );
nand \U$64714 ( \65063 , \65061 , \65062 );
_DC ge638 ( \65064_nGe638 , \65063 , \65019 );
buf \U$64715 ( \65065 , \65064_nGe638 );
xor \U$64716 ( \65066 , \64055 , \64056 );
xor \U$64717 ( \65067 , \65066 , \64699 );
_DC ge441 ( \65068_nGe441 , \65067 , \65019 );
buf \U$64718 ( \65069 , \65068_nGe441 );
xnor \U$64719 ( \65070 , \64059 , \64058 );
not \U$64720 ( \65071 , \65070 );
not \U$64721 ( \65072 , \64689 );
or \U$64722 ( \65073 , \65071 , \65072 );
or \U$64723 ( \65074 , \64689 , \65070 );
nand \U$64724 ( \65075 , \65073 , \65074 );
_DC ge060 ( \65076_nGe060 , \65075 , \65019 );
buf \U$64725 ( \65077 , \65076_nGe060 );
xnor \U$64726 ( \65078 , \64675 , \64674 );
not \U$64727 ( \65079 , \65078 );
not \U$64728 ( \65080 , \64669 );
or \U$64729 ( \65081 , \65079 , \65080 );
or \U$64730 ( \65082 , \64669 , \65078 );
nand \U$64731 ( \65083 , \65081 , \65082 );
_DC gd9de ( \65084_nGd9de , \65083 , \65019 );
buf \U$64732 ( \65085 , \65084_nGd9de );
xor \U$64733 ( \65086 , \64071 , \64072 );
xor \U$64734 ( \65087 , \65086 , \64666 );
_DC gd7a2 ( \65088_nGd7a2 , \65087 , \65019 );
buf \U$64735 ( \65089 , \65088_nGd7a2 );
xor \U$64736 ( \65090 , \64074 , \64075 );
xor \U$64737 ( \65091 , \65090 , \64663 );
_DC gd59f ( \65092_nGd59f , \65091 , \65019 );
buf \U$64738 ( \65093 , \65092_nGd59f );
xor \U$64739 ( \65094 , \64077 , \64078 );
xor \U$64740 ( \65095 , \65094 , \64660 );
_DC gd368 ( \65096_nGd368 , \65095 , \65019 );
buf \U$64741 ( \65097 , \65096_nGd368 );
xnor \U$64742 ( \65098 , \64649 , \64647 );
not \U$64743 ( \65099 , \65098 );
not \U$64744 ( \65100 , \64646 );
or \U$64745 ( \65101 , \65099 , \65100 );
or \U$64746 ( \65102 , \64646 , \65098 );
nand \U$64747 ( \65103 , \65101 , \65102 );
_DC gcebb ( \65104_nGcebb , \65103 , \65019 );
buf \U$64748 ( \65105 , \65104_nGcebb );
xor \U$64749 ( \65106 , \64080 , \64081 );
xor \U$64750 ( \65107 , \65106 , \64643 );
_DC gcc44 ( \65108_nGcc44 , \65107 , \65019 );
buf \U$64751 ( \65109 , \65108_nGcc44 );
xor \U$64752 ( \65110 , \64083 , \64084 );
xor \U$64753 ( \65111 , \65110 , \64640 );
_DC gc9e1 ( \65112_nGc9e1 , \65111 , \65019 );
buf \U$64754 ( \65113 , \65112_nGc9e1 );
xnor \U$64755 ( \65114 , \64628 , \64627 );
not \U$64756 ( \65115 , \65114 );
not \U$64757 ( \65116 , \64626 );
or \U$64758 ( \65117 , \65115 , \65116 );
or \U$64759 ( \65118 , \64626 , \65114 );
nand \U$64760 ( \65119 , \65117 , \65118 );
_DC gc4a5 ( \65120_nGc4a5 , \65119 , \65019 );
buf \U$64761 ( \65121 , \65120_nGc4a5 );
xor \U$64762 ( \65122 , \64086 , \64087 );
xor \U$64763 ( \65123 , \65122 , \64623 );
_DC gc1e2 ( \65124_nGc1e2 , \65123 , \65019 );
buf \U$64764 ( \65125 , \65124_nGc1e2 );
xnor \U$64765 ( \65126 , \64610 , \64612 );
not \U$64766 ( \65127 , \65126 );
not \U$64767 ( \65128 , \64609 );
or \U$64768 ( \65129 , \65127 , \65128 );
or \U$64769 ( \65130 , \64609 , \65126 );
nand \U$64770 ( \65131 , \65129 , \65130 );
_DC gbc0f ( \65132_nGbc0f , \65131 , \65019 );
buf \U$64771 ( \65133 , \65132_nGbc0f );
xor \U$64772 ( \65134 , \64089 , \64090 );
xor \U$64773 ( \65135 , \65134 , \64606 );
_DC gb8f8 ( \65136_nGb8f8 , \65135 , \65019 );
buf \U$64774 ( \65137 , \65136_nGb8f8 );
xor \U$64775 ( \65138 , \64092 , \64093 );
xor \U$64776 ( \65139 , \65138 , \64603 );
_DC gb5fc ( \65140_nGb5fc , \65139 , \65019 );
buf \U$64777 ( \65141 , \65140_nGb5fc );
xor \U$64778 ( \65142 , \64095 , \64096 );
xor \U$64779 ( \65143 , \65142 , \64600 );
_DC gb31e ( \65144_nGb31e , \65143 , \65019 );
buf \U$64780 ( \65145 , \65144_nGb31e );
not \U$64781 ( \65146 , \64572 );
xnor \U$64782 ( \65147 , \64574 , \64573 );
not \U$64783 ( \65148 , \65147 );
or \U$64784 ( \65149 , \65146 , \65148 );
or \U$64785 ( \65150 , \65147 , \64572 );
nand \U$64786 ( \65151 , \65149 , \65150 );
_DC ga763 ( \65152_nGa763 , \65151 , \65019 );
buf \U$64787 ( \65153 , \65152_nGa763 );
xor \U$64788 ( \65154 , \64098 , \64099 );
xor \U$64789 ( \65155 , \65154 , \64569 );
_DC ga455 ( \65156_nGa455 , \65155 , \65019 );
buf \U$64790 ( \65157 , \65156_nGa455 );
xor \U$64791 ( \65158 , \64101 , \64102 );
xor \U$64792 ( \65159 , \65158 , \64566 );
_DC ga121 ( \65160_nGa121 , \65159 , \65019 );
buf \U$64793 ( \65161 , \65160_nGa121 );
xor \U$64794 ( \65162 , \64108 , \64109 );
xor \U$64795 ( \65163 , \65162 , \64563 );
_DC g9e06 ( \65164_nG9e06 , \65163 , \65019 );
buf \U$64796 ( \65165 , \65164_nG9e06 );
xor \U$64797 ( \65166 , \64111 , \64112 );
xor \U$64798 ( \65167 , \65166 , \64560 );
_DC g9ab5 ( \65168_nG9ab5 , \65167 , \65019 );
buf \U$64799 ( \65169 , \65168_nG9ab5 );
not \U$64800 ( \65170 , \64549 );
xnor \U$64801 ( \65171 , \64119 , \64118 );
not \U$64802 ( \65172 , \65171 );
or \U$64803 ( \65173 , \65170 , \65172 );
or \U$64804 ( \65174 , \65171 , \64549 );
nand \U$64805 ( \65175 , \65173 , \65174 );
_DC g93cf ( \65176_nG93cf , \65175 , \65019 );
buf \U$64806 ( \65177 , \65176_nG93cf );
not \U$64807 ( \65178 , \64535 );
xnor \U$64808 ( \65179 , \64537 , \64536 );
not \U$64809 ( \65180 , \65179 );
or \U$64810 ( \65181 , \65178 , \65180 );
or \U$64811 ( \65182 , \65179 , \64535 );
nand \U$64812 ( \65183 , \65181 , \65182 );
_DC g8c6c ( \65184_nG8c6c , \65183 , \65019 );
buf \U$64813 ( \65185 , \65184_nG8c6c );
xor \U$64814 ( \65186 , \64122 , \64123 );
xor \U$64815 ( \65187 , \65186 , \64532 );
_DC g88da ( \65188_nG88da , \65187 , \65019 );
buf \U$64816 ( \65189 , \65188_nG88da );
xor \U$64817 ( \65190 , \64125 , \64126 );
xor \U$64818 ( \65191 , \65190 , \64529 );
_DC g84f5 ( \65192_nG84f5 , \65191 , \65019 );
buf \U$64819 ( \65193 , \65192_nG84f5 );
xor \U$64820 ( \65194 , \64131 , \64132 );
xor \U$64821 ( \65195 , \65194 , \64526 );
_DC g80db ( \65196_nG80db , \65195 , \65019 );
buf \U$64822 ( \65197 , \65196_nG80db );
xor \U$64823 ( \65198 , \64134 , \64135 );
xor \U$64824 ( \65199 , \65198 , \64523 );
_DC g7cdd ( \65200_nG7cdd , \65199 , \65019 );
buf \U$64825 ( \65201 , \65200_nG7cdd );
not \U$64826 ( \65202 , \64511 );
xnor \U$64827 ( \65203 , \64138 , \64137 );
not \U$64828 ( \65204 , \65203 );
or \U$64829 ( \65205 , \65202 , \65204 );
or \U$64830 ( \65206 , \65203 , \64511 );
nand \U$64831 ( \65207 , \65205 , \65206 );
_DC g7550 ( \65208_nG7550 , \65207 , \65019 );
buf \U$64832 ( \65209 , \65208_nG7550 );
xor \U$64833 ( \65210 , \64140 , \64141 );
xor \U$64834 ( \65211 , \65210 , \64508 );
_DC g71d5 ( \65212_nG71d5 , \65211 , \65019 );
buf \U$64835 ( \65213 , \65212_nG71d5 );
xor \U$64836 ( \65214 , \64143 , \64144 );
xor \U$64837 ( \65215 , \65214 , \64505 );
_DC g6e56 ( \65216_nG6e56 , \65215 , \65019 );
buf \U$64838 ( \65217 , \65216_nG6e56 );
xor \U$64839 ( \65218 , \64146 , \64147 );
xor \U$64840 ( \65219 , \65218 , \64502 );
_DC g6aad ( \65220_nG6aad , \65219 , \65019 );
buf \U$64841 ( \65221 , \65220_nG6aad );
xor \U$64842 ( \65222 , \64149 , \64150 );
xor \U$64843 ( \65223 , \65222 , \64499 );
_DC g6724 ( \65224_nG6724 , \65223 , \65019 );
buf \U$64844 ( \65225 , \65224_nG6724 );
xor \U$64845 ( \65226 , \64152 , \64153 );
xor \U$64846 ( \65227 , \65226 , \64496 );
_DC g63c0 ( \65228_nG63c0 , \65227 , \65019 );
buf \U$64847 ( \65229 , \65228_nG63c0 );
xor \U$64848 ( \65230 , \64155 , \64156 );
xor \U$64849 ( \65231 , \65230 , \64493 );
_DC g6058 ( \65232_nG6058 , \65231 , \65019 );
buf \U$64850 ( \65233 , \65232_nG6058 );
xor \U$64851 ( \65234 , \64158 , \64159 );
xor \U$64852 ( \65235 , \65234 , \64490 );
_DC g5ce5 ( \65236_nG5ce5 , \65235 , \65019 );
buf \U$64853 ( \65237 , \65236_nG5ce5 );
xor \U$64854 ( \65238 , \64161 , \64162 );
xor \U$64855 ( \65239 , \65238 , \64487 );
_DC g59a6 ( \65240_nG59a6 , \65239 , \65019 );
buf \U$64856 ( \65241 , \65240_nG59a6 );
xor \U$64857 ( \65242 , \64164 , \64165 );
xor \U$64858 ( \65243 , \65242 , \64484 );
_DC g5674 ( \65244_nG5674 , \65243 , \65019 );
buf \U$64859 ( \65245 , \65244_nG5674 );
xor \U$64860 ( \65246 , \64167 , \64168 );
xor \U$64861 ( \65247 , \65246 , \64481 );
_DC g5358 ( \65248_nG5358 , \65247 , \65019 );
buf \U$64862 ( \65249 , \65248_nG5358 );
xor \U$64863 ( \65250 , \64170 , \64171 );
xor \U$64864 ( \65251 , \65250 , \64478 );
_DC g5053 ( \65252_nG5053 , \65251 , \65019 );
buf \U$64865 ( \65253 , \65252_nG5053 );
xor \U$64866 ( \65254 , \64173 , \64174 );
xor \U$64867 ( \65255 , \65254 , \64475 );
_DC g4d41 ( \65256_nG4d41 , \65255 , \65019 );
buf \U$64868 ( \65257 , \65256_nG4d41 );
xor \U$64869 ( \65258 , \64176 , \64177 );
xor \U$64870 ( \65259 , \65258 , \64472 );
_DC g4a68 ( \65260_nG4a68 , \65259 , \65019 );
buf \U$64871 ( \65261 , \65260_nG4a68 );
xor \U$64872 ( \65262 , \64179 , \64180 );
xor \U$64873 ( \65263 , \65262 , \64469 );
_DC g4793 ( \65264_nG4793 , \65263 , \65019 );
buf \U$64874 ( \65265 , \65264_nG4793 );
xor \U$64875 ( \65266 , \64182 , \64183 );
xor \U$64876 ( \65267 , \65266 , \64466 );
_DC g44bd ( \65268_nG44bd , \65267 , \65019 );
buf \U$64877 ( \65269 , \65268_nG44bd );
xor \U$64878 ( \65270 , \64185 , \64186 );
xor \U$64879 ( \65271 , \65270 , \64463 );
_DC g41fa ( \65272_nG41fa , \65271 , \65019 );
buf \U$64880 ( \65273 , \65272_nG41fa );
xor \U$64881 ( \65274 , \64188 , \64189 );
xor \U$64882 ( \65275 , \65274 , \64460 );
_DC g3f43 ( \65276_nG3f43 , \65275 , \65019 );
buf \U$64883 ( \65277 , \65276_nG3f43 );
xor \U$64884 ( \65278 , \64191 , \64192 );
xor \U$64885 ( \65279 , \65278 , \64457 );
_DC g3cb4 ( \65280_nG3cb4 , \65279 , \65019 );
buf \U$64886 ( \65281 , \65280_nG3cb4 );
xor \U$64887 ( \65282 , \64194 , \64195 );
xor \U$64888 ( \65283 , \65282 , \64454 );
_DC g3a4a ( \65284_nG3a4a , \65283 , \65019 );
buf \U$64889 ( \65285 , \65284_nG3a4a );
xor \U$64890 ( \65286 , \64197 , \64198 );
xor \U$64891 ( \65287 , \65286 , \64451 );
_DC g37e1 ( \65288_nG37e1 , \65287 , \65019 );
buf \U$64892 ( \65289 , \65288_nG37e1 );
xor \U$64893 ( \65290 , \64200 , \64201 );
xor \U$64894 ( \65291 , \65290 , \64448 );
_DC g358f ( \65292_nG358f , \65291 , \65019 );
buf \U$64895 ( \65293 , \65292_nG358f );
xor \U$64896 ( \65294 , \64203 , \64204 );
xor \U$64897 ( \65295 , \65294 , \64445 );
_DC g332f ( \65296_nG332f , \65295 , \65019 );
buf \U$64898 ( \65297 , \65296_nG332f );
xor \U$64899 ( \65298 , \64206 , \64207 );
xor \U$64900 ( \65299 , \65298 , \64442 );
_DC g30bf ( \65300_nG30bf , \65299 , \65019 );
buf \U$64901 ( \65301 , \65300_nG30bf );
xor \U$64902 ( \65302 , \64209 , \64210 );
xor \U$64903 ( \65303 , \65302 , \64439 );
_DC g2e68 ( \65304_nG2e68 , \65303 , \65019 );
buf \U$64904 ( \65305 , \65304_nG2e68 );
xor \U$64905 ( \65306 , \64212 , \64213 );
xor \U$64906 ( \65307 , \65306 , \64436 );
_DC g2bfd ( \65308_nG2bfd , \65307 , \65019 );
buf \U$64907 ( \65309 , \65308_nG2bfd );
xor \U$64908 ( \65310 , \64215 , \64216 );
xor \U$64909 ( \65311 , \65310 , \64433 );
_DC g29b2 ( \65312_nG29b2 , \65311 , \65019 );
buf \U$64910 ( \65313 , \65312_nG29b2 );
xor \U$64911 ( \65314 , \64218 , \64219 );
xor \U$64912 ( \65315 , \65314 , \64430 );
_DC g276d ( \65316_nG276d , \65315 , \65019 );
buf \U$64913 ( \65317 , \65316_nG276d );
xor \U$64914 ( \65318 , \64221 , \64222 );
xor \U$64915 ( \65319 , \65318 , \64427 );
_DC g2549 ( \65320_nG2549 , \65319 , \65019 );
buf \U$64916 ( \65321 , \65320_nG2549 );
xor \U$64917 ( \65322 , \64224 , \64225 );
xor \U$64918 ( \65323 , \65322 , \64424 );
_DC g2359 ( \65324_nG2359 , \65323 , \65019 );
buf \U$64919 ( \65325 , \65324_nG2359 );
xor \U$64920 ( \65326 , \64227 , \64228 );
xor \U$64921 ( \65327 , \65326 , \64421 );
_DC g2175 ( \65328_nG2175 , \65327 , \65019 );
buf \U$64922 ( \65329 , \65328_nG2175 );
xor \U$64923 ( \65330 , \64230 , \64231 );
xor \U$64924 ( \65331 , \65330 , \64418 );
_DC g1f9c ( \65332_nG1f9c , \65331 , \65019 );
buf \U$64925 ( \65333 , \65332_nG1f9c );
xor \U$64926 ( \65334 , \64233 , \64234 );
xor \U$64927 ( \65335 , \65334 , \64415 );
_DC g1dda ( \65336_nG1dda , \65335 , \65019 );
buf \U$64928 ( \65337 , \65336_nG1dda );
xor \U$64929 ( \65338 , \64236 , \64237 );
xor \U$64930 ( \65339 , \65338 , \64412 );
_DC g1c2e ( \65340_nG1c2e , \65339 , \65019 );
buf \U$64931 ( \65341 , \65340_nG1c2e );
xor \U$64932 ( \65342 , \64239 , \64240 );
xor \U$64933 ( \65343 , \65342 , \64409 );
_DC g1a7f ( \65344_nG1a7f , \65343 , \65019 );
buf \U$64934 ( \65345 , \65344_nG1a7f );
xor \U$64935 ( \65346 , \64242 , \64243 );
xor \U$64936 ( \65347 , \65346 , \64406 );
_DC g18e2 ( \65348_nG18e2 , \65347 , \65019 );
buf \U$64937 ( \65349 , \65348_nG18e2 );
xor \U$64938 ( \65350 , \64245 , \64246 );
xor \U$64939 ( \65351 , \65350 , \64403 );
_DC g173e ( \65352_nG173e , \65351 , \65019 );
buf \U$64940 ( \65353 , \65352_nG173e );
xor \U$64941 ( \65354 , \64248 , \64249 );
xor \U$64942 ( \65355 , \65354 , \64400 );
_DC gff30 ( \65356_nGff30 , \65355 , \65019 );
buf \U$64943 ( \65357 , \65356_nGff30 );
xor \U$64944 ( \65358 , \64251 , \64252 );
xor \U$64945 ( \65359 , \65358 , \64397 );
_DC gff2d ( \65360_nGff2d , \65359 , \65019 );
buf \U$64946 ( \65361 , \65360_nGff2d );
xor \U$64947 ( \65362 , \64254 , \64255 );
xor \U$64948 ( \65363 , \65362 , \64394 );
_DC gff2a ( \65364_nGff2a , \65363 , \65019 );
buf \U$64949 ( \65365 , \65364_nGff2a );
xor \U$64950 ( \65366 , \64257 , \64258 );
xor \U$64951 ( \65367 , \65366 , \64391 );
_DC gff27 ( \65368_nGff27 , \65367 , \65019 );
buf \U$64952 ( \65369 , \65368_nGff27 );
xor \U$64953 ( \65370 , \64260 , \64261 );
xor \U$64954 ( \65371 , \65370 , \64388 );
_DC gff24 ( \65372_nGff24 , \65371 , \65019 );
buf \U$64955 ( \65373 , \65372_nGff24 );
xor \U$64956 ( \65374 , \64263 , \64264 );
xor \U$64957 ( \65375 , \65374 , \64385 );
_DC gff21 ( \65376_nGff21 , \65375 , \65019 );
buf \U$64958 ( \65377 , \65376_nGff21 );
xor \U$64959 ( \65378 , \64266 , \64267 );
xor \U$64960 ( \65379 , \65378 , \64382 );
_DC gec14 ( \65380_nGec14 , \65379 , \65019 );
buf \U$64961 ( \65381 , \65380_nGec14 );
xor \U$64962 ( \65382 , \64269 , \64270 );
xor \U$64963 ( \65383 , \65382 , \64379 );
_DC gd7a5 ( \65384_nGd7a5 , \65383 , \65019 );
buf \U$64964 ( \65385 , \65384_nGd7a5 );
xor \U$64965 ( \65386 , \64272 , \64273 );
xor \U$64966 ( \65387 , \65386 , \64376 );
_DC gc4a8 ( \65388_nGc4a8 , \65387 , \65019 );
buf \U$64967 ( \65389 , \65388_nGc4a8 );
xor \U$64968 ( \65390 , \64275 , \64276 );
xor \U$64969 ( \65391 , \65390 , \64373 );
_DC gb321 ( \65392_nGb321 , \65391 , \65019 );
buf \U$64970 ( \65393 , \65392_nGb321 );
xor \U$64971 ( \65394 , \64278 , \64279 );
xor \U$64972 ( \65395 , \65394 , \64370 );
_DC ga458 ( \65396_nGa458 , \65395 , \65019 );
buf \U$64973 ( \65397 , \65396_nGa458 );
xor \U$64974 ( \65398 , \64281 , \64282 );
xor \U$64975 ( \65399 , \65398 , \64367 );
_DC g93d2 ( \65400_nG93d2 , \65399 , \65019 );
buf \U$64976 ( \65401 , \65400_nG93d2 );
xor \U$64977 ( \65402 , \64284 , \64285 );
xor \U$64978 ( \65403 , \65402 , \64364 );
_DC g88dd ( \65404_nG88dd , \65403 , \65019 );
buf \U$64979 ( \65405 , \65404_nG88dd );
xor \U$64980 ( \65406 , \64287 , \64288 );
xor \U$64981 ( \65407 , \65406 , \64361 );
_DC g7553 ( \65408_nG7553 , \65407 , \65019 );
buf \U$64982 ( \65409 , \65408_nG7553 );
xor \U$64983 ( \65410 , \64290 , \64291 );
xor \U$64984 ( \65411 , \65410 , \64358 );
_DC g6e59 ( \65412_nG6e59 , \65411 , \65019 );
buf \U$64985 ( \65413 , \65412_nG6e59 );
endmodule

